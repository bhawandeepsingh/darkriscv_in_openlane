VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO darkriscv
  CLASS BLOCK ;
  FOREIGN darkriscv ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.835 BY 515.955 ;
  PIN BE[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.100 511.955 480.380 515.955 ;
    END
  END BE[0]
  PIN BE[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.900 511.955 89.180 515.955 ;
    END
  END BE[1]
  PIN BE[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.470 4.000 415.070 ;
    END
  END BE[2]
  PIN BE[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.500 0.000 278.780 4.000 ;
    END
  END BE[3]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 499.570 500.835 500.170 ;
    END
  END CLK
  PIN DADDR[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.870 4.000 89.470 ;
    END
  END DADDR[0]
  PIN DADDR[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.700 511.955 441.980 515.955 ;
    END
  END DADDR[10]
  PIN DADDR[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.900 0.000 353.180 4.000 ;
    END
  END DADDR[11]
  PIN DADDR[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.100 511.955 108.380 515.955 ;
    END
  END DADDR[12]
  PIN DADDR[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.500 0.000 182.780 4.000 ;
    END
  END DADDR[13]
  PIN DADDR[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.500 511.955 422.780 515.955 ;
    END
  END DADDR[14]
  PIN DADDR[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 469.970 500.835 470.570 ;
    END
  END DADDR[15]
  PIN DADDR[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.700 0.000 249.980 4.000 ;
    END
  END DADDR[16]
  PIN DADDR[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 14.870 500.835 15.470 ;
    END
  END DADDR[17]
  PIN DADDR[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.870 4.000 385.470 ;
    END
  END DADDR[18]
  PIN DADDR[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.900 511.955 269.180 515.955 ;
    END
  END DADDR[19]
  PIN DADDR[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.670 4.000 252.270 ;
    END
  END DADDR[1]
  PIN DADDR[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.900 0.000 77.180 4.000 ;
    END
  END DADDR[20]
  PIN DADDR[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.500 0.000 410.780 4.000 ;
    END
  END DADDR[21]
  PIN DADDR[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.270 4.000 207.870 ;
    END
  END DADDR[22]
  PIN DADDR[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.100 511.955 336.380 515.955 ;
    END
  END DADDR[23]
  PIN DADDR[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.500 511.955 146.780 515.955 ;
    END
  END DADDR[24]
  PIN DADDR[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.100 511.955 432.380 515.955 ;
    END
  END DADDR[25]
  PIN DADDR[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.300 511.955 403.580 515.955 ;
    END
  END DADDR[26]
  PIN DADDR[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.670 4.000 104.270 ;
    END
  END DADDR[27]
  PIN DADDR[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.500 0.000 362.780 4.000 ;
    END
  END DADDR[28]
  PIN DADDR[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.900 511.955 41.180 515.955 ;
    END
  END DADDR[29]
  PIN DADDR[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.100 511.955 60.380 515.955 ;
    END
  END DADDR[2]
  PIN DADDR[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.500 0.000 314.780 4.000 ;
    END
  END DADDR[30]
  PIN DADDR[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.270 4.000 59.870 ;
    END
  END DADDR[31]
  PIN DADDR[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.900 511.955 365.180 515.955 ;
    END
  END DADDR[3]
  PIN DADDR[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 292.370 500.835 292.970 ;
    END
  END DADDR[4]
  PIN DADDR[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 99.970 500.835 100.570 ;
    END
  END DADDR[5]
  PIN DADDR[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 440.370 500.835 440.970 ;
    END
  END DADDR[6]
  PIN DADDR[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.270 4.000 355.870 ;
    END
  END DADDR[7]
  PIN DADDR[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.300 0.000 391.580 4.000 ;
    END
  END DADDR[8]
  PIN DADDR[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 395.970 500.835 396.570 ;
    END
  END DADDR[9]
  PIN DATAI[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.070 4.000 296.670 ;
    END
  END DATAI[0]
  PIN DATAI[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 144.370 500.835 144.970 ;
    END
  END DATAI[10]
  PIN DATAI[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.900 511.955 137.180 515.955 ;
    END
  END DATAI[11]
  PIN DATAI[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.700 511.955 21.980 515.955 ;
    END
  END DATAI[12]
  PIN DATAI[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.500 511.955 2.780 515.955 ;
    END
  END DATAI[13]
  PIN DATAI[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.300 0.000 211.580 4.000 ;
    END
  END DATAI[14]
  PIN DATAI[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.100 0.000 420.380 4.000 ;
    END
  END DATAI[15]
  PIN DATAI[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.370 4.000 440.970 ;
    END
  END DATAI[16]
  PIN DATAI[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 425.570 500.835 426.170 ;
    END
  END DATAI[17]
  PIN DATAI[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.300 0.000 163.580 4.000 ;
    END
  END DATAI[18]
  PIN DATAI[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.700 0.000 477.980 4.000 ;
    END
  END DATAI[19]
  PIN DATAI[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.700 0.000 333.980 4.000 ;
    END
  END DATAI[1]
  PIN DATAI[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 410.770 500.835 411.370 ;
    END
  END DATAI[20]
  PIN DATAI[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.500 511.955 98.780 515.955 ;
    END
  END DATAI[21]
  PIN DATAI[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.670 4.000 400.270 ;
    END
  END DATAI[22]
  PIN DATAI[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.300 0.000 295.580 4.000 ;
    END
  END DATAI[23]
  PIN DATAI[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.100 511.955 240.380 515.955 ;
    END
  END DATAI[24]
  PIN DATAI[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.870 4.000 15.470 ;
    END
  END DATAI[25]
  PIN DATAI[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.970 4.000 470.570 ;
    END
  END DATAI[26]
  PIN DATAI[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.270 4.000 281.870 ;
    END
  END DATAI[27]
  PIN DATAI[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.300 511.955 127.580 515.955 ;
    END
  END DATAI[28]
  PIN DATAI[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 88.870 500.835 89.470 ;
    END
  END DATAI[29]
  PIN DATAI[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.500 0.000 38.780 4.000 ;
    END
  END DATAI[2]
  PIN DATAI[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.900 0.000 497.180 4.000 ;
    END
  END DATAI[30]
  PIN DATAI[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 114.770 500.835 115.370 ;
    END
  END DATAI[31]
  PIN DATAI[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.300 511.955 175.580 515.955 ;
    END
  END DATAI[3]
  PIN DATAI[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.300 511.955 355.580 515.955 ;
    END
  END DATAI[4]
  PIN DATAI[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.900 0.000 305.180 4.000 ;
    END
  END DATAI[5]
  PIN DATAI[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.100 0.000 192.380 4.000 ;
    END
  END DATAI[6]
  PIN DATAI[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.300 511.955 259.580 515.955 ;
    END
  END DATAI[7]
  PIN DATAI[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.500 0.000 458.780 4.000 ;
    END
  END DATAI[8]
  PIN DATAI[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.300 0.000 19.580 4.000 ;
    END
  END DATAI[9]
  PIN DATAO[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.470 4.000 267.070 ;
    END
  END DATAO[0]
  PIN DATAO[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.870 4.000 163.470 ;
    END
  END DATAO[10]
  PIN DATAO[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 233.170 500.835 233.770 ;
    END
  END DATAO[11]
  PIN DATAO[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.700 511.955 345.980 515.955 ;
    END
  END DATAO[12]
  PIN DATAO[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.900 511.955 185.180 515.955 ;
    END
  END DATAO[13]
  PIN DATAO[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.500 0.000 230.780 4.000 ;
    END
  END DATAO[14]
  PIN DATAO[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.900 0.000 401.180 4.000 ;
    END
  END DATAO[15]
  PIN DATAO[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.700 0.000 153.980 4.000 ;
    END
  END DATAO[16]
  PIN DATAO[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.300 0.000 439.580 4.000 ;
    END
  END DATAO[17]
  PIN DATAO[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.100 511.955 12.380 515.955 ;
    END
  END DATAO[18]
  PIN DATAO[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.500 511.955 374.780 515.955 ;
    END
  END DATAO[19]
  PIN DATAO[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.100 0.000 144.380 4.000 ;
    END
  END DATAO[1]
  PIN DATAO[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.070 4.000 148.670 ;
    END
  END DATAO[20]
  PIN DATAO[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.070 4.000 370.670 ;
    END
  END DATAO[21]
  PIN DATAO[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.700 511.955 165.980 515.955 ;
    END
  END DATAO[22]
  PIN DATAO[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.100 511.955 156.380 515.955 ;
    END
  END DATAO[23]
  PIN DATAO[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.100 0.000 468.380 4.000 ;
    END
  END DATAO[24]
  PIN DATAO[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.100 0.000 48.380 4.000 ;
    END
  END DATAO[25]
  PIN DATAO[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.100 0.000 324.380 4.000 ;
    END
  END DATAO[26]
  PIN DATAO[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.500 511.955 470.780 515.955 ;
    END
  END DATAO[27]
  PIN DATAO[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 262.770 500.835 263.370 ;
    END
  END DATAO[28]
  PIN DATAO[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.300 0.000 343.580 4.000 ;
    END
  END DATAO[29]
  PIN DATAO[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.700 0.000 285.980 4.000 ;
    END
  END DATAO[2]
  PIN DATAO[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.500 0.000 86.780 4.000 ;
    END
  END DATAO[30]
  PIN DATAO[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.700 0.000 201.980 4.000 ;
    END
  END DATAO[31]
  PIN DATAO[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 351.570 500.835 352.170 ;
    END
  END DATAO[3]
  PIN DATAO[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 59.270 500.835 59.870 ;
    END
  END DATAO[4]
  PIN DATAO[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.900 0.000 449.180 4.000 ;
    END
  END DATAO[5]
  PIN DATAO[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.300 511.955 79.580 515.955 ;
    END
  END DATAO[6]
  PIN DATAO[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.900 0.000 173.180 4.000 ;
    END
  END DATAO[7]
  PIN DATAO[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.670 4.000 178.270 ;
    END
  END DATAO[8]
  PIN DATAO[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 277.570 500.835 278.170 ;
    END
  END DATAO[9]
  PIN DEBUG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.900 0.000 125.180 4.000 ;
    END
  END DEBUG[0]
  PIN DEBUG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.070 4.000 222.670 ;
    END
  END DEBUG[1]
  PIN DEBUG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.300 0.000 259.580 4.000 ;
    END
  END DEBUG[2]
  PIN DEBUG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.670 4.000 326.270 ;
    END
  END DEBUG[3]
  PIN HLT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.470 4.000 193.070 ;
    END
  END HLT
  PIN IADDR[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 203.570 500.835 204.170 ;
    END
  END IADDR[0]
  PIN IADDR[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.700 511.955 249.980 515.955 ;
    END
  END IADDR[10]
  PIN IADDR[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.870 4.000 237.470 ;
    END
  END IADDR[11]
  PIN IADDR[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.500 511.955 278.780 515.955 ;
    END
  END IADDR[12]
  PIN IADDR[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.900 511.955 497.180 515.955 ;
    END
  END IADDR[13]
  PIN IADDR[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.470 4.000 45.070 ;
    END
  END IADDR[14]
  PIN IADDR[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 218.370 500.835 218.970 ;
    END
  END IADDR[15]
  PIN IADDR[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.570 4.000 500.170 ;
    END
  END IADDR[16]
  PIN IADDR[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.900 0.000 29.180 4.000 ;
    END
  END IADDR[17]
  PIN IADDR[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.700 0.000 9.980 4.000 ;
    END
  END IADDR[18]
  PIN IADDR[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.270 4.000 133.870 ;
    END
  END IADDR[19]
  PIN IADDR[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 188.770 500.835 189.370 ;
    END
  END IADDR[1]
  PIN IADDR[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.500 511.955 326.780 515.955 ;
    END
  END IADDR[20]
  PIN IADDR[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 307.170 500.835 307.770 ;
    END
  END IADDR[21]
  PIN IADDR[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 484.770 500.835 485.370 ;
    END
  END IADDR[22]
  PIN IADDR[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.900 0.000 269.180 4.000 ;
    END
  END IADDR[23]
  PIN IADDR[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.100 0.000 372.380 4.000 ;
    END
  END IADDR[24]
  PIN IADDR[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 129.570 500.835 130.170 ;
    END
  END IADDR[25]
  PIN IADDR[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 74.070 500.835 74.670 ;
    END
  END IADDR[26]
  PIN IADDR[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.500 511.955 194.780 515.955 ;
    END
  END IADDR[27]
  PIN IADDR[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.700 511.955 69.980 515.955 ;
    END
  END IADDR[28]
  PIN IADDR[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.500 511.955 50.780 515.955 ;
    END
  END IADDR[29]
  PIN IADDR[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.700 511.955 393.980 515.955 ;
    END
  END IADDR[2]
  PIN IADDR[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.500 0.000 134.780 4.000 ;
    END
  END IADDR[30]
  PIN IADDR[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 321.970 500.835 322.570 ;
    END
  END IADDR[31]
  PIN IADDR[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.470 4.000 341.070 ;
    END
  END IADDR[3]
  PIN IADDR[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.300 511.955 31.580 515.955 ;
    END
  END IADDR[4]
  PIN IADDR[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.700 511.955 117.980 515.955 ;
    END
  END IADDR[5]
  PIN IADDR[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.100 0.000 240.380 4.000 ;
    END
  END IADDR[6]
  PIN IADDR[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.700 511.955 489.980 515.955 ;
    END
  END IADDR[7]
  PIN IADDR[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 159.170 500.835 159.770 ;
    END
  END IADDR[8]
  PIN IADDR[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.070 4.000 74.670 ;
    END
  END IADDR[9]
  PIN IDATA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.500 511.955 230.780 515.955 ;
    END
  END IDATA[0]
  PIN IDATA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.470 4.000 119.070 ;
    END
  END IDATA[10]
  PIN IDATA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.300 0.000 115.580 4.000 ;
    END
  END IDATA[11]
  PIN IDATA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 381.170 500.835 381.770 ;
    END
  END IDATA[12]
  PIN IDATA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 336.770 500.835 337.370 ;
    END
  END IDATA[13]
  PIN IDATA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.300 0.000 67.580 4.000 ;
    END
  END IDATA[14]
  PIN IDATA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.900 511.955 413.180 515.955 ;
    END
  END IDATA[15]
  PIN IDATA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.700 0.000 57.980 4.000 ;
    END
  END IDATA[16]
  PIN IDATA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 44.470 500.835 45.070 ;
    END
  END IDATA[17]
  PIN IDATA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.700 511.955 213.980 515.955 ;
    END
  END IDATA[18]
  PIN IDATA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 247.970 500.835 248.570 ;
    END
  END IDATA[19]
  PIN IDATA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 366.370 500.835 366.970 ;
    END
  END IDATA[1]
  PIN IDATA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.300 511.955 451.580 515.955 ;
    END
  END IDATA[20]
  PIN IDATA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.100 511.955 384.380 515.955 ;
    END
  END IDATA[21]
  PIN IDATA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.500 0.000 2.780 4.000 ;
    END
  END IDATA[22]
  PIN IDATA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.700 0.000 105.980 4.000 ;
    END
  END IDATA[23]
  PIN IDATA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.900 0.000 221.180 4.000 ;
    END
  END IDATA[24]
  PIN IDATA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.700 511.955 297.980 515.955 ;
    END
  END IDATA[25]
  PIN IDATA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.100 0.000 96.380 4.000 ;
    END
  END IDATA[26]
  PIN IDATA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.670 4.000 30.270 ;
    END
  END IDATA[27]
  PIN IDATA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.900 511.955 461.180 515.955 ;
    END
  END IDATA[28]
  PIN IDATA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.100 511.955 204.380 515.955 ;
    END
  END IDATA[29]
  PIN IDATA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 173.970 500.835 174.570 ;
    END
  END IDATA[2]
  PIN IDATA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.870 4.000 311.470 ;
    END
  END IDATA[30]
  PIN IDATA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.300 511.955 307.580 515.955 ;
    END
  END IDATA[31]
  PIN IDATA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 29.670 500.835 30.270 ;
    END
  END IDATA[3]
  PIN IDATA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.300 0.000 487.580 4.000 ;
    END
  END IDATA[4]
  PIN IDATA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.100 511.955 288.380 515.955 ;
    END
  END IDATA[5]
  PIN IDATA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.770 4.000 485.370 ;
    END
  END IDATA[6]
  PIN IDATA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.570 4.000 426.170 ;
    END
  END IDATA[7]
  PIN IDATA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.900 511.955 221.180 515.955 ;
    END
  END IDATA[8]
  PIN IDATA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.900 511.955 317.180 515.955 ;
    END
  END IDATA[9]
  PIN IDLE
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.700 0.000 429.980 4.000 ;
    END
  END IDLE
  PIN RD
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.835 455.170 500.835 455.770 ;
    END
  END RD
  PIN RES
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.170 4.000 455.770 ;
    END
  END RES
  PIN WR
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.700 0.000 381.980 4.000 ;
    END
  END WR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 482.080 13.080 483.680 499.740 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.480 13.080 330.080 499.740 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.880 13.080 176.480 499.740 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.280 13.080 22.880 499.740 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.280 13.080 406.880 499.740 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.680 13.080 253.280 499.740 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 98.080 13.080 99.680 499.740 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.760 13.235 494.880 499.585 ;
      LAYER met1 ;
        RECT 2.480 12.635 497.200 500.555 ;
      LAYER met2 ;
        RECT 3.060 511.675 11.820 511.955 ;
        RECT 12.660 511.675 21.420 511.955 ;
        RECT 22.260 511.675 31.020 511.955 ;
        RECT 31.860 511.675 40.620 511.955 ;
        RECT 41.460 511.675 50.220 511.955 ;
        RECT 51.060 511.675 59.820 511.955 ;
        RECT 60.660 511.675 69.420 511.955 ;
        RECT 70.260 511.675 79.020 511.955 ;
        RECT 79.860 511.675 88.620 511.955 ;
        RECT 89.460 511.675 98.220 511.955 ;
        RECT 99.060 511.675 107.820 511.955 ;
        RECT 108.660 511.675 117.420 511.955 ;
        RECT 118.260 511.675 127.020 511.955 ;
        RECT 127.860 511.675 136.620 511.955 ;
        RECT 137.460 511.675 146.220 511.955 ;
        RECT 147.060 511.675 155.820 511.955 ;
        RECT 156.660 511.675 165.420 511.955 ;
        RECT 166.260 511.675 175.020 511.955 ;
        RECT 175.860 511.675 184.620 511.955 ;
        RECT 185.460 511.675 194.220 511.955 ;
        RECT 195.060 511.675 203.820 511.955 ;
        RECT 204.660 511.675 213.420 511.955 ;
        RECT 214.260 511.675 220.620 511.955 ;
        RECT 221.460 511.675 230.220 511.955 ;
        RECT 231.060 511.675 239.820 511.955 ;
        RECT 240.660 511.675 249.420 511.955 ;
        RECT 250.260 511.675 259.020 511.955 ;
        RECT 259.860 511.675 268.620 511.955 ;
        RECT 269.460 511.675 278.220 511.955 ;
        RECT 279.060 511.675 287.820 511.955 ;
        RECT 288.660 511.675 297.420 511.955 ;
        RECT 298.260 511.675 307.020 511.955 ;
        RECT 307.860 511.675 316.620 511.955 ;
        RECT 317.460 511.675 326.220 511.955 ;
        RECT 327.060 511.675 335.820 511.955 ;
        RECT 336.660 511.675 345.420 511.955 ;
        RECT 346.260 511.675 355.020 511.955 ;
        RECT 355.860 511.675 364.620 511.955 ;
        RECT 365.460 511.675 374.220 511.955 ;
        RECT 375.060 511.675 383.820 511.955 ;
        RECT 384.660 511.675 393.420 511.955 ;
        RECT 394.260 511.675 403.020 511.955 ;
        RECT 403.860 511.675 412.620 511.955 ;
        RECT 413.460 511.675 422.220 511.955 ;
        RECT 423.060 511.675 431.820 511.955 ;
        RECT 432.660 511.675 441.420 511.955 ;
        RECT 442.260 511.675 451.020 511.955 ;
        RECT 451.860 511.675 460.620 511.955 ;
        RECT 461.460 511.675 470.220 511.955 ;
        RECT 471.060 511.675 479.820 511.955 ;
        RECT 480.660 511.675 489.420 511.955 ;
        RECT 490.260 511.675 496.620 511.955 ;
        RECT 2.510 4.280 497.170 511.675 ;
        RECT 3.060 4.000 9.420 4.280 ;
        RECT 10.260 4.000 19.020 4.280 ;
        RECT 19.860 4.000 28.620 4.280 ;
        RECT 29.460 4.000 38.220 4.280 ;
        RECT 39.060 4.000 47.820 4.280 ;
        RECT 48.660 4.000 57.420 4.280 ;
        RECT 58.260 4.000 67.020 4.280 ;
        RECT 67.860 4.000 76.620 4.280 ;
        RECT 77.460 4.000 86.220 4.280 ;
        RECT 87.060 4.000 95.820 4.280 ;
        RECT 96.660 4.000 105.420 4.280 ;
        RECT 106.260 4.000 115.020 4.280 ;
        RECT 115.860 4.000 124.620 4.280 ;
        RECT 125.460 4.000 134.220 4.280 ;
        RECT 135.060 4.000 143.820 4.280 ;
        RECT 144.660 4.000 153.420 4.280 ;
        RECT 154.260 4.000 163.020 4.280 ;
        RECT 163.860 4.000 172.620 4.280 ;
        RECT 173.460 4.000 182.220 4.280 ;
        RECT 183.060 4.000 191.820 4.280 ;
        RECT 192.660 4.000 201.420 4.280 ;
        RECT 202.260 4.000 211.020 4.280 ;
        RECT 211.860 4.000 220.620 4.280 ;
        RECT 221.460 4.000 230.220 4.280 ;
        RECT 231.060 4.000 239.820 4.280 ;
        RECT 240.660 4.000 249.420 4.280 ;
        RECT 250.260 4.000 259.020 4.280 ;
        RECT 259.860 4.000 268.620 4.280 ;
        RECT 269.460 4.000 278.220 4.280 ;
        RECT 279.060 4.000 285.420 4.280 ;
        RECT 286.260 4.000 295.020 4.280 ;
        RECT 295.860 4.000 304.620 4.280 ;
        RECT 305.460 4.000 314.220 4.280 ;
        RECT 315.060 4.000 323.820 4.280 ;
        RECT 324.660 4.000 333.420 4.280 ;
        RECT 334.260 4.000 343.020 4.280 ;
        RECT 343.860 4.000 352.620 4.280 ;
        RECT 353.460 4.000 362.220 4.280 ;
        RECT 363.060 4.000 371.820 4.280 ;
        RECT 372.660 4.000 381.420 4.280 ;
        RECT 382.260 4.000 391.020 4.280 ;
        RECT 391.860 4.000 400.620 4.280 ;
        RECT 401.460 4.000 410.220 4.280 ;
        RECT 411.060 4.000 419.820 4.280 ;
        RECT 420.660 4.000 429.420 4.280 ;
        RECT 430.260 4.000 439.020 4.280 ;
        RECT 439.860 4.000 448.620 4.280 ;
        RECT 449.460 4.000 458.220 4.280 ;
        RECT 459.060 4.000 467.820 4.280 ;
        RECT 468.660 4.000 477.420 4.280 ;
        RECT 478.260 4.000 487.020 4.280 ;
        RECT 487.860 4.000 496.620 4.280 ;
      LAYER met3 ;
        RECT 4.400 499.170 496.435 500.035 ;
        RECT 4.000 485.770 496.835 499.170 ;
        RECT 4.400 484.370 496.435 485.770 ;
        RECT 4.000 470.970 496.835 484.370 ;
        RECT 4.400 469.570 496.435 470.970 ;
        RECT 4.000 456.170 496.835 469.570 ;
        RECT 4.400 454.770 496.435 456.170 ;
        RECT 4.000 441.370 496.835 454.770 ;
        RECT 4.400 439.970 496.435 441.370 ;
        RECT 4.000 426.570 496.835 439.970 ;
        RECT 4.400 425.170 496.435 426.570 ;
        RECT 4.000 415.470 496.835 425.170 ;
        RECT 4.400 414.070 496.835 415.470 ;
        RECT 4.000 411.770 496.835 414.070 ;
        RECT 4.000 410.370 496.435 411.770 ;
        RECT 4.000 400.670 496.835 410.370 ;
        RECT 4.400 399.270 496.835 400.670 ;
        RECT 4.000 396.970 496.835 399.270 ;
        RECT 4.000 395.570 496.435 396.970 ;
        RECT 4.000 385.870 496.835 395.570 ;
        RECT 4.400 384.470 496.835 385.870 ;
        RECT 4.000 382.170 496.835 384.470 ;
        RECT 4.000 380.770 496.435 382.170 ;
        RECT 4.000 371.070 496.835 380.770 ;
        RECT 4.400 369.670 496.835 371.070 ;
        RECT 4.000 367.370 496.835 369.670 ;
        RECT 4.000 365.970 496.435 367.370 ;
        RECT 4.000 356.270 496.835 365.970 ;
        RECT 4.400 354.870 496.835 356.270 ;
        RECT 4.000 352.570 496.835 354.870 ;
        RECT 4.000 351.170 496.435 352.570 ;
        RECT 4.000 341.470 496.835 351.170 ;
        RECT 4.400 340.070 496.835 341.470 ;
        RECT 4.000 337.770 496.835 340.070 ;
        RECT 4.000 336.370 496.435 337.770 ;
        RECT 4.000 326.670 496.835 336.370 ;
        RECT 4.400 325.270 496.835 326.670 ;
        RECT 4.000 322.970 496.835 325.270 ;
        RECT 4.000 321.570 496.435 322.970 ;
        RECT 4.000 311.870 496.835 321.570 ;
        RECT 4.400 310.470 496.835 311.870 ;
        RECT 4.000 308.170 496.835 310.470 ;
        RECT 4.000 306.770 496.435 308.170 ;
        RECT 4.000 297.070 496.835 306.770 ;
        RECT 4.400 295.670 496.835 297.070 ;
        RECT 4.000 293.370 496.835 295.670 ;
        RECT 4.000 291.970 496.435 293.370 ;
        RECT 4.000 282.270 496.835 291.970 ;
        RECT 4.400 280.870 496.835 282.270 ;
        RECT 4.000 278.570 496.835 280.870 ;
        RECT 4.000 277.170 496.435 278.570 ;
        RECT 4.000 267.470 496.835 277.170 ;
        RECT 4.400 266.070 496.835 267.470 ;
        RECT 4.000 263.770 496.835 266.070 ;
        RECT 4.000 262.370 496.435 263.770 ;
        RECT 4.000 252.670 496.835 262.370 ;
        RECT 4.400 251.270 496.835 252.670 ;
        RECT 4.000 248.970 496.835 251.270 ;
        RECT 4.000 247.570 496.435 248.970 ;
        RECT 4.000 237.870 496.835 247.570 ;
        RECT 4.400 236.470 496.835 237.870 ;
        RECT 4.000 234.170 496.835 236.470 ;
        RECT 4.000 232.770 496.435 234.170 ;
        RECT 4.000 223.070 496.835 232.770 ;
        RECT 4.400 221.670 496.835 223.070 ;
        RECT 4.000 219.370 496.835 221.670 ;
        RECT 4.000 217.970 496.435 219.370 ;
        RECT 4.000 208.270 496.835 217.970 ;
        RECT 4.400 206.870 496.835 208.270 ;
        RECT 4.000 204.570 496.835 206.870 ;
        RECT 4.000 203.170 496.435 204.570 ;
        RECT 4.000 193.470 496.835 203.170 ;
        RECT 4.400 192.070 496.835 193.470 ;
        RECT 4.000 189.770 496.835 192.070 ;
        RECT 4.000 188.370 496.435 189.770 ;
        RECT 4.000 178.670 496.835 188.370 ;
        RECT 4.400 177.270 496.835 178.670 ;
        RECT 4.000 174.970 496.835 177.270 ;
        RECT 4.000 173.570 496.435 174.970 ;
        RECT 4.000 163.870 496.835 173.570 ;
        RECT 4.400 162.470 496.835 163.870 ;
        RECT 4.000 160.170 496.835 162.470 ;
        RECT 4.000 158.770 496.435 160.170 ;
        RECT 4.000 149.070 496.835 158.770 ;
        RECT 4.400 147.670 496.835 149.070 ;
        RECT 4.000 145.370 496.835 147.670 ;
        RECT 4.000 143.970 496.435 145.370 ;
        RECT 4.000 134.270 496.835 143.970 ;
        RECT 4.400 132.870 496.835 134.270 ;
        RECT 4.000 130.570 496.835 132.870 ;
        RECT 4.000 129.170 496.435 130.570 ;
        RECT 4.000 119.470 496.835 129.170 ;
        RECT 4.400 118.070 496.835 119.470 ;
        RECT 4.000 115.770 496.835 118.070 ;
        RECT 4.000 114.370 496.435 115.770 ;
        RECT 4.000 104.670 496.835 114.370 ;
        RECT 4.400 103.270 496.835 104.670 ;
        RECT 4.000 100.970 496.835 103.270 ;
        RECT 4.000 99.570 496.435 100.970 ;
        RECT 4.000 89.870 496.835 99.570 ;
        RECT 4.400 88.470 496.435 89.870 ;
        RECT 4.000 75.070 496.835 88.470 ;
        RECT 4.400 73.670 496.435 75.070 ;
        RECT 4.000 60.270 496.835 73.670 ;
        RECT 4.400 58.870 496.435 60.270 ;
        RECT 4.000 45.470 496.835 58.870 ;
        RECT 4.400 44.070 496.435 45.470 ;
        RECT 4.000 30.670 496.835 44.070 ;
        RECT 4.400 29.270 496.435 30.670 ;
        RECT 4.000 15.870 496.835 29.270 ;
        RECT 4.400 14.470 496.435 15.870 ;
        RECT 4.000 13.155 496.835 14.470 ;
      LAYER met4 ;
        RECT 23.355 14.265 97.680 498.555 ;
        RECT 100.080 14.265 174.480 498.555 ;
        RECT 176.880 14.265 251.280 498.555 ;
        RECT 253.680 14.265 328.080 498.555 ;
        RECT 330.480 14.265 404.880 498.555 ;
        RECT 407.280 14.265 481.680 498.555 ;
        RECT 484.080 14.265 489.285 498.555 ;
  END
END darkriscv
END LIBRARY

