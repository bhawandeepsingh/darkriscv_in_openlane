module user_project_wrapper (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    vccd1,
    vssd1,
    vccd2,
    vssd2,
    vdda1,
    vssa1,
    vdda2,
    vssa2,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input vccd1;
 input vssd1;
 input vccd2;
 input vssd2;
 input vdda1;
 input vssa1;
 input vdda2;
 input vssa2;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 sky130_fd_sc_hd__inv_2 _07037_ (.A(\design_top.DACK[0] ),
    .Y(_01111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07038_ (.A(\design_top.core0.FLUSH[1] ),
    .Y(_04615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07039_ (.A(\design_top.core0.FLUSH[0] ),
    .Y(_04616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _07040_ (.A(_04615_),
    .B(_04616_),
    .C(\design_top.core0.XLCC ),
    .X(_04617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07041_ (.A(_04617_),
    .X(io_out[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07042_ (.A1(_01111_),
    .A2(\design_top.DACK[1] ),
    .B1(io_out[12]),
    .Y(_04618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07043_ (.A(_04618_),
    .Y(_04619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07044_ (.A(_04619_),
    .X(_04620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07045_ (.A(\design_top.core0.XJALR ),
    .Y(_04621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07046_ (.A(\design_top.core0.XJAL ),
    .Y(_04622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07047_ (.A(_00900_),
    .Y(_04623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07048_ (.A(\design_top.core0.FCT3[2] ),
    .Y(_04624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07049_ (.A(\design_top.core0.FCT3[1] ),
    .B(\design_top.core0.FCT3[0] ),
    .X(_04625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07050_ (.A(_04625_),
    .X(_00539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07051_ (.A(_00304_),
    .Y(_04626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07052_ (.A1(_00323_),
    .A2(_04626_),
    .B1(_00320_),
    .B2(_00304_),
    .X(_04627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _07053_ (.A(_00833_),
    .B(_04627_),
    .Y(_01587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _07054_ (.A1(_00833_),
    .A2(_04627_),
    .B1(_01587_),
    .Y(_04628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07055_ (.A(_04628_),
    .X(_04629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07056_ (.A(_00756_),
    .B(_00500_),
    .X(_04630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07057_ (.A(_00756_),
    .B(_00500_),
    .Y(_00758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07058_ (.A(_04630_),
    .B(_00758_),
    .Y(_00876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07059_ (.A(_00876_),
    .Y(_04631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07060_ (.A(_00512_),
    .X(_04632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _07061_ (.A(_00772_),
    .B(_04632_),
    .Y(_00773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _07062_ (.A1(_00772_),
    .A2(_04632_),
    .B1(_00773_),
    .Y(_04633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07063_ (.A(_00518_),
    .X(_04634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07064_ (.A(_04634_),
    .B(_00781_),
    .Y(_01914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07065_ (.A1(_04634_),
    .A2(_00781_),
    .B1(_01914_),
    .Y(_00873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07066_ (.A(_00873_),
    .Y(_04635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _07067_ (.A(_00506_),
    .B(_00765_),
    .Y(_00766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07068_ (.A(_00506_),
    .B(_00765_),
    .Y(_01960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07069_ (.A(_01960_),
    .Y(_04636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07070_ (.A(_00766_),
    .B(_04636_),
    .X(_04637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07071_ (.A(_04637_),
    .Y(_04638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07072_ (.A(_04631_),
    .B(_04633_),
    .C(_04635_),
    .D(_04638_),
    .X(_04639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07073_ (.A(_00530_),
    .B(_00792_),
    .Y(_01845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07074_ (.A1(_00530_),
    .A2(_00792_),
    .B1(_01845_),
    .Y(_04640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07075_ (.A(_04640_),
    .Y(_04641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07076_ (.A(_00359_),
    .X(_04642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _07077_ (.A(_00799_),
    .B(_04642_),
    .Y(_00800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _07078_ (.A1(_00799_),
    .A2(_04642_),
    .B1(_00800_),
    .Y(_04643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07079_ (.A(_00352_),
    .X(_04644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07080_ (.A(_04644_),
    .B(_00808_),
    .Y(_01758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07081_ (.A1(_04644_),
    .A2(_00808_),
    .B1(_01758_),
    .Y(_04645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07082_ (.A(_04645_),
    .Y(_04646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _07083_ (.A(_00524_),
    .B(_00783_),
    .Y(_00784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _07084_ (.A1(_00524_),
    .A2(_00783_),
    .B1(_00784_),
    .Y(_04647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07085_ (.A(_04641_),
    .B(_04643_),
    .C(_04646_),
    .D(_04647_),
    .X(_04648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07086_ (.A(_00816_),
    .X(_04649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07087_ (.A1(_00341_),
    .A2(_04626_),
    .B1(_00338_),
    .B2(_00304_),
    .X(_04650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _07088_ (.A(_00816_),
    .B(_04650_),
    .Y(_00817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _07089_ (.A1(_04649_),
    .A2(_04650_),
    .B1(_00817_),
    .Y(_04651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07090_ (.A(_04629_),
    .B(_04639_),
    .C(_04648_),
    .D(_04651_),
    .X(_04652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07091_ (.A(_00482_),
    .B(_00732_),
    .Y(_02053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07092_ (.A1(_00482_),
    .A2(_00732_),
    .B1(_02053_),
    .Y(_04653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07093_ (.A(_04653_),
    .X(_02054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07094_ (.A(_02054_),
    .Y(_04654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07095_ (.A(_00488_),
    .X(_04655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07096_ (.A(_04655_),
    .X(_04656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07097_ (.A(_04655_),
    .B(_00740_),
    .Y(_00742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07098_ (.A1(_04656_),
    .A2(_00740_),
    .B1(_00742_),
    .Y(_00878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07099_ (.A(_00878_),
    .Y(_04657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07100_ (.A(_00494_),
    .X(_04658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07101_ (.A(_04658_),
    .B(_00749_),
    .Y(_02005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07102_ (.A1(_04658_),
    .A2(_00749_),
    .B1(_02005_),
    .Y(_04659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07103_ (.A(_04659_),
    .X(_00877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07104_ (.A(_00877_),
    .Y(_04660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07105_ (.A(_00825_),
    .Y(_04661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07106_ (.A(_00317_),
    .Y(_04662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07107_ (.A(_04662_),
    .X(_04663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07108_ (.A1(_00825_),
    .A2(_00317_),
    .B1(_04661_),
    .B2(_04663_),
    .X(_04664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07109_ (.A(_00476_),
    .X(_04665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07110_ (.A(_04665_),
    .B(_00723_),
    .Y(_00725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07111_ (.A1(_04665_),
    .A2(_00723_),
    .B1(_00725_),
    .Y(_00879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07112_ (.A(_00879_),
    .Y(_04666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07113_ (.A(_04664_),
    .B(_04666_),
    .X(_04667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07114_ (.A(_04654_),
    .B(_04657_),
    .C(_04660_),
    .D(_04667_),
    .X(_04668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07115_ (.A(_00404_),
    .B(_00626_),
    .Y(_00628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07116_ (.A1(_00404_),
    .A2(_00626_),
    .B1(_00628_),
    .Y(_00890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07117_ (.A(_00890_),
    .Y(_04669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07118_ (.A(_00410_),
    .B(_00635_),
    .Y(_02302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07119_ (.A1(_00410_),
    .A2(_00635_),
    .B1(_02302_),
    .Y(_04670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07120_ (.A(_04670_),
    .Y(_04671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07121_ (.A(_00416_),
    .X(_04672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07122_ (.A(_04672_),
    .B(_00643_),
    .Y(_00645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07123_ (.A1(_04672_),
    .A2(_00643_),
    .B1(_00645_),
    .Y(_00888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07124_ (.A(_00888_),
    .Y(_04673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07125_ (.A(_00422_),
    .X(_04674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07126_ (.A(_04674_),
    .B(_00652_),
    .Y(_02260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07127_ (.A1(_04674_),
    .A2(_00652_),
    .B1(_02260_),
    .Y(_04675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4b_2 _07128_ (.A(_04669_),
    .B(_04671_),
    .C(_04673_),
    .D_N(_04675_),
    .X(_04676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07129_ (.A(_00464_),
    .X(_04677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07130_ (.A(_04677_),
    .X(_04678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07131_ (.A(_04677_),
    .B(_00711_),
    .Y(_00713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07132_ (.A1(_04678_),
    .A2(_00711_),
    .B1(_00713_),
    .Y(_00881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07133_ (.A(_00881_),
    .Y(_04679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07134_ (.A(_00452_),
    .X(_04680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07135_ (.A(_04680_),
    .B(_00694_),
    .Y(_00696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07136_ (.A1(_04680_),
    .A2(_00694_),
    .B1(_00696_),
    .Y(_00882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07137_ (.A(_00882_),
    .Y(_04681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07138_ (.A(_00470_),
    .X(_04682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07139_ (.A(_00720_),
    .B(_00470_),
    .Y(_02094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07140_ (.A1(_00720_),
    .A2(_04682_),
    .B1(_02094_),
    .Y(_00880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07141_ (.A(_00880_),
    .Y(_04683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _07142_ (.A(_00458_),
    .B(_00703_),
    .Y(_00704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07143_ (.A(_00458_),
    .B(_00703_),
    .Y(_02136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07144_ (.A(_02136_),
    .Y(_04684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07145_ (.A(_00704_),
    .B(_04684_),
    .X(_04685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07146_ (.A(_04685_),
    .Y(_04686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07147_ (.A(_04679_),
    .B(_04681_),
    .C(_04683_),
    .D(_04686_),
    .X(_04687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07148_ (.A(_00434_),
    .X(_04688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07149_ (.A(_04688_),
    .B(_00669_),
    .Y(_02220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07150_ (.A1(_04688_),
    .A2(_00669_),
    .B1(_02220_),
    .Y(_04689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07151_ (.A(_04689_),
    .Y(_04690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07152_ (.A(_00428_),
    .X(_04691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07153_ (.A(_04691_),
    .B(_00660_),
    .Y(_00662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07154_ (.A1(_04691_),
    .A2(_00660_),
    .B1(_00662_),
    .Y(_00886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07155_ (.A(_00886_),
    .Y(_04692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07156_ (.A(_00446_),
    .X(_04693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07157_ (.A(_04693_),
    .B(_00686_),
    .Y(_02178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07158_ (.A1(_04693_),
    .A2(_00686_),
    .B1(_02178_),
    .Y(_04694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07159_ (.A(_04694_),
    .Y(_04695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07160_ (.A(_00440_),
    .X(_04696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07161_ (.A(_04696_),
    .X(_04697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07162_ (.A(_04696_),
    .B(_00677_),
    .Y(_00679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07163_ (.A1(_04697_),
    .A2(_00677_),
    .B1(_00679_),
    .Y(_00884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07164_ (.A(_00884_),
    .Y(_04698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07165_ (.A(_04690_),
    .B(_04692_),
    .C(_04695_),
    .D(_04698_),
    .X(_04699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07166_ (.A(_00386_),
    .B(_00600_),
    .Y(_00602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07167_ (.A1(_00386_),
    .A2(_00600_),
    .B1(_00602_),
    .Y(_00893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07168_ (.A(_00893_),
    .Y(_04700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07169_ (.A(_00381_),
    .Y(_04701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _07170_ (.A(_04701_),
    .B(_00591_),
    .Y(_00592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _07171_ (.A1(_04701_),
    .A2(_00591_),
    .B1(_00592_),
    .Y(_04702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _07172_ (.A(_00398_),
    .B(_00618_),
    .Y(_00619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _07173_ (.A1(_00398_),
    .A2(_00618_),
    .B1(_00619_),
    .Y(_04703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07174_ (.A(_00392_),
    .X(_04704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07175_ (.A(_00392_),
    .B(_00609_),
    .Y(_00611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07176_ (.A1(_04704_),
    .A2(_00609_),
    .B1(_00611_),
    .Y(_00892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07177_ (.A(_00892_),
    .Y(_04705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07178_ (.A(_04700_),
    .B(_04702_),
    .C(_04703_),
    .D(_04705_),
    .X(_04706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07179_ (.A(_04676_),
    .B(_04687_),
    .C(_04699_),
    .D(_04706_),
    .X(_04707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _07180_ (.A(_04652_),
    .B(_04668_),
    .C(_04707_),
    .X(_04708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _07181_ (.A(_04624_),
    .B(_00539_),
    .C(_04708_),
    .X(_04709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07182_ (.A1(_04623_),
    .A2(_04709_),
    .B1(\design_top.core0.XBCC ),
    .Y(_04710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07183_ (.A(\design_top.core0.FLUSH[1] ),
    .B(\design_top.core0.FLUSH[0] ),
    .X(_04711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _07184_ (.A1(_04621_),
    .A2(_04622_),
    .A3(_04710_),
    .B1(_04711_),
    .X(_00901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07185_ (.A(_04620_),
    .B(_00901_),
    .X(_04712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07186_ (.A(_04712_),
    .Y(_04713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07187_ (.A(_02403_),
    .Y(_04714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07188_ (.A(\design_top.core0.XRES ),
    .Y(_04715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07189_ (.A(_04715_),
    .X(_04716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07190_ (.A(_04716_),
    .X(_04717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _07191_ (.A1(io_out[16]),
    .A2(_04713_),
    .B1(_04714_),
    .B2(_04712_),
    .C1(_04717_),
    .X(_04436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07192_ (.A(\design_top.DATAO[31] ),
    .Y(_04718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07193_ (.A(_04718_),
    .X(_04719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07194_ (.A(_04711_),
    .Y(_00309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _07195_ (.A(\design_top.core0.XSCC ),
    .B(_00309_),
    .Y(_04720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07196_ (.A(\design_top.core0.SIMM[30] ),
    .Y(_00387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07197_ (.A(_00386_),
    .X(_04721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07198_ (.A(_04721_),
    .Y(_04722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _07199_ (.A1(\design_top.core0.SIMM[30] ),
    .A2(_04721_),
    .B1(_00387_),
    .B2(_04722_),
    .X(_04723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07200_ (.A(\design_top.core0.SIMM[29] ),
    .X(_04724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _07201_ (.A(\design_top.core0.SIMM[29] ),
    .B(_00392_),
    .Y(_04725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _07202_ (.A1(_04724_),
    .A2(_04704_),
    .B1(_04725_),
    .Y(_04726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07203_ (.A(_04726_),
    .Y(_04727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07204_ (.A(\design_top.core0.SIMM[28] ),
    .Y(_00399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07205_ (.A(_00398_),
    .Y(_04728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07206_ (.A(\design_top.core0.SIMM[28] ),
    .X(_04729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07207_ (.A1(_00399_),
    .A2(_04728_),
    .B1(_04729_),
    .B2(_00398_),
    .X(_04730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07208_ (.A(_04730_),
    .Y(_04731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07209_ (.A(\design_top.core0.SIMM[27] ),
    .Y(_04732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07210_ (.A(_04732_),
    .X(_00405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07211_ (.A(_00404_),
    .Y(_04733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07212_ (.A(\design_top.core0.SIMM[26] ),
    .Y(_04734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07213_ (.A(_00410_),
    .Y(_04735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _07214_ (.A1(_04732_),
    .A2(_04733_),
    .B1(_04734_),
    .C1(_04735_),
    .X(_04736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _07215_ (.A1(\design_top.core0.SIMM[27] ),
    .A2(_00404_),
    .B1(_04732_),
    .B2(_04733_),
    .X(_04737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _07216_ (.A1(\design_top.core0.SIMM[26] ),
    .A2(_00410_),
    .B1(_04734_),
    .B2(_04735_),
    .X(_04738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07217_ (.A(_04737_),
    .B(_04738_),
    .X(_04739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _07218_ (.A1(\design_top.core0.SIMM[25] ),
    .A2(_00416_),
    .B1(\design_top.core0.SIMM[24] ),
    .B2(_04674_),
    .X(_04740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07219_ (.A1(\design_top.core0.SIMM[25] ),
    .A2(_00416_),
    .B1(_04740_),
    .Y(_04741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07220_ (.A(_04739_),
    .B(_04741_),
    .X(_04742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07221_ (.A(\design_top.core0.SIMM[25] ),
    .Y(_00417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07222_ (.A(_00416_),
    .Y(_04743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07223_ (.A1(_00417_),
    .A2(_04743_),
    .B1(\design_top.core0.SIMM[25] ),
    .B2(_00416_),
    .X(_04744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07224_ (.A(_04744_),
    .Y(_04745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07225_ (.A(\design_top.core0.SIMM[24] ),
    .Y(_00423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07226_ (.A(_00422_),
    .Y(_04746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07227_ (.A1(_00423_),
    .A2(_04746_),
    .B1(\design_top.core0.SIMM[24] ),
    .B2(_00422_),
    .X(_04747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07228_ (.A(_04747_),
    .Y(_04748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07229_ (.A(\design_top.core0.SIMM[18] ),
    .Y(_00459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07230_ (.A(_00458_),
    .Y(_04749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07231_ (.A(_04749_),
    .X(_04750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07232_ (.A(\design_top.core0.SIMM[18] ),
    .X(_04751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07233_ (.A1(_00459_),
    .A2(_04750_),
    .B1(_04751_),
    .B2(_00458_),
    .X(_04752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07234_ (.A(\design_top.core0.SIMM[19] ),
    .X(_04753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _07235_ (.A(\design_top.core0.SIMM[19] ),
    .B(_00452_),
    .Y(_04754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _07236_ (.A1(_04753_),
    .A2(_00452_),
    .B1(_04754_),
    .Y(_04755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07237_ (.A(\design_top.core0.SIMM[17] ),
    .Y(_00465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07238_ (.A(_04677_),
    .Y(_04756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07239_ (.A1(\design_top.core0.SIMM[17] ),
    .A2(_04677_),
    .B1(_00465_),
    .B2(_04756_),
    .X(_04757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07240_ (.A(\design_top.core0.SIMM[16] ),
    .Y(_00471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07241_ (.A(_00470_),
    .Y(_04758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07242_ (.A1(_00471_),
    .A2(_04758_),
    .B1(\design_top.core0.SIMM[16] ),
    .B2(_00470_),
    .X(_04759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and4_2 _07243_ (.A(_04752_),
    .B(_04755_),
    .C(_04757_),
    .D(_04759_),
    .X(_04760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07244_ (.A(\design_top.core0.SIMM[21] ),
    .Y(_00441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07245_ (.A(_04696_),
    .Y(_04761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07246_ (.A1(\design_top.core0.SIMM[21] ),
    .A2(_04696_),
    .B1(_00441_),
    .B2(_04761_),
    .X(_04762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07247_ (.A(_04762_),
    .Y(_04763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07248_ (.A(\design_top.core0.SIMM[20] ),
    .Y(_00447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07249_ (.A(_00446_),
    .Y(_04764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07250_ (.A(\design_top.core0.SIMM[20] ),
    .X(_04765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07251_ (.A1(_00447_),
    .A2(_04764_),
    .B1(_04765_),
    .B2(_00446_),
    .X(_04766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07252_ (.A(_04766_),
    .Y(_04767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07253_ (.A(\design_top.core0.SIMM[22] ),
    .Y(_00435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07254_ (.A(_00434_),
    .Y(_04768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07255_ (.A(\design_top.core0.SIMM[22] ),
    .X(_04769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _07256_ (.A1(_00435_),
    .A2(_04768_),
    .B1(_04769_),
    .B2(_04688_),
    .X(_04770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07257_ (.A(\design_top.core0.SIMM[23] ),
    .Y(_00429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07258_ (.A(_00428_),
    .Y(_04771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _07259_ (.A1(_00429_),
    .A2(_04771_),
    .B1(\design_top.core0.SIMM[23] ),
    .B2(_00428_),
    .X(_04772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor4_2 _07260_ (.A(_04763_),
    .B(_04767_),
    .C(_04770_),
    .D(_04772_),
    .Y(_04773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07261_ (.A(\design_top.core0.SIMM[14] ),
    .Y(_04774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07262_ (.A(_00482_),
    .Y(_04775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07263_ (.A(\design_top.core0.SIMM[14] ),
    .X(_04776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07264_ (.A1(_04774_),
    .A2(_04775_),
    .B1(_04776_),
    .B2(_00482_),
    .X(_04777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07265_ (.A(_04777_),
    .Y(_04778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _07266_ (.A(\design_top.core0.SIMM[15] ),
    .B(_00476_),
    .Y(_04779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _07267_ (.A1(\design_top.core0.SIMM[15] ),
    .A2(_00476_),
    .B1(_04779_),
    .Y(_04780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07268_ (.A(_04780_),
    .Y(_04781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07269_ (.A(\design_top.core0.SIMM[13] ),
    .Y(_00489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07270_ (.A(_00488_),
    .Y(_04782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07271_ (.A1(_00489_),
    .A2(_04782_),
    .B1(\design_top.core0.SIMM[13] ),
    .B2(_04655_),
    .X(_04783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07272_ (.A(_04783_),
    .Y(_04784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07273_ (.A(\design_top.core0.SIMM[12] ),
    .Y(_00495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07274_ (.A(_00494_),
    .Y(_04785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07275_ (.A(\design_top.core0.SIMM[12] ),
    .X(_04786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07276_ (.A1(_00495_),
    .A2(_04785_),
    .B1(_04786_),
    .B2(_00494_),
    .X(_04787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07277_ (.A(_04787_),
    .Y(_04788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07278_ (.A(_04778_),
    .B(_04781_),
    .C(_04784_),
    .D(_04788_),
    .X(_04789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07279_ (.A(\design_top.core0.SIMM[10] ),
    .Y(_04790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07280_ (.A(_00506_),
    .Y(_04791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07281_ (.A1(_04790_),
    .A2(_04791_),
    .B1(\design_top.core0.SIMM[10] ),
    .B2(_00506_),
    .X(_04792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07282_ (.A(_04792_),
    .Y(_04793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _07283_ (.A(\design_top.core0.SIMM[11] ),
    .B(_00500_),
    .Y(_04794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _07284_ (.A1(\design_top.core0.SIMM[11] ),
    .A2(_00500_),
    .B1(_04794_),
    .Y(_04795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07285_ (.A(_04795_),
    .Y(_04796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _07286_ (.A1(\design_top.core0.SIMM[9] ),
    .A2(_00512_),
    .B1(\design_top.core0.SIMM[8] ),
    .B2(_00518_),
    .X(_04797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07287_ (.A1(\design_top.core0.SIMM[9] ),
    .A2(_00512_),
    .B1(_04797_),
    .Y(_04798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07288_ (.A(_04790_),
    .X(_00507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07289_ (.A(\design_top.core0.SIMM[11] ),
    .X(_04799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07290_ (.A(_04799_),
    .Y(_00501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07291_ (.A(_00500_),
    .Y(_01383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _07292_ (.A1(_00507_),
    .A2(_04791_),
    .A3(_04794_),
    .B1(_00501_),
    .B2(_01383_),
    .X(_04800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _07293_ (.A1(_04793_),
    .A2(_04796_),
    .A3(_04798_),
    .B1(_04800_),
    .X(_04801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07294_ (.A(\design_top.core0.SIMM[4] ),
    .Y(_00347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07295_ (.A(_04644_),
    .Y(_04802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _07296_ (.A1(\design_top.core0.SIMM[4] ),
    .A2(_04644_),
    .B1(_00347_),
    .B2(_04802_),
    .X(_04803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07297_ (.A(\design_top.core0.SIMM[5] ),
    .Y(_00354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07298_ (.A(_00359_),
    .Y(_04804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _07299_ (.A1(\design_top.core0.SIMM[5] ),
    .A2(_04642_),
    .B1(_00354_),
    .B2(_04804_),
    .X(_04805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07300_ (.A(\design_top.core0.SIMM[7] ),
    .Y(_00525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07301_ (.A(_00524_),
    .Y(_04806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _07302_ (.A1(\design_top.core0.SIMM[7] ),
    .A2(_00524_),
    .B1(_00525_),
    .B2(_04806_),
    .X(_04807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07303_ (.A(\design_top.core0.SIMM[6] ),
    .Y(_00531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07304_ (.A(_00530_),
    .Y(_04808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _07305_ (.A1(\design_top.core0.SIMM[6] ),
    .A2(_00530_),
    .B1(_00531_),
    .B2(_04808_),
    .X(_04809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07306_ (.A(_04807_),
    .B(_04809_),
    .X(_04810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07307_ (.A(\design_top.core0.SIMM[3] ),
    .X(_04811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _07308_ (.A(\design_top.core0.SIMM[3] ),
    .B(_00342_),
    .Y(_04812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _07309_ (.A1(_04811_),
    .A2(_00342_),
    .B1(_04812_),
    .X(_04813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07310_ (.A(\design_top.core0.SIMM[2] ),
    .Y(_00310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07311_ (.A(\design_top.core0.SIMM[2] ),
    .X(_04814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07312_ (.A1(_00310_),
    .A2(_04662_),
    .B1(_04814_),
    .B2(_00317_),
    .X(_04815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07313_ (.A(_04815_),
    .Y(_04816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07314_ (.A(\design_top.core0.SIMM[1] ),
    .X(_04817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07315_ (.A(\design_top.core0.SIMM[0] ),
    .Y(_04818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07316_ (.A(_00333_),
    .Y(_04819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _07317_ (.A(_04818_),
    .B(_04819_),
    .Y(_04820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07318_ (.A(\design_top.core0.SIMM[1] ),
    .Y(_00325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07319_ (.A(_00324_),
    .Y(_04821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07320_ (.A1(_00325_),
    .A2(_04821_),
    .B1(\design_top.core0.SIMM[1] ),
    .B2(_00324_),
    .X(_04822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _07321_ (.A1(_04817_),
    .A2(_00324_),
    .B1(_04820_),
    .B2(_04822_),
    .X(_04823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07322_ (.A(_04823_),
    .Y(_04824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07323_ (.A(\design_top.core0.SIMM[3] ),
    .Y(_00335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07324_ (.A(_00342_),
    .Y(_04825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _07325_ (.A1(_00310_),
    .A2(_04662_),
    .A3(_04812_),
    .B1(_00335_),
    .B2(_04825_),
    .X(_04826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _07326_ (.A1(_04813_),
    .A2(_04816_),
    .A3(_04824_),
    .B1(_04826_),
    .X(_04827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _07327_ (.A1(\design_top.core0.SIMM[4] ),
    .A2(_00352_),
    .B1(\design_top.core0.SIMM[5] ),
    .B2(_00359_),
    .X(_04828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07328_ (.A1(\design_top.core0.SIMM[5] ),
    .A2(_04642_),
    .B1(_04828_),
    .Y(_04829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _07329_ (.A1(_00525_),
    .A2(_04806_),
    .B1(_00531_),
    .C1(_04808_),
    .X(_04830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _07330_ (.A1(_00525_),
    .A2(_04806_),
    .B1(_04810_),
    .B2(_04829_),
    .C1(_04830_),
    .X(_04831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o41a_2 _07331_ (.A1(_04803_),
    .A2(_04805_),
    .A3(_04810_),
    .A4(_04827_),
    .B1(_04831_),
    .X(_04832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07332_ (.A(\design_top.core0.SIMM[9] ),
    .Y(_00513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07333_ (.A(_00512_),
    .Y(_01385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07334_ (.A1(_00513_),
    .A2(_01385_),
    .B1(\design_top.core0.SIMM[9] ),
    .B2(_00512_),
    .X(_04833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07335_ (.A(_04833_),
    .Y(_04834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07336_ (.A(\design_top.core0.SIMM[8] ),
    .Y(_00519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07337_ (.A(_00518_),
    .Y(_00775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07338_ (.A1(_00519_),
    .A2(_00775_),
    .B1(\design_top.core0.SIMM[8] ),
    .B2(_00518_),
    .X(_04835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07339_ (.A(_04835_),
    .Y(_04836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07340_ (.A(_04793_),
    .B(_04796_),
    .C(_04834_),
    .D(_04836_),
    .X(_04837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07341_ (.A(_04789_),
    .B(_04837_),
    .X(_04838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _07342_ (.A1(\design_top.core0.SIMM[13] ),
    .A2(_04655_),
    .B1(_04786_),
    .B2(_04658_),
    .X(_04839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _07343_ (.A1(\design_top.core0.SIMM[13] ),
    .A2(_04655_),
    .B1(_04839_),
    .Y(_04840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07344_ (.A(_04774_),
    .X(_00483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07345_ (.A(\design_top.core0.SIMM[15] ),
    .X(_04841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07346_ (.A(_04841_),
    .Y(_00477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07347_ (.A(_04665_),
    .Y(_04842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _07348_ (.A1(_00483_),
    .A2(_04775_),
    .A3(_04779_),
    .B1(_00477_),
    .B2(_04842_),
    .X(_04843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _07349_ (.A1(_04778_),
    .A2(_04781_),
    .A3(_04840_),
    .B1(_04843_),
    .X(_04844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221ai_2 _07350_ (.A1(_04789_),
    .A2(_04801_),
    .B1(_04832_),
    .B2(_04838_),
    .C1(_04844_),
    .Y(_04845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07351_ (.A(\design_top.core0.SIMM[23] ),
    .X(_04846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _07352_ (.A1(\design_top.core0.SIMM[17] ),
    .A2(_00464_),
    .B1(\design_top.core0.SIMM[16] ),
    .B2(_00470_),
    .X(_04847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _07353_ (.A1(\design_top.core0.SIMM[17] ),
    .A2(_04677_),
    .B1(_04847_),
    .X(_04848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07354_ (.A(\design_top.core0.SIMM[19] ),
    .Y(_00453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07355_ (.A(_00452_),
    .Y(_04849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _07356_ (.A1(_00459_),
    .A2(_04749_),
    .A3(_04754_),
    .B1(_00453_),
    .B2(_04849_),
    .X(_04850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07357_ (.A(_04850_),
    .Y(_04851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _07358_ (.A1(_04752_),
    .A2(_04755_),
    .A3(_04848_),
    .B1(_04851_),
    .X(_04852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _07359_ (.A1(\design_top.core0.SIMM[21] ),
    .A2(_00440_),
    .B1(_04765_),
    .B2(_00446_),
    .X(_04853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _07360_ (.A1(\design_top.core0.SIMM[21] ),
    .A2(_04696_),
    .B1(_04853_),
    .X(_04854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _07361_ (.A1(_04762_),
    .A2(_04766_),
    .A3(_04852_),
    .B1(_04854_),
    .X(_04855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _07362_ (.A1(\design_top.core0.SIMM[22] ),
    .A2(_00434_),
    .B1(_04855_),
    .X(_04856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _07363_ (.A1(\design_top.core0.SIMM[23] ),
    .A2(_00428_),
    .B1(\design_top.core0.SIMM[22] ),
    .B2(_04688_),
    .X(_04857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07364_ (.A1(_04846_),
    .A2(_00428_),
    .B1(_04856_),
    .B2(_04857_),
    .X(_04858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _07365_ (.A1(_04760_),
    .A2(_04773_),
    .A3(_04845_),
    .B1(_04858_),
    .X(_04859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07366_ (.A(_04859_),
    .Y(_04860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07367_ (.A(_04745_),
    .B(_04748_),
    .C(_04739_),
    .D(_04860_),
    .X(_04861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2111a_2 _07368_ (.A1(_00405_),
    .A2(_04733_),
    .B1(_04736_),
    .C1(_04742_),
    .D1(_04861_),
    .X(_04862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07369_ (.A(\design_top.core0.SIMM[29] ),
    .Y(_00393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07370_ (.A(_00392_),
    .Y(_04863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _07371_ (.A1(_00399_),
    .A2(_04728_),
    .A3(_04725_),
    .B1(_00393_),
    .B2(_04863_),
    .X(_04864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _07372_ (.A1(_04727_),
    .A2(_04731_),
    .A3(_04862_),
    .B1(_04864_),
    .X(_04865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _07373_ (.A1(_00387_),
    .A2(_04722_),
    .B1(_04723_),
    .B2(_04865_),
    .Y(_04866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07374_ (.A(_04701_),
    .X(_04867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07375_ (.A(\design_top.core0.SIMM[31] ),
    .Y(_01360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _07376_ (.A1(\design_top.core0.SIMM[31] ),
    .A2(_04867_),
    .B1(_01360_),
    .B2(_00381_),
    .X(_04868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07377_ (.A1_N(_04866_),
    .A2_N(_04868_),
    .B1(_04866_),
    .B2(_04868_),
    .X(\design_top.DADDR[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _07378_ (.A(_04619_),
    .B(_04720_),
    .C(\design_top.DADDR[31] ),
    .X(_04869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07379_ (.A(_00553_),
    .B(_04869_),
    .X(_04870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07380_ (.A(_04870_),
    .X(_04871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07381_ (.A1(_00310_),
    .A2(_04663_),
    .B1(_04824_),
    .B2(_04816_),
    .X(_04872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07382_ (.A1_N(_04813_),
    .A2_N(_04872_),
    .B1(_04813_),
    .B2(_04872_),
    .X(_00343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07383_ (.A(_00343_),
    .Y(\design_top.DADDR[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07384_ (.A1(_04824_),
    .A2(_04816_),
    .B1(_04823_),
    .B2(_04815_),
    .X(\design_top.DADDR[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07385_ (.A(\design_top.DADDR[2] ),
    .Y(_00334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07386_ (.A(\design_top.DADDR[3] ),
    .B(_00334_),
    .X(_04873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07387_ (.A1_N(_04827_),
    .A2_N(_04803_),
    .B1(_04827_),
    .B2(_04803_),
    .X(_00353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07388_ (.A(_00353_),
    .Y(_00543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _07389_ (.A1(_00347_),
    .A2(_04802_),
    .B1(_04827_),
    .B2(_04803_),
    .X(_04874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07390_ (.A1_N(_04805_),
    .A2_N(_04874_),
    .B1(_04805_),
    .B2(_04874_),
    .X(_00360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07391_ (.A(_00543_),
    .B(_00360_),
    .X(_04875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07392_ (.A(_04873_),
    .B(_04875_),
    .X(_04876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07393_ (.A(_04871_),
    .B(_04876_),
    .X(_04877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07394_ (.A(_04877_),
    .X(_04878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07395_ (.A(wbs_adr_i[0]),
    .X(_04879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07396_ (.A(wbs_adr_i[1]),
    .Y(_04880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07397_ (.A(_04880_),
    .X(_04881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07398_ (.A(\design_top.XRES ),
    .Y(_04882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07399_ (.A(_04882_),
    .X(_04883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07400_ (.A(wbs_we_i),
    .Y(_04884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _07401_ (.A(_04883_),
    .B(_04884_),
    .C_N(wbs_sel_i[1]),
    .X(_04885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _07402_ (.A(_04879_),
    .B(_04881_),
    .C(_04885_),
    .Y(_04886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07403_ (.A(_04886_),
    .B_N(_04877_),
    .Y(_04887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07404_ (.A(_04887_),
    .X(_04888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07405_ (.A1_N(_04719_),
    .A2_N(_04878_),
    .B1(\design_top.MEM[9][31] ),
    .B2(_04888_),
    .X(_04435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07406_ (.A(\design_top.DATAO[30] ),
    .Y(_04889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07407_ (.A(_04889_),
    .X(_04890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07408_ (.A1_N(_04890_),
    .A2_N(_04878_),
    .B1(\design_top.MEM[9][30] ),
    .B2(_04888_),
    .X(_04434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07409_ (.A(\design_top.DATAO[29] ),
    .Y(_04891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07410_ (.A(_04891_),
    .X(_04892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07411_ (.A1_N(_04892_),
    .A2_N(_04878_),
    .B1(\design_top.MEM[9][29] ),
    .B2(_04888_),
    .X(_04433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07412_ (.A(\design_top.DATAO[28] ),
    .Y(_04893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07413_ (.A(_04893_),
    .X(_04894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07414_ (.A1_N(_04894_),
    .A2_N(_04878_),
    .B1(\design_top.MEM[9][28] ),
    .B2(_04888_),
    .X(_04432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07415_ (.A(\design_top.DATAO[27] ),
    .Y(_04895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07416_ (.A(_04895_),
    .X(_04896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07417_ (.A1_N(_04896_),
    .A2_N(_04878_),
    .B1(\design_top.MEM[9][27] ),
    .B2(_04888_),
    .X(_04431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07418_ (.A(\design_top.DATAO[26] ),
    .Y(_04897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07419_ (.A(_04897_),
    .X(_04898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07420_ (.A1_N(_04898_),
    .A2_N(_04877_),
    .B1(\design_top.MEM[9][26] ),
    .B2(_04887_),
    .X(_04430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07421_ (.A(\design_top.DATAO[25] ),
    .Y(_04899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07422_ (.A(_04899_),
    .X(_04900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07423_ (.A1_N(_04900_),
    .A2_N(_04877_),
    .B1(\design_top.MEM[9][25] ),
    .B2(_04887_),
    .X(_04429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07424_ (.A(\design_top.DATAO[24] ),
    .Y(_04901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07425_ (.A(_04901_),
    .X(_04902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07426_ (.A1_N(_04902_),
    .A2_N(_04877_),
    .B1(\design_top.MEM[9][24] ),
    .B2(_04887_),
    .X(_04428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07427_ (.A(\design_top.DATAO[15] ),
    .Y(_04903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07428_ (.A(_04903_),
    .X(_04904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07429_ (.A(_00353_),
    .B(_00360_),
    .X(_04905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07430_ (.A(_00343_),
    .B(\design_top.DADDR[2] ),
    .X(_04906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07431_ (.A(_04905_),
    .B(_04906_),
    .X(_04907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07432_ (.A(_00547_),
    .B(_04869_),
    .X(_04908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07433_ (.A(_04908_),
    .X(_04909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07434_ (.A(_04907_),
    .B(_04909_),
    .X(_04910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07435_ (.A(_04910_),
    .X(_04911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07436_ (.A(wbs_adr_i[0]),
    .Y(_04912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07437_ (.A(_04912_),
    .X(_04913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _07438_ (.A(_04882_),
    .B(_04884_),
    .C_N(wbs_sel_i[2]),
    .X(_04914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _07439_ (.A(_04913_),
    .B(_04881_),
    .C(_04914_),
    .Y(_04915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07440_ (.A(_04915_),
    .B_N(_04910_),
    .Y(_04916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07441_ (.A(_04916_),
    .X(_04917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07442_ (.A1_N(_04904_),
    .A2_N(_04911_),
    .B1(\design_top.MEM[14][15] ),
    .B2(_04917_),
    .X(_04427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07443_ (.A(\design_top.DATAO[14] ),
    .Y(_04918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07444_ (.A(_04918_),
    .X(_04919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07445_ (.A1_N(_04919_),
    .A2_N(_04911_),
    .B1(\design_top.MEM[14][14] ),
    .B2(_04917_),
    .X(_04426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07446_ (.A(\design_top.DATAO[13] ),
    .Y(_04920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07447_ (.A(_04920_),
    .X(_04921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07448_ (.A1_N(_04921_),
    .A2_N(_04911_),
    .B1(\design_top.MEM[14][13] ),
    .B2(_04917_),
    .X(_04425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07449_ (.A(\design_top.DATAO[12] ),
    .Y(_04922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07450_ (.A(_04922_),
    .X(_04923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07451_ (.A1_N(_04923_),
    .A2_N(_04911_),
    .B1(\design_top.MEM[14][12] ),
    .B2(_04917_),
    .X(_04424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07452_ (.A(\design_top.DATAO[11] ),
    .Y(_04924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07453_ (.A(_04924_),
    .X(_04925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07454_ (.A1_N(_04925_),
    .A2_N(_04911_),
    .B1(\design_top.MEM[14][11] ),
    .B2(_04917_),
    .X(_04423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07455_ (.A(\design_top.DATAO[10] ),
    .Y(_04926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07456_ (.A(_04926_),
    .X(_04927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07457_ (.A1_N(_04927_),
    .A2_N(_04910_),
    .B1(\design_top.MEM[14][10] ),
    .B2(_04916_),
    .X(_04422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07458_ (.A(\design_top.DATAO[9] ),
    .Y(_04928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07459_ (.A(_04928_),
    .X(_04929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07460_ (.A1_N(_04929_),
    .A2_N(_04910_),
    .B1(\design_top.MEM[14][9] ),
    .B2(_04916_),
    .X(_04421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07461_ (.A(\design_top.DATAO[8] ),
    .Y(_04930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07462_ (.A(_04930_),
    .X(_04931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07463_ (.A1_N(_04931_),
    .A2_N(_04910_),
    .B1(\design_top.MEM[14][8] ),
    .B2(_04916_),
    .X(_04420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07464_ (.A(_04871_),
    .B(_04907_),
    .X(_04932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07465_ (.A(_04932_),
    .X(_04933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07466_ (.A(_04915_),
    .B_N(_04932_),
    .Y(_04934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07467_ (.A(_04934_),
    .X(_04935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07468_ (.A1_N(_04719_),
    .A2_N(_04933_),
    .B1(\design_top.MEM[14][31] ),
    .B2(_04935_),
    .X(_04419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07469_ (.A1_N(_04890_),
    .A2_N(_04933_),
    .B1(\design_top.MEM[14][30] ),
    .B2(_04935_),
    .X(_04418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07470_ (.A1_N(_04892_),
    .A2_N(_04933_),
    .B1(\design_top.MEM[14][29] ),
    .B2(_04935_),
    .X(_04417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07471_ (.A1_N(_04894_),
    .A2_N(_04933_),
    .B1(\design_top.MEM[14][28] ),
    .B2(_04935_),
    .X(_04416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07472_ (.A1_N(_04896_),
    .A2_N(_04933_),
    .B1(\design_top.MEM[14][27] ),
    .B2(_04935_),
    .X(_04415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07473_ (.A1_N(_04898_),
    .A2_N(_04932_),
    .B1(\design_top.MEM[14][26] ),
    .B2(_04934_),
    .X(_04414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07474_ (.A1_N(_04900_),
    .A2_N(_04932_),
    .B1(\design_top.MEM[14][25] ),
    .B2(_04934_),
    .X(_04413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07475_ (.A1_N(_04902_),
    .A2_N(_04932_),
    .B1(\design_top.MEM[14][24] ),
    .B2(_04934_),
    .X(_04412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07476_ (.A(\design_top.DATAO[23] ),
    .Y(_04936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07477_ (.A(_04936_),
    .X(_04937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07478_ (.A(_00542_),
    .B(_04869_),
    .X(_04938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07479_ (.A(_04938_),
    .X(_04939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07480_ (.A(_04907_),
    .B(_04939_),
    .X(_04940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07481_ (.A(_04940_),
    .X(_04941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07482_ (.A(_04915_),
    .B_N(_04940_),
    .Y(_04942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07483_ (.A(_04942_),
    .X(_04943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07484_ (.A1_N(_04937_),
    .A2_N(_04941_),
    .B1(\design_top.MEM[14][23] ),
    .B2(_04943_),
    .X(_04411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07485_ (.A(\design_top.DATAO[22] ),
    .Y(_04944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07486_ (.A(_04944_),
    .X(_04945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07487_ (.A1_N(_04945_),
    .A2_N(_04941_),
    .B1(\design_top.MEM[14][22] ),
    .B2(_04943_),
    .X(_04410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07488_ (.A(\design_top.DATAO[21] ),
    .Y(_04946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07489_ (.A(_04946_),
    .X(_04947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07490_ (.A1_N(_04947_),
    .A2_N(_04941_),
    .B1(\design_top.MEM[14][21] ),
    .B2(_04943_),
    .X(_04409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07491_ (.A(\design_top.DATAO[20] ),
    .Y(_04948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07492_ (.A(_04948_),
    .X(_04949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07493_ (.A1_N(_04949_),
    .A2_N(_04941_),
    .B1(\design_top.MEM[14][20] ),
    .B2(_04943_),
    .X(_04408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07494_ (.A(\design_top.DATAO[19] ),
    .Y(_04950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07495_ (.A(_04950_),
    .X(_04951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07496_ (.A1_N(_04951_),
    .A2_N(_04941_),
    .B1(\design_top.MEM[14][19] ),
    .B2(_04943_),
    .X(_04407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07497_ (.A(\design_top.DATAO[18] ),
    .Y(_04952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07498_ (.A(_04952_),
    .X(_04953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07499_ (.A1_N(_04953_),
    .A2_N(_04940_),
    .B1(\design_top.MEM[14][18] ),
    .B2(_04942_),
    .X(_04406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07500_ (.A(\design_top.DATAO[17] ),
    .Y(_04954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07501_ (.A(_04954_),
    .X(_04955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07502_ (.A1_N(_04955_),
    .A2_N(_04940_),
    .B1(\design_top.MEM[14][17] ),
    .B2(_04942_),
    .X(_04405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07503_ (.A(\design_top.DATAO[16] ),
    .Y(_04956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07504_ (.A(_04956_),
    .X(_04957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07505_ (.A1_N(_04957_),
    .A2_N(_04940_),
    .B1(\design_top.MEM[14][16] ),
    .B2(_04942_),
    .X(_04404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07506_ (.A(\design_top.DADDR[3] ),
    .B(\design_top.DADDR[2] ),
    .X(_04958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07507_ (.A(_00360_),
    .Y(_02415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07508_ (.A(_00543_),
    .B(_02415_),
    .X(_04959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07509_ (.A(_04958_),
    .B(_04959_),
    .X(_04960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07510_ (.A(_04871_),
    .B(_04960_),
    .X(_04961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07511_ (.A(_04961_),
    .X(_04962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07512_ (.A(wbs_adr_i[1]),
    .X(_04963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _07513_ (.A(_04882_),
    .B(_04884_),
    .C_N(wbs_sel_i[0]),
    .X(_04964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _07514_ (.A(_04879_),
    .B(_04963_),
    .C(_04964_),
    .Y(_04965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07515_ (.A(_04965_),
    .B_N(_04961_),
    .Y(_04966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07516_ (.A(_04966_),
    .X(_04967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07517_ (.A1_N(_04719_),
    .A2_N(_04962_),
    .B1(\design_top.MEM[0][31] ),
    .B2(_04967_),
    .X(_04403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07518_ (.A1_N(_04890_),
    .A2_N(_04962_),
    .B1(\design_top.MEM[0][30] ),
    .B2(_04967_),
    .X(_04402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07519_ (.A1_N(_04892_),
    .A2_N(_04962_),
    .B1(\design_top.MEM[0][29] ),
    .B2(_04967_),
    .X(_04401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07520_ (.A1_N(_04894_),
    .A2_N(_04962_),
    .B1(\design_top.MEM[0][28] ),
    .B2(_04967_),
    .X(_04400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07521_ (.A1_N(_04896_),
    .A2_N(_04962_),
    .B1(\design_top.MEM[0][27] ),
    .B2(_04967_),
    .X(_04399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07522_ (.A1_N(_04898_),
    .A2_N(_04961_),
    .B1(\design_top.MEM[0][26] ),
    .B2(_04966_),
    .X(_04398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07523_ (.A1_N(_04900_),
    .A2_N(_04961_),
    .B1(\design_top.MEM[0][25] ),
    .B2(_04966_),
    .X(_04397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07524_ (.A1_N(_04902_),
    .A2_N(_04961_),
    .B1(\design_top.MEM[0][24] ),
    .B2(_04966_),
    .X(_04396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07525_ (.A(_04939_),
    .B(_04960_),
    .X(_04968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07526_ (.A(_04968_),
    .X(_04969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07527_ (.A(_04965_),
    .B_N(_04968_),
    .Y(_04970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07528_ (.A(_04970_),
    .X(_04971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07529_ (.A1_N(_04937_),
    .A2_N(_04969_),
    .B1(\design_top.MEM[0][23] ),
    .B2(_04971_),
    .X(_04395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07530_ (.A1_N(_04945_),
    .A2_N(_04969_),
    .B1(\design_top.MEM[0][22] ),
    .B2(_04971_),
    .X(_04394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07531_ (.A1_N(_04947_),
    .A2_N(_04969_),
    .B1(\design_top.MEM[0][21] ),
    .B2(_04971_),
    .X(_04393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07532_ (.A1_N(_04949_),
    .A2_N(_04969_),
    .B1(\design_top.MEM[0][20] ),
    .B2(_04971_),
    .X(_04392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07533_ (.A1_N(_04951_),
    .A2_N(_04969_),
    .B1(\design_top.MEM[0][19] ),
    .B2(_04971_),
    .X(_04391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07534_ (.A1_N(_04953_),
    .A2_N(_04968_),
    .B1(\design_top.MEM[0][18] ),
    .B2(_04970_),
    .X(_04390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07535_ (.A1_N(_04955_),
    .A2_N(_04968_),
    .B1(\design_top.MEM[0][17] ),
    .B2(_04970_),
    .X(_04389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07536_ (.A1_N(_04957_),
    .A2_N(_04968_),
    .B1(\design_top.MEM[0][16] ),
    .B2(_04970_),
    .X(_04388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07537_ (.A(_04909_),
    .B(_04960_),
    .X(_04972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07538_ (.A(_04972_),
    .X(_04973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07539_ (.A(_04965_),
    .B_N(_04972_),
    .Y(_04974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07540_ (.A(_04974_),
    .X(_04975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07541_ (.A1_N(_04904_),
    .A2_N(_04973_),
    .B1(\design_top.MEM[0][15] ),
    .B2(_04975_),
    .X(_04387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07542_ (.A1_N(_04919_),
    .A2_N(_04973_),
    .B1(\design_top.MEM[0][14] ),
    .B2(_04975_),
    .X(_04386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07543_ (.A1_N(_04921_),
    .A2_N(_04973_),
    .B1(\design_top.MEM[0][13] ),
    .B2(_04975_),
    .X(_04385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07544_ (.A1_N(_04923_),
    .A2_N(_04973_),
    .B1(\design_top.MEM[0][12] ),
    .B2(_04975_),
    .X(_04384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07545_ (.A1_N(_04925_),
    .A2_N(_04973_),
    .B1(\design_top.MEM[0][11] ),
    .B2(_04975_),
    .X(_04383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07546_ (.A1_N(_04927_),
    .A2_N(_04972_),
    .B1(\design_top.MEM[0][10] ),
    .B2(_04974_),
    .X(_04382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07547_ (.A1_N(_04929_),
    .A2_N(_04972_),
    .B1(\design_top.MEM[0][9] ),
    .B2(_04974_),
    .X(_04381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07548_ (.A1_N(_04931_),
    .A2_N(_04972_),
    .B1(\design_top.MEM[0][8] ),
    .B2(_04974_),
    .X(_04380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07549_ (.A(_04875_),
    .B(_04906_),
    .X(_04976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07550_ (.A(_04909_),
    .B(_04976_),
    .X(_04977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07551_ (.A(_04977_),
    .X(_04978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _07552_ (.A(_04879_),
    .B(_04881_),
    .C(_04914_),
    .Y(_04979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07553_ (.A(_04979_),
    .B_N(_04977_),
    .Y(_04980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07554_ (.A(_04980_),
    .X(_04981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07555_ (.A1_N(_04904_),
    .A2_N(_04978_),
    .B1(\design_top.MEM[10][15] ),
    .B2(_04981_),
    .X(_04379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07556_ (.A1_N(_04919_),
    .A2_N(_04978_),
    .B1(\design_top.MEM[10][14] ),
    .B2(_04981_),
    .X(_04378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07557_ (.A1_N(_04921_),
    .A2_N(_04978_),
    .B1(\design_top.MEM[10][13] ),
    .B2(_04981_),
    .X(_04377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07558_ (.A1_N(_04923_),
    .A2_N(_04978_),
    .B1(\design_top.MEM[10][12] ),
    .B2(_04981_),
    .X(_04376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07559_ (.A1_N(_04925_),
    .A2_N(_04978_),
    .B1(\design_top.MEM[10][11] ),
    .B2(_04981_),
    .X(_04375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07560_ (.A1_N(_04927_),
    .A2_N(_04977_),
    .B1(\design_top.MEM[10][10] ),
    .B2(_04980_),
    .X(_04374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07561_ (.A1_N(_04929_),
    .A2_N(_04977_),
    .B1(\design_top.MEM[10][9] ),
    .B2(_04980_),
    .X(_04373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07562_ (.A1_N(_04931_),
    .A2_N(_04977_),
    .B1(\design_top.MEM[10][8] ),
    .B2(_04980_),
    .X(_04372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07563_ (.A(_04939_),
    .B(_04976_),
    .X(_04982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07564_ (.A(_04982_),
    .X(_04983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07565_ (.A(_04979_),
    .B_N(_04982_),
    .Y(_04984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07566_ (.A(_04984_),
    .X(_04985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07567_ (.A1_N(_04937_),
    .A2_N(_04983_),
    .B1(\design_top.MEM[10][23] ),
    .B2(_04985_),
    .X(_04371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07568_ (.A1_N(_04945_),
    .A2_N(_04983_),
    .B1(\design_top.MEM[10][22] ),
    .B2(_04985_),
    .X(_04370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07569_ (.A1_N(_04947_),
    .A2_N(_04983_),
    .B1(\design_top.MEM[10][21] ),
    .B2(_04985_),
    .X(_04369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07570_ (.A1_N(_04949_),
    .A2_N(_04983_),
    .B1(\design_top.MEM[10][20] ),
    .B2(_04985_),
    .X(_04368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07571_ (.A1_N(_04951_),
    .A2_N(_04983_),
    .B1(\design_top.MEM[10][19] ),
    .B2(_04985_),
    .X(_04367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07572_ (.A1_N(_04953_),
    .A2_N(_04982_),
    .B1(\design_top.MEM[10][18] ),
    .B2(_04984_),
    .X(_04366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07573_ (.A1_N(_04955_),
    .A2_N(_04982_),
    .B1(\design_top.MEM[10][17] ),
    .B2(_04984_),
    .X(_04365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07574_ (.A1_N(_04957_),
    .A2_N(_04982_),
    .B1(\design_top.MEM[10][16] ),
    .B2(_04984_),
    .X(_04364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07575_ (.A(_04871_),
    .B(_04976_),
    .X(_04986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07576_ (.A(_04986_),
    .X(_04987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07577_ (.A(_04979_),
    .B_N(_04986_),
    .Y(_04988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07578_ (.A(_04988_),
    .X(_04989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07579_ (.A1_N(_04719_),
    .A2_N(_04987_),
    .B1(\design_top.MEM[10][31] ),
    .B2(_04989_),
    .X(_04363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07580_ (.A1_N(_04890_),
    .A2_N(_04987_),
    .B1(\design_top.MEM[10][30] ),
    .B2(_04989_),
    .X(_04362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07581_ (.A1_N(_04892_),
    .A2_N(_04987_),
    .B1(\design_top.MEM[10][29] ),
    .B2(_04989_),
    .X(_04361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07582_ (.A1_N(_04894_),
    .A2_N(_04987_),
    .B1(\design_top.MEM[10][28] ),
    .B2(_04989_),
    .X(_04360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07583_ (.A1_N(_04896_),
    .A2_N(_04987_),
    .B1(\design_top.MEM[10][27] ),
    .B2(_04989_),
    .X(_04359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07584_ (.A1_N(_04898_),
    .A2_N(_04986_),
    .B1(\design_top.MEM[10][26] ),
    .B2(_04988_),
    .X(_04358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07585_ (.A1_N(_04900_),
    .A2_N(_04986_),
    .B1(\design_top.MEM[10][25] ),
    .B2(_04988_),
    .X(_04357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07586_ (.A1_N(_04902_),
    .A2_N(_04986_),
    .B1(\design_top.MEM[10][24] ),
    .B2(_04988_),
    .X(_04356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07587_ (.A(_00343_),
    .B(_00334_),
    .X(_04990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07588_ (.A(_04875_),
    .B(_04990_),
    .X(_04991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07589_ (.A(_04939_),
    .B(_04991_),
    .X(_04992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07590_ (.A(_04992_),
    .X(_04993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _07591_ (.A(_04882_),
    .B(_04884_),
    .C_N(wbs_sel_i[3]),
    .X(_04994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _07592_ (.A(_04879_),
    .B(_04881_),
    .C(_04994_),
    .Y(_04995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07593_ (.A(_04995_),
    .B_N(_04992_),
    .Y(_04996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07594_ (.A(_04996_),
    .X(_04997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07595_ (.A1_N(_04937_),
    .A2_N(_04993_),
    .B1(\design_top.MEM[11][23] ),
    .B2(_04997_),
    .X(_04355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07596_ (.A1_N(_04945_),
    .A2_N(_04993_),
    .B1(\design_top.MEM[11][22] ),
    .B2(_04997_),
    .X(_04354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07597_ (.A1_N(_04947_),
    .A2_N(_04993_),
    .B1(\design_top.MEM[11][21] ),
    .B2(_04997_),
    .X(_04353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07598_ (.A1_N(_04949_),
    .A2_N(_04993_),
    .B1(\design_top.MEM[11][20] ),
    .B2(_04997_),
    .X(_04352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07599_ (.A1_N(_04951_),
    .A2_N(_04993_),
    .B1(\design_top.MEM[11][19] ),
    .B2(_04997_),
    .X(_04351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07600_ (.A1_N(_04953_),
    .A2_N(_04992_),
    .B1(\design_top.MEM[11][18] ),
    .B2(_04996_),
    .X(_04350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07601_ (.A1_N(_04955_),
    .A2_N(_04992_),
    .B1(\design_top.MEM[11][17] ),
    .B2(_04996_),
    .X(_04349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07602_ (.A1_N(_04957_),
    .A2_N(_04992_),
    .B1(\design_top.MEM[11][16] ),
    .B2(_04996_),
    .X(_04348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07603_ (.A(_04871_),
    .B(_04991_),
    .X(_04998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07604_ (.A(_04998_),
    .X(_04999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07605_ (.A(_04995_),
    .B_N(_04998_),
    .Y(_05000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07606_ (.A(_05000_),
    .X(_05001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07607_ (.A1_N(_04719_),
    .A2_N(_04999_),
    .B1(\design_top.MEM[11][31] ),
    .B2(_05001_),
    .X(_04347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07608_ (.A1_N(_04890_),
    .A2_N(_04999_),
    .B1(\design_top.MEM[11][30] ),
    .B2(_05001_),
    .X(_04346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07609_ (.A1_N(_04892_),
    .A2_N(_04999_),
    .B1(\design_top.MEM[11][29] ),
    .B2(_05001_),
    .X(_04345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07610_ (.A1_N(_04894_),
    .A2_N(_04999_),
    .B1(\design_top.MEM[11][28] ),
    .B2(_05001_),
    .X(_04344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07611_ (.A1_N(_04896_),
    .A2_N(_04999_),
    .B1(\design_top.MEM[11][27] ),
    .B2(_05001_),
    .X(_04343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07612_ (.A1_N(_04898_),
    .A2_N(_04998_),
    .B1(\design_top.MEM[11][26] ),
    .B2(_05000_),
    .X(_04342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07613_ (.A1_N(_04900_),
    .A2_N(_04998_),
    .B1(\design_top.MEM[11][25] ),
    .B2(_05000_),
    .X(_04341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07614_ (.A1_N(_04902_),
    .A2_N(_04998_),
    .B1(\design_top.MEM[11][24] ),
    .B2(_05000_),
    .X(_04340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07615_ (.A(_04909_),
    .B(_04991_),
    .X(_05002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07616_ (.A(_05002_),
    .X(_05003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07617_ (.A(_04995_),
    .B_N(_05002_),
    .Y(_05004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07618_ (.A(_05004_),
    .X(_05005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07619_ (.A1_N(_04904_),
    .A2_N(_05003_),
    .B1(\design_top.MEM[11][15] ),
    .B2(_05005_),
    .X(_04339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07620_ (.A1_N(_04919_),
    .A2_N(_05003_),
    .B1(\design_top.MEM[11][14] ),
    .B2(_05005_),
    .X(_04338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07621_ (.A1_N(_04921_),
    .A2_N(_05003_),
    .B1(\design_top.MEM[11][13] ),
    .B2(_05005_),
    .X(_04337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07622_ (.A1_N(_04923_),
    .A2_N(_05003_),
    .B1(\design_top.MEM[11][12] ),
    .B2(_05005_),
    .X(_04336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07623_ (.A1_N(_04925_),
    .A2_N(_05003_),
    .B1(\design_top.MEM[11][11] ),
    .B2(_05005_),
    .X(_04335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07624_ (.A1_N(_04927_),
    .A2_N(_05002_),
    .B1(\design_top.MEM[11][10] ),
    .B2(_05004_),
    .X(_04334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07625_ (.A1_N(_04929_),
    .A2_N(_05002_),
    .B1(\design_top.MEM[11][9] ),
    .B2(_05004_),
    .X(_04333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07626_ (.A1_N(_04931_),
    .A2_N(_05002_),
    .B1(\design_top.MEM[11][8] ),
    .B2(_05004_),
    .X(_04332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07627_ (.A(_04908_),
    .X(_05006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07628_ (.A(_04905_),
    .B(_04958_),
    .X(_05007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07629_ (.A(_05006_),
    .B(_05007_),
    .X(_05008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07630_ (.A(_05008_),
    .X(_05009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _07631_ (.A(_04913_),
    .B(_04881_),
    .C(_04964_),
    .Y(_05010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07632_ (.A(_05010_),
    .B_N(_05008_),
    .Y(_05011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07633_ (.A(_05011_),
    .X(_05012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07634_ (.A1_N(_04904_),
    .A2_N(_05009_),
    .B1(\design_top.MEM[12][15] ),
    .B2(_05012_),
    .X(_04331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07635_ (.A1_N(_04919_),
    .A2_N(_05009_),
    .B1(\design_top.MEM[12][14] ),
    .B2(_05012_),
    .X(_04330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07636_ (.A1_N(_04921_),
    .A2_N(_05009_),
    .B1(\design_top.MEM[12][13] ),
    .B2(_05012_),
    .X(_04329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07637_ (.A1_N(_04923_),
    .A2_N(_05009_),
    .B1(\design_top.MEM[12][12] ),
    .B2(_05012_),
    .X(_04328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07638_ (.A1_N(_04925_),
    .A2_N(_05009_),
    .B1(\design_top.MEM[12][11] ),
    .B2(_05012_),
    .X(_04327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07639_ (.A1_N(_04927_),
    .A2_N(_05008_),
    .B1(\design_top.MEM[12][10] ),
    .B2(_05011_),
    .X(_04326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07640_ (.A1_N(_04929_),
    .A2_N(_05008_),
    .B1(\design_top.MEM[12][9] ),
    .B2(_05011_),
    .X(_04325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07641_ (.A1_N(_04931_),
    .A2_N(_05008_),
    .B1(\design_top.MEM[12][8] ),
    .B2(_05011_),
    .X(_04324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07642_ (.A(_04822_),
    .Y(_05013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07643_ (.A(_04818_),
    .X(_00326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _07644_ (.A1(_00326_),
    .A2(_04819_),
    .B1(_04820_),
    .Y(_05014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07645_ (.A(_05014_),
    .Y(_05015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07646_ (.A(_05013_),
    .B(_05015_),
    .X(_05016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07647_ (.A(\design_top.DADDR[31] ),
    .Y(_05017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07648_ (.A(_04720_),
    .B(_05017_),
    .X(_05018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07649_ (.A(_04718_),
    .B(_05016_),
    .C(_04958_),
    .D(_05018_),
    .X(_05019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07650_ (.A(_05019_),
    .Y(_05020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07651_ (.A(\design_top.IRES[7] ),
    .Y(_05021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07652_ (.A(_05021_),
    .X(_05022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07653_ (.A(_05022_),
    .X(_05023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _07654_ (.A1(\design_top.IREQ[7] ),
    .A2(_05019_),
    .B1(\design_top.IACK[7] ),
    .B2(_05020_),
    .C1(_05023_),
    .X(_04323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07655_ (.A(\design_top.IOMUX[3][11] ),
    .B(\design_top.IOMUX[3][10] ),
    .C(\design_top.IOMUX[3][9] ),
    .D(\design_top.IOMUX[3][8] ),
    .X(_05024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07656_ (.A(\design_top.IOMUX[3][15] ),
    .B(\design_top.IOMUX[3][14] ),
    .C(\design_top.IOMUX[3][13] ),
    .D(\design_top.IOMUX[3][12] ),
    .X(_05025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07657_ (.A(\design_top.IOMUX[3][3] ),
    .B(\design_top.IOMUX[3][2] ),
    .C(\design_top.IOMUX[3][1] ),
    .D(\design_top.IOMUX[3][0] ),
    .X(_05026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07658_ (.A(\design_top.IOMUX[3][7] ),
    .B(\design_top.IOMUX[3][6] ),
    .C(\design_top.IOMUX[3][5] ),
    .D(\design_top.IOMUX[3][4] ),
    .X(_05027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07659_ (.A(_05024_),
    .B(_05025_),
    .C(_05026_),
    .D(_05027_),
    .X(_05028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07660_ (.A(\design_top.IOMUX[3][27] ),
    .B(\design_top.IOMUX[3][26] ),
    .C(\design_top.IOMUX[3][25] ),
    .D(\design_top.IOMUX[3][24] ),
    .X(_05029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07661_ (.A(\design_top.IOMUX[3][31] ),
    .B(\design_top.IOMUX[3][30] ),
    .C(\design_top.IOMUX[3][29] ),
    .D(\design_top.IOMUX[3][28] ),
    .X(_05030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07662_ (.A(\design_top.IOMUX[3][19] ),
    .B(\design_top.IOMUX[3][18] ),
    .C(\design_top.IOMUX[3][17] ),
    .D(\design_top.IOMUX[3][16] ),
    .X(_05031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07663_ (.A(\design_top.IOMUX[3][23] ),
    .B(\design_top.IOMUX[3][22] ),
    .C(\design_top.IOMUX[3][21] ),
    .D(\design_top.IOMUX[3][20] ),
    .X(_05032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07664_ (.A(_05029_),
    .B(_05030_),
    .C(_05031_),
    .D(_05032_),
    .X(_05033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _07665_ (.A(_05028_),
    .B(_05033_),
    .Y(_05034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07666_ (.A(\design_top.TIMER[31] ),
    .B(\design_top.TIMER[30] ),
    .X(_05035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07667_ (.A(\design_top.TIMER[19] ),
    .B(\design_top.TIMER[18] ),
    .X(_05036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07668_ (.A(\design_top.TIMER[1] ),
    .B(\design_top.TIMER[0] ),
    .X(_05037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07669_ (.A(\design_top.TIMER[2] ),
    .B(_05037_),
    .X(_05038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07670_ (.A(\design_top.TIMER[3] ),
    .B(_05038_),
    .X(_05039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07671_ (.A(\design_top.TIMER[4] ),
    .B(_05039_),
    .X(_05040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07672_ (.A(\design_top.TIMER[5] ),
    .B(_05040_),
    .X(_05041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07673_ (.A(\design_top.TIMER[6] ),
    .B(_05041_),
    .X(_05042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07674_ (.A(\design_top.TIMER[7] ),
    .B(_05042_),
    .X(_05043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07675_ (.A(\design_top.TIMER[8] ),
    .B(_05043_),
    .X(_05044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07676_ (.A(\design_top.TIMER[9] ),
    .B(_05044_),
    .X(_05045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07677_ (.A(\design_top.TIMER[10] ),
    .B(_05045_),
    .X(_05046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07678_ (.A(\design_top.TIMER[11] ),
    .B(_05046_),
    .X(_05047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07679_ (.A(\design_top.TIMER[12] ),
    .B(_05047_),
    .X(_05048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07680_ (.A(\design_top.TIMER[13] ),
    .B(_05048_),
    .X(_05049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07681_ (.A(\design_top.TIMER[14] ),
    .B(_05049_),
    .X(_05050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07682_ (.A(\design_top.TIMER[15] ),
    .B(_05050_),
    .X(_05051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07683_ (.A(\design_top.TIMER[17] ),
    .B(\design_top.TIMER[16] ),
    .C(_05036_),
    .D(_05051_),
    .X(_05052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _07684_ (.A(\design_top.TIMER[21] ),
    .B(\design_top.TIMER[20] ),
    .C(_05052_),
    .X(_05053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _07685_ (.A(\design_top.TIMER[23] ),
    .B(\design_top.TIMER[22] ),
    .C(_05053_),
    .X(_05054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _07686_ (.A(\design_top.TIMER[25] ),
    .B(\design_top.TIMER[24] ),
    .C(_05054_),
    .X(_05055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07687_ (.A(\design_top.TIMER[26] ),
    .B(_05055_),
    .X(_05056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07688_ (.A(\design_top.TIMER[27] ),
    .B(_05056_),
    .X(_05057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _07689_ (.A(\design_top.TIMER[29] ),
    .B(\design_top.TIMER[28] ),
    .C(_05035_),
    .D(_05057_),
    .X(_05058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07690_ (.A(_05034_),
    .B(_05058_),
    .X(_05059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07691_ (.A(_05059_),
    .Y(_05060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _07692_ (.A(\design_top.IACK[7] ),
    .Y(_05061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07693_ (.A(_05021_),
    .X(_05062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07694_ (.A(_05062_),
    .X(_05063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _07695_ (.A1(\design_top.IREQ[7] ),
    .A2(_05060_),
    .B1(_05061_),
    .B2(_05059_),
    .C1(_05063_),
    .X(_04322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07696_ (.A(_04938_),
    .X(_05064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07697_ (.A(_05064_),
    .B(_05007_),
    .X(_05065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07698_ (.A(_05065_),
    .X(_05066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07699_ (.A(_05010_),
    .B_N(_05065_),
    .Y(_05067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07700_ (.A(_05067_),
    .X(_05068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07701_ (.A1_N(_04937_),
    .A2_N(_05066_),
    .B1(\design_top.MEM[12][23] ),
    .B2(_05068_),
    .X(_04321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07702_ (.A1_N(_04945_),
    .A2_N(_05066_),
    .B1(\design_top.MEM[12][22] ),
    .B2(_05068_),
    .X(_04320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07703_ (.A1_N(_04947_),
    .A2_N(_05066_),
    .B1(\design_top.MEM[12][21] ),
    .B2(_05068_),
    .X(_04319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07704_ (.A1_N(_04949_),
    .A2_N(_05066_),
    .B1(\design_top.MEM[12][20] ),
    .B2(_05068_),
    .X(_04318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07705_ (.A1_N(_04951_),
    .A2_N(_05066_),
    .B1(\design_top.MEM[12][19] ),
    .B2(_05068_),
    .X(_04317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07706_ (.A1_N(_04953_),
    .A2_N(_05065_),
    .B1(\design_top.MEM[12][18] ),
    .B2(_05067_),
    .X(_04316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07707_ (.A1_N(_04955_),
    .A2_N(_05065_),
    .B1(\design_top.MEM[12][17] ),
    .B2(_05067_),
    .X(_04315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07708_ (.A1_N(_04957_),
    .A2_N(_05065_),
    .B1(\design_top.MEM[12][16] ),
    .B2(_05067_),
    .X(_04314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07709_ (.A(_04718_),
    .X(_05069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07710_ (.A(_04870_),
    .X(_05070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07711_ (.A(_05070_),
    .B(_05007_),
    .X(_05071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07712_ (.A(_05071_),
    .X(_05072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07713_ (.A(_05010_),
    .B_N(_05071_),
    .Y(_05073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07714_ (.A(_05073_),
    .X(_05074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07715_ (.A1_N(_05069_),
    .A2_N(_05072_),
    .B1(\design_top.MEM[12][31] ),
    .B2(_05074_),
    .X(_04313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07716_ (.A(_04889_),
    .X(_05075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07717_ (.A1_N(_05075_),
    .A2_N(_05072_),
    .B1(\design_top.MEM[12][30] ),
    .B2(_05074_),
    .X(_04312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07718_ (.A(_04891_),
    .X(_05076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07719_ (.A1_N(_05076_),
    .A2_N(_05072_),
    .B1(\design_top.MEM[12][29] ),
    .B2(_05074_),
    .X(_04311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07720_ (.A(_04893_),
    .X(_05077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07721_ (.A1_N(_05077_),
    .A2_N(_05072_),
    .B1(\design_top.MEM[12][28] ),
    .B2(_05074_),
    .X(_04310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07722_ (.A(_04895_),
    .X(_05078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07723_ (.A1_N(_05078_),
    .A2_N(_05072_),
    .B1(\design_top.MEM[12][27] ),
    .B2(_05074_),
    .X(_04309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07724_ (.A(_04897_),
    .X(_05079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07725_ (.A1_N(_05079_),
    .A2_N(_05071_),
    .B1(\design_top.MEM[12][26] ),
    .B2(_05073_),
    .X(_04308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07726_ (.A(_04899_),
    .X(_05080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07727_ (.A1_N(_05080_),
    .A2_N(_05071_),
    .B1(\design_top.MEM[12][25] ),
    .B2(_05073_),
    .X(_04307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07728_ (.A(_04901_),
    .X(_05081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07729_ (.A1_N(_05081_),
    .A2_N(_05071_),
    .B1(\design_top.MEM[12][24] ),
    .B2(_05073_),
    .X(_04306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07730_ (.A(_04903_),
    .X(_05082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07731_ (.A(_04873_),
    .B(_04905_),
    .X(_05083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07732_ (.A(_05006_),
    .B(_05083_),
    .X(_05084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07733_ (.A(_05084_),
    .X(_05085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _07734_ (.A(_04913_),
    .B(_04880_),
    .C(_04885_),
    .Y(_05086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07735_ (.A(_05086_),
    .B_N(_05084_),
    .Y(_05087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07736_ (.A(_05087_),
    .X(_05088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07737_ (.A1_N(_05082_),
    .A2_N(_05085_),
    .B1(\design_top.MEM[13][15] ),
    .B2(_05088_),
    .X(_04305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07738_ (.A(_04918_),
    .X(_05089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07739_ (.A1_N(_05089_),
    .A2_N(_05085_),
    .B1(\design_top.MEM[13][14] ),
    .B2(_05088_),
    .X(_04304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07740_ (.A(_04920_),
    .X(_05090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07741_ (.A1_N(_05090_),
    .A2_N(_05085_),
    .B1(\design_top.MEM[13][13] ),
    .B2(_05088_),
    .X(_04303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07742_ (.A(_04922_),
    .X(_05091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07743_ (.A1_N(_05091_),
    .A2_N(_05085_),
    .B1(\design_top.MEM[13][12] ),
    .B2(_05088_),
    .X(_04302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07744_ (.A(_04924_),
    .X(_05092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07745_ (.A1_N(_05092_),
    .A2_N(_05085_),
    .B1(\design_top.MEM[13][11] ),
    .B2(_05088_),
    .X(_04301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07746_ (.A(_04926_),
    .X(_05093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07747_ (.A1_N(_05093_),
    .A2_N(_05084_),
    .B1(\design_top.MEM[13][10] ),
    .B2(_05087_),
    .X(_04300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07748_ (.A(_04928_),
    .X(_05094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07749_ (.A1_N(_05094_),
    .A2_N(_05084_),
    .B1(\design_top.MEM[13][9] ),
    .B2(_05087_),
    .X(_04299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07750_ (.A(_04930_),
    .X(_05095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07751_ (.A1_N(_05095_),
    .A2_N(_05084_),
    .B1(\design_top.MEM[13][8] ),
    .B2(_05087_),
    .X(_04298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07752_ (.A(_04936_),
    .X(_05096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07753_ (.A(_05064_),
    .B(_05083_),
    .X(_05097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07754_ (.A(_05097_),
    .X(_05098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07755_ (.A(_05086_),
    .B_N(_05097_),
    .Y(_05099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07756_ (.A(_05099_),
    .X(_05100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07757_ (.A1_N(_05096_),
    .A2_N(_05098_),
    .B1(\design_top.MEM[13][23] ),
    .B2(_05100_),
    .X(_04297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07758_ (.A(_04944_),
    .X(_05101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07759_ (.A1_N(_05101_),
    .A2_N(_05098_),
    .B1(\design_top.MEM[13][22] ),
    .B2(_05100_),
    .X(_04296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07760_ (.A(_04946_),
    .X(_05102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07761_ (.A1_N(_05102_),
    .A2_N(_05098_),
    .B1(\design_top.MEM[13][21] ),
    .B2(_05100_),
    .X(_04295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07762_ (.A(_04948_),
    .X(_05103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07763_ (.A1_N(_05103_),
    .A2_N(_05098_),
    .B1(\design_top.MEM[13][20] ),
    .B2(_05100_),
    .X(_04294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07764_ (.A(_04950_),
    .X(_05104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07765_ (.A1_N(_05104_),
    .A2_N(_05098_),
    .B1(\design_top.MEM[13][19] ),
    .B2(_05100_),
    .X(_04293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07766_ (.A(_04952_),
    .X(_05105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07767_ (.A1_N(_05105_),
    .A2_N(_05097_),
    .B1(\design_top.MEM[13][18] ),
    .B2(_05099_),
    .X(_04292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07768_ (.A(_04954_),
    .X(_05106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07769_ (.A1_N(_05106_),
    .A2_N(_05097_),
    .B1(\design_top.MEM[13][17] ),
    .B2(_05099_),
    .X(_04291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07770_ (.A(_04956_),
    .X(_05107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07771_ (.A1_N(_05107_),
    .A2_N(_05097_),
    .B1(\design_top.MEM[13][16] ),
    .B2(_05099_),
    .X(_04290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07772_ (.A(_04905_),
    .B(_04990_),
    .X(_05108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07773_ (.A(_05006_),
    .B(_05108_),
    .X(_05109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07774_ (.A(_05109_),
    .X(_05110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _07775_ (.A(_04913_),
    .B(_04880_),
    .C(_04994_),
    .Y(_05111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07776_ (.A(_05111_),
    .B_N(_05109_),
    .Y(_05112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07777_ (.A(_05112_),
    .X(_05113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07778_ (.A1_N(_05082_),
    .A2_N(_05110_),
    .B1(\design_top.MEM[15][15] ),
    .B2(_05113_),
    .X(_04289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07779_ (.A1_N(_05089_),
    .A2_N(_05110_),
    .B1(\design_top.MEM[15][14] ),
    .B2(_05113_),
    .X(_04288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07780_ (.A1_N(_05090_),
    .A2_N(_05110_),
    .B1(\design_top.MEM[15][13] ),
    .B2(_05113_),
    .X(_04287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07781_ (.A1_N(_05091_),
    .A2_N(_05110_),
    .B1(\design_top.MEM[15][12] ),
    .B2(_05113_),
    .X(_04286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07782_ (.A1_N(_05092_),
    .A2_N(_05110_),
    .B1(\design_top.MEM[15][11] ),
    .B2(_05113_),
    .X(_04285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07783_ (.A1_N(_05093_),
    .A2_N(_05109_),
    .B1(\design_top.MEM[15][10] ),
    .B2(_05112_),
    .X(_04284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07784_ (.A1_N(_05094_),
    .A2_N(_05109_),
    .B1(\design_top.MEM[15][9] ),
    .B2(_05112_),
    .X(_04283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07785_ (.A1_N(_05095_),
    .A2_N(_05109_),
    .B1(\design_top.MEM[15][8] ),
    .B2(_05112_),
    .X(_04282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07786_ (.A(_05064_),
    .B(_05108_),
    .X(_05114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07787_ (.A(_05114_),
    .X(_05115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07788_ (.A(_05111_),
    .B_N(_05114_),
    .Y(_05116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07789_ (.A(_05116_),
    .X(_05117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07790_ (.A1_N(_05096_),
    .A2_N(_05115_),
    .B1(\design_top.MEM[15][23] ),
    .B2(_05117_),
    .X(_04281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07791_ (.A1_N(_05101_),
    .A2_N(_05115_),
    .B1(\design_top.MEM[15][22] ),
    .B2(_05117_),
    .X(_04280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07792_ (.A1_N(_05102_),
    .A2_N(_05115_),
    .B1(\design_top.MEM[15][21] ),
    .B2(_05117_),
    .X(_04279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07793_ (.A1_N(_05103_),
    .A2_N(_05115_),
    .B1(\design_top.MEM[15][20] ),
    .B2(_05117_),
    .X(_04278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07794_ (.A1_N(_05104_),
    .A2_N(_05115_),
    .B1(\design_top.MEM[15][19] ),
    .B2(_05117_),
    .X(_04277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07795_ (.A1_N(_05105_),
    .A2_N(_05114_),
    .B1(\design_top.MEM[15][18] ),
    .B2(_05116_),
    .X(_04276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07796_ (.A1_N(_05106_),
    .A2_N(_05114_),
    .B1(\design_top.MEM[15][17] ),
    .B2(_05116_),
    .X(_04275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07797_ (.A1_N(_05107_),
    .A2_N(_05114_),
    .B1(\design_top.MEM[15][16] ),
    .B2(_05116_),
    .X(_04274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07798_ (.A(_05070_),
    .B(_05108_),
    .X(_05118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07799_ (.A(_05118_),
    .X(_05119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07800_ (.A(_05111_),
    .B_N(_05118_),
    .Y(_05120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07801_ (.A(_05120_),
    .X(_05121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07802_ (.A1_N(_05069_),
    .A2_N(_05119_),
    .B1(\design_top.MEM[15][31] ),
    .B2(_05121_),
    .X(_04273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07803_ (.A1_N(_05075_),
    .A2_N(_05119_),
    .B1(\design_top.MEM[15][30] ),
    .B2(_05121_),
    .X(_04272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07804_ (.A1_N(_05076_),
    .A2_N(_05119_),
    .B1(\design_top.MEM[15][29] ),
    .B2(_05121_),
    .X(_04271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07805_ (.A1_N(_05077_),
    .A2_N(_05119_),
    .B1(\design_top.MEM[15][28] ),
    .B2(_05121_),
    .X(_04270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07806_ (.A1_N(_05078_),
    .A2_N(_05119_),
    .B1(\design_top.MEM[15][27] ),
    .B2(_05121_),
    .X(_04269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07807_ (.A1_N(_05079_),
    .A2_N(_05118_),
    .B1(\design_top.MEM[15][26] ),
    .B2(_05120_),
    .X(_04268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07808_ (.A1_N(_05080_),
    .A2_N(_05118_),
    .B1(\design_top.MEM[15][25] ),
    .B2(_05120_),
    .X(_04267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07809_ (.A1_N(_05081_),
    .A2_N(_05118_),
    .B1(\design_top.MEM[15][24] ),
    .B2(_05120_),
    .X(_04266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07810_ (.A(_04873_),
    .B(_04959_),
    .X(_05122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07811_ (.A(_05064_),
    .B(_05122_),
    .X(_05123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07812_ (.A(_05123_),
    .X(_05124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _07813_ (.A(_04879_),
    .B(_04963_),
    .C(_04885_),
    .Y(_05125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07814_ (.A(_05125_),
    .B_N(_05123_),
    .Y(_05126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07815_ (.A(_05126_),
    .X(_05127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07816_ (.A1_N(_05096_),
    .A2_N(_05124_),
    .B1(\design_top.MEM[1][23] ),
    .B2(_05127_),
    .X(_04265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07817_ (.A1_N(_05101_),
    .A2_N(_05124_),
    .B1(\design_top.MEM[1][22] ),
    .B2(_05127_),
    .X(_04264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07818_ (.A1_N(_05102_),
    .A2_N(_05124_),
    .B1(\design_top.MEM[1][21] ),
    .B2(_05127_),
    .X(_04263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07819_ (.A1_N(_05103_),
    .A2_N(_05124_),
    .B1(\design_top.MEM[1][20] ),
    .B2(_05127_),
    .X(_04262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07820_ (.A1_N(_05104_),
    .A2_N(_05124_),
    .B1(\design_top.MEM[1][19] ),
    .B2(_05127_),
    .X(_04261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07821_ (.A1_N(_05105_),
    .A2_N(_05123_),
    .B1(\design_top.MEM[1][18] ),
    .B2(_05126_),
    .X(_04260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07822_ (.A1_N(_05106_),
    .A2_N(_05123_),
    .B1(\design_top.MEM[1][17] ),
    .B2(_05126_),
    .X(_04259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07823_ (.A1_N(_05107_),
    .A2_N(_05123_),
    .B1(\design_top.MEM[1][16] ),
    .B2(_05126_),
    .X(_04258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07824_ (.A(_05070_),
    .B(_05122_),
    .X(_05128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07825_ (.A(_05128_),
    .X(_05129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07826_ (.A(_05125_),
    .B_N(_05128_),
    .Y(_05130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07827_ (.A(_05130_),
    .X(_05131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07828_ (.A1_N(_05069_),
    .A2_N(_05129_),
    .B1(\design_top.MEM[1][31] ),
    .B2(_05131_),
    .X(_04257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07829_ (.A1_N(_05075_),
    .A2_N(_05129_),
    .B1(\design_top.MEM[1][30] ),
    .B2(_05131_),
    .X(_04256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07830_ (.A1_N(_05076_),
    .A2_N(_05129_),
    .B1(\design_top.MEM[1][29] ),
    .B2(_05131_),
    .X(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07831_ (.A1_N(_05077_),
    .A2_N(_05129_),
    .B1(\design_top.MEM[1][28] ),
    .B2(_05131_),
    .X(_04254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07832_ (.A1_N(_05078_),
    .A2_N(_05129_),
    .B1(\design_top.MEM[1][27] ),
    .B2(_05131_),
    .X(_04253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07833_ (.A1_N(_05079_),
    .A2_N(_05128_),
    .B1(\design_top.MEM[1][26] ),
    .B2(_05130_),
    .X(_04252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07834_ (.A1_N(_05080_),
    .A2_N(_05128_),
    .B1(\design_top.MEM[1][25] ),
    .B2(_05130_),
    .X(_04251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07835_ (.A1_N(_05081_),
    .A2_N(_05128_),
    .B1(\design_top.MEM[1][24] ),
    .B2(_05130_),
    .X(_04250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07836_ (.A(_05006_),
    .B(_05122_),
    .X(_05132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07837_ (.A(_05132_),
    .X(_05133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07838_ (.A(_05125_),
    .B_N(_05132_),
    .Y(_05134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07839_ (.A(_05134_),
    .X(_05135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07840_ (.A1_N(_05082_),
    .A2_N(_05133_),
    .B1(\design_top.MEM[1][15] ),
    .B2(_05135_),
    .X(_04249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07841_ (.A1_N(_05089_),
    .A2_N(_05133_),
    .B1(\design_top.MEM[1][14] ),
    .B2(_05135_),
    .X(_04248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07842_ (.A1_N(_05090_),
    .A2_N(_05133_),
    .B1(\design_top.MEM[1][13] ),
    .B2(_05135_),
    .X(_04247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07843_ (.A1_N(_05091_),
    .A2_N(_05133_),
    .B1(\design_top.MEM[1][12] ),
    .B2(_05135_),
    .X(_04246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07844_ (.A1_N(_05092_),
    .A2_N(_05133_),
    .B1(\design_top.MEM[1][11] ),
    .B2(_05135_),
    .X(_04245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07845_ (.A1_N(_05093_),
    .A2_N(_05132_),
    .B1(\design_top.MEM[1][10] ),
    .B2(_05134_),
    .X(_04244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07846_ (.A1_N(_05094_),
    .A2_N(_05132_),
    .B1(\design_top.MEM[1][9] ),
    .B2(_05134_),
    .X(_04243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07847_ (.A1_N(_05095_),
    .A2_N(_05132_),
    .B1(\design_top.MEM[1][8] ),
    .B2(_05134_),
    .X(_04242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07848_ (.A(_04906_),
    .B(_04959_),
    .X(_05136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07849_ (.A(_05006_),
    .B(_05136_),
    .X(_05137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07850_ (.A(_05137_),
    .X(_05138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _07851_ (.A(wbs_adr_i[0]),
    .B(_04963_),
    .C(_04914_),
    .Y(_05139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07852_ (.A(_05139_),
    .B_N(_05137_),
    .Y(_05140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07853_ (.A(_05140_),
    .X(_05141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07854_ (.A1_N(_05082_),
    .A2_N(_05138_),
    .B1(\design_top.MEM[2][15] ),
    .B2(_05141_),
    .X(_04241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07855_ (.A1_N(_05089_),
    .A2_N(_05138_),
    .B1(\design_top.MEM[2][14] ),
    .B2(_05141_),
    .X(_04240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07856_ (.A1_N(_05090_),
    .A2_N(_05138_),
    .B1(\design_top.MEM[2][13] ),
    .B2(_05141_),
    .X(_04239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07857_ (.A1_N(_05091_),
    .A2_N(_05138_),
    .B1(\design_top.MEM[2][12] ),
    .B2(_05141_),
    .X(_04238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07858_ (.A1_N(_05092_),
    .A2_N(_05138_),
    .B1(\design_top.MEM[2][11] ),
    .B2(_05141_),
    .X(_04237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07859_ (.A1_N(_05093_),
    .A2_N(_05137_),
    .B1(\design_top.MEM[2][10] ),
    .B2(_05140_),
    .X(_04236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07860_ (.A1_N(_05094_),
    .A2_N(_05137_),
    .B1(\design_top.MEM[2][9] ),
    .B2(_05140_),
    .X(_04235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07861_ (.A1_N(_05095_),
    .A2_N(_05137_),
    .B1(\design_top.MEM[2][8] ),
    .B2(_05140_),
    .X(_04234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07862_ (.A(_05064_),
    .B(_05136_),
    .X(_05142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07863_ (.A(_05142_),
    .X(_05143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07864_ (.A(_05139_),
    .B_N(_05142_),
    .Y(_05144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07865_ (.A(_05144_),
    .X(_05145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07866_ (.A1_N(_05096_),
    .A2_N(_05143_),
    .B1(\design_top.MEM[2][23] ),
    .B2(_05145_),
    .X(_04233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07867_ (.A1_N(_05101_),
    .A2_N(_05143_),
    .B1(\design_top.MEM[2][22] ),
    .B2(_05145_),
    .X(_04232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07868_ (.A1_N(_05102_),
    .A2_N(_05143_),
    .B1(\design_top.MEM[2][21] ),
    .B2(_05145_),
    .X(_04231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07869_ (.A1_N(_05103_),
    .A2_N(_05143_),
    .B1(\design_top.MEM[2][20] ),
    .B2(_05145_),
    .X(_04230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07870_ (.A1_N(_05104_),
    .A2_N(_05143_),
    .B1(\design_top.MEM[2][19] ),
    .B2(_05145_),
    .X(_04229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07871_ (.A1_N(_05105_),
    .A2_N(_05142_),
    .B1(\design_top.MEM[2][18] ),
    .B2(_05144_),
    .X(_04228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07872_ (.A1_N(_05106_),
    .A2_N(_05142_),
    .B1(\design_top.MEM[2][17] ),
    .B2(_05144_),
    .X(_04227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07873_ (.A1_N(_05107_),
    .A2_N(_05142_),
    .B1(\design_top.MEM[2][16] ),
    .B2(_05144_),
    .X(_04226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07874_ (.A(_05070_),
    .B(_05136_),
    .X(_05146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07875_ (.A(_05146_),
    .X(_05147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07876_ (.A(_05139_),
    .B_N(_05146_),
    .Y(_05148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07877_ (.A(_05148_),
    .X(_05149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07878_ (.A1_N(_05069_),
    .A2_N(_05147_),
    .B1(\design_top.MEM[2][31] ),
    .B2(_05149_),
    .X(_04225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07879_ (.A1_N(_05075_),
    .A2_N(_05147_),
    .B1(\design_top.MEM[2][30] ),
    .B2(_05149_),
    .X(_04224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07880_ (.A1_N(_05076_),
    .A2_N(_05147_),
    .B1(\design_top.MEM[2][29] ),
    .B2(_05149_),
    .X(_04223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07881_ (.A1_N(_05077_),
    .A2_N(_05147_),
    .B1(\design_top.MEM[2][28] ),
    .B2(_05149_),
    .X(_04222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07882_ (.A1_N(_05078_),
    .A2_N(_05147_),
    .B1(\design_top.MEM[2][27] ),
    .B2(_05149_),
    .X(_04221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07883_ (.A1_N(_05079_),
    .A2_N(_05146_),
    .B1(\design_top.MEM[2][26] ),
    .B2(_05148_),
    .X(_04220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07884_ (.A1_N(_05080_),
    .A2_N(_05146_),
    .B1(\design_top.MEM[2][25] ),
    .B2(_05148_),
    .X(_04219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07885_ (.A1_N(_05081_),
    .A2_N(_05146_),
    .B1(\design_top.MEM[2][24] ),
    .B2(_05148_),
    .X(_04218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07886_ (.A(_04908_),
    .X(_05150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07887_ (.A(_04959_),
    .B(_04990_),
    .X(_05151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07888_ (.A(_05150_),
    .B(_05151_),
    .X(_05152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07889_ (.A(_05152_),
    .X(_05153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _07890_ (.A(wbs_adr_i[0]),
    .B(_04963_),
    .C(_04994_),
    .Y(_05154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07891_ (.A(_05154_),
    .B_N(_05152_),
    .Y(_05155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07892_ (.A(_05155_),
    .X(_05156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07893_ (.A1_N(_05082_),
    .A2_N(_05153_),
    .B1(\design_top.MEM[3][15] ),
    .B2(_05156_),
    .X(_04217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07894_ (.A1_N(_05089_),
    .A2_N(_05153_),
    .B1(\design_top.MEM[3][14] ),
    .B2(_05156_),
    .X(_04216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07895_ (.A1_N(_05090_),
    .A2_N(_05153_),
    .B1(\design_top.MEM[3][13] ),
    .B2(_05156_),
    .X(_04215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07896_ (.A1_N(_05091_),
    .A2_N(_05153_),
    .B1(\design_top.MEM[3][12] ),
    .B2(_05156_),
    .X(_04214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07897_ (.A1_N(_05092_),
    .A2_N(_05153_),
    .B1(\design_top.MEM[3][11] ),
    .B2(_05156_),
    .X(_04213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07898_ (.A1_N(_05093_),
    .A2_N(_05152_),
    .B1(\design_top.MEM[3][10] ),
    .B2(_05155_),
    .X(_04212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07899_ (.A1_N(_05094_),
    .A2_N(_05152_),
    .B1(\design_top.MEM[3][9] ),
    .B2(_05155_),
    .X(_04211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07900_ (.A1_N(_05095_),
    .A2_N(_05152_),
    .B1(\design_top.MEM[3][8] ),
    .B2(_05155_),
    .X(_04210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07901_ (.A(_04938_),
    .X(_05157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07902_ (.A(_05157_),
    .B(_05151_),
    .X(_05158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07903_ (.A(_05158_),
    .X(_05159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07904_ (.A(_05154_),
    .B_N(_05158_),
    .Y(_05160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07905_ (.A(_05160_),
    .X(_05161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07906_ (.A1_N(_05096_),
    .A2_N(_05159_),
    .B1(\design_top.MEM[3][23] ),
    .B2(_05161_),
    .X(_04209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07907_ (.A1_N(_05101_),
    .A2_N(_05159_),
    .B1(\design_top.MEM[3][22] ),
    .B2(_05161_),
    .X(_04208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07908_ (.A1_N(_05102_),
    .A2_N(_05159_),
    .B1(\design_top.MEM[3][21] ),
    .B2(_05161_),
    .X(_04207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07909_ (.A1_N(_05103_),
    .A2_N(_05159_),
    .B1(\design_top.MEM[3][20] ),
    .B2(_05161_),
    .X(_04206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07910_ (.A1_N(_05104_),
    .A2_N(_05159_),
    .B1(\design_top.MEM[3][19] ),
    .B2(_05161_),
    .X(_04205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07911_ (.A1_N(_05105_),
    .A2_N(_05158_),
    .B1(\design_top.MEM[3][18] ),
    .B2(_05160_),
    .X(_04204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07912_ (.A1_N(_05106_),
    .A2_N(_05158_),
    .B1(\design_top.MEM[3][17] ),
    .B2(_05160_),
    .X(_04203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07913_ (.A1_N(_05107_),
    .A2_N(_05158_),
    .B1(\design_top.MEM[3][16] ),
    .B2(_05160_),
    .X(_04202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07914_ (.A(_05070_),
    .B(_05151_),
    .X(_05162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07915_ (.A(_05162_),
    .X(_05163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07916_ (.A(_05154_),
    .B_N(_05162_),
    .Y(_05164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07917_ (.A(_05164_),
    .X(_05165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07918_ (.A1_N(_05069_),
    .A2_N(_05163_),
    .B1(\design_top.MEM[3][31] ),
    .B2(_05165_),
    .X(_04201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07919_ (.A1_N(_05075_),
    .A2_N(_05163_),
    .B1(\design_top.MEM[3][30] ),
    .B2(_05165_),
    .X(_04200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07920_ (.A1_N(_05076_),
    .A2_N(_05163_),
    .B1(\design_top.MEM[3][29] ),
    .B2(_05165_),
    .X(_04199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07921_ (.A1_N(_05077_),
    .A2_N(_05163_),
    .B1(\design_top.MEM[3][28] ),
    .B2(_05165_),
    .X(_04198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07922_ (.A1_N(_05078_),
    .A2_N(_05163_),
    .B1(\design_top.MEM[3][27] ),
    .B2(_05165_),
    .X(_04197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07923_ (.A1_N(_05079_),
    .A2_N(_05162_),
    .B1(\design_top.MEM[3][26] ),
    .B2(_05164_),
    .X(_04196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07924_ (.A1_N(_05080_),
    .A2_N(_05162_),
    .B1(\design_top.MEM[3][25] ),
    .B2(_05164_),
    .X(_04195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07925_ (.A1_N(_05081_),
    .A2_N(_05162_),
    .B1(\design_top.MEM[3][24] ),
    .B2(_05164_),
    .X(_04194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07926_ (.A(_04903_),
    .X(_05166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07927_ (.A(_00353_),
    .B(_02415_),
    .X(_05167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07928_ (.A(_04958_),
    .B(_05167_),
    .X(_05168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07929_ (.A(_05150_),
    .B(_05168_),
    .X(_05169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07930_ (.A(_05169_),
    .X(_05170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _07931_ (.A(_04913_),
    .B(_04963_),
    .C(_04964_),
    .Y(_05171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07932_ (.A(_05171_),
    .B_N(_05169_),
    .Y(_05172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07933_ (.A(_05172_),
    .X(_05173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07934_ (.A1_N(_05166_),
    .A2_N(_05170_),
    .B1(\design_top.MEM[4][15] ),
    .B2(_05173_),
    .X(_04193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07935_ (.A(_04918_),
    .X(_05174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07936_ (.A1_N(_05174_),
    .A2_N(_05170_),
    .B1(\design_top.MEM[4][14] ),
    .B2(_05173_),
    .X(_04192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07937_ (.A(_04920_),
    .X(_05175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07938_ (.A1_N(_05175_),
    .A2_N(_05170_),
    .B1(\design_top.MEM[4][13] ),
    .B2(_05173_),
    .X(_04191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07939_ (.A(_04922_),
    .X(_05176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07940_ (.A1_N(_05176_),
    .A2_N(_05170_),
    .B1(\design_top.MEM[4][12] ),
    .B2(_05173_),
    .X(_04190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07941_ (.A(_04924_),
    .X(_05177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07942_ (.A1_N(_05177_),
    .A2_N(_05170_),
    .B1(\design_top.MEM[4][11] ),
    .B2(_05173_),
    .X(_04189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07943_ (.A(_04926_),
    .X(_05178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07944_ (.A1_N(_05178_),
    .A2_N(_05169_),
    .B1(\design_top.MEM[4][10] ),
    .B2(_05172_),
    .X(_04188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07945_ (.A(_04928_),
    .X(_05179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07946_ (.A1_N(_05179_),
    .A2_N(_05169_),
    .B1(\design_top.MEM[4][9] ),
    .B2(_05172_),
    .X(_04187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07947_ (.A(_04930_),
    .X(_05180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07948_ (.A1_N(_05180_),
    .A2_N(_05169_),
    .B1(\design_top.MEM[4][8] ),
    .B2(_05172_),
    .X(_04186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07949_ (.A(_04936_),
    .X(_05181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07950_ (.A(_05157_),
    .B(_05168_),
    .X(_05182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07951_ (.A(_05182_),
    .X(_05183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07952_ (.A(_05171_),
    .B_N(_05182_),
    .Y(_05184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07953_ (.A(_05184_),
    .X(_05185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07954_ (.A1_N(_05181_),
    .A2_N(_05183_),
    .B1(\design_top.MEM[4][23] ),
    .B2(_05185_),
    .X(_04185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07955_ (.A(_04944_),
    .X(_05186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07956_ (.A1_N(_05186_),
    .A2_N(_05183_),
    .B1(\design_top.MEM[4][22] ),
    .B2(_05185_),
    .X(_04184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07957_ (.A(_04946_),
    .X(_05187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07958_ (.A1_N(_05187_),
    .A2_N(_05183_),
    .B1(\design_top.MEM[4][21] ),
    .B2(_05185_),
    .X(_04183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07959_ (.A(_04948_),
    .X(_05188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07960_ (.A1_N(_05188_),
    .A2_N(_05183_),
    .B1(\design_top.MEM[4][20] ),
    .B2(_05185_),
    .X(_04182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07961_ (.A(_04950_),
    .X(_05189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07962_ (.A1_N(_05189_),
    .A2_N(_05183_),
    .B1(\design_top.MEM[4][19] ),
    .B2(_05185_),
    .X(_04181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07963_ (.A(_04952_),
    .X(_05190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07964_ (.A1_N(_05190_),
    .A2_N(_05182_),
    .B1(\design_top.MEM[4][18] ),
    .B2(_05184_),
    .X(_04180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07965_ (.A(_04954_),
    .X(_05191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07966_ (.A1_N(_05191_),
    .A2_N(_05182_),
    .B1(\design_top.MEM[4][17] ),
    .B2(_05184_),
    .X(_04179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07967_ (.A(_04956_),
    .X(_05192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07968_ (.A1_N(_05192_),
    .A2_N(_05182_),
    .B1(\design_top.MEM[4][16] ),
    .B2(_05184_),
    .X(_04178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07969_ (.A(_04718_),
    .X(_05193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07970_ (.A(_04870_),
    .X(_05194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07971_ (.A(_05194_),
    .B(_05168_),
    .X(_05195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07972_ (.A(_05195_),
    .X(_05196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07973_ (.A(_05171_),
    .B_N(_05195_),
    .Y(_05197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07974_ (.A(_05197_),
    .X(_05198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07975_ (.A1_N(_05193_),
    .A2_N(_05196_),
    .B1(\design_top.MEM[4][31] ),
    .B2(_05198_),
    .X(_04177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07976_ (.A(_04889_),
    .X(_05199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07977_ (.A1_N(_05199_),
    .A2_N(_05196_),
    .B1(\design_top.MEM[4][30] ),
    .B2(_05198_),
    .X(_04176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07978_ (.A(_04891_),
    .X(_05200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07979_ (.A1_N(_05200_),
    .A2_N(_05196_),
    .B1(\design_top.MEM[4][29] ),
    .B2(_05198_),
    .X(_04175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07980_ (.A(_04893_),
    .X(_05201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07981_ (.A1_N(_05201_),
    .A2_N(_05196_),
    .B1(\design_top.MEM[4][28] ),
    .B2(_05198_),
    .X(_04174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07982_ (.A(_04895_),
    .X(_05202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07983_ (.A1_N(_05202_),
    .A2_N(_05196_),
    .B1(\design_top.MEM[4][27] ),
    .B2(_05198_),
    .X(_04173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07984_ (.A(_04897_),
    .X(_05203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07985_ (.A1_N(_05203_),
    .A2_N(_05195_),
    .B1(\design_top.MEM[4][26] ),
    .B2(_05197_),
    .X(_04172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07986_ (.A(_04899_),
    .X(_05204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07987_ (.A1_N(_05204_),
    .A2_N(_05195_),
    .B1(\design_top.MEM[4][25] ),
    .B2(_05197_),
    .X(_04171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07988_ (.A(_04901_),
    .X(_05205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07989_ (.A1_N(_05205_),
    .A2_N(_05195_),
    .B1(\design_top.MEM[4][24] ),
    .B2(_05197_),
    .X(_04170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07990_ (.A(_04873_),
    .B(_05167_),
    .X(_05206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _07991_ (.A(_05150_),
    .B(_05206_),
    .X(_05207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07992_ (.A(_05207_),
    .X(_05208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _07993_ (.A(_04912_),
    .B(wbs_adr_i[1]),
    .C(_04885_),
    .Y(_05209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _07994_ (.A(_05209_),
    .B_N(_05207_),
    .Y(_05210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _07995_ (.A(_05210_),
    .X(_05211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07996_ (.A1_N(_05166_),
    .A2_N(_05208_),
    .B1(\design_top.MEM[5][15] ),
    .B2(_05211_),
    .X(_04169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07997_ (.A1_N(_05174_),
    .A2_N(_05208_),
    .B1(\design_top.MEM[5][14] ),
    .B2(_05211_),
    .X(_04168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07998_ (.A1_N(_05175_),
    .A2_N(_05208_),
    .B1(\design_top.MEM[5][13] ),
    .B2(_05211_),
    .X(_04167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _07999_ (.A1_N(_05176_),
    .A2_N(_05208_),
    .B1(\design_top.MEM[5][12] ),
    .B2(_05211_),
    .X(_04166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08000_ (.A1_N(_05177_),
    .A2_N(_05208_),
    .B1(\design_top.MEM[5][11] ),
    .B2(_05211_),
    .X(_04165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08001_ (.A1_N(_05178_),
    .A2_N(_05207_),
    .B1(\design_top.MEM[5][10] ),
    .B2(_05210_),
    .X(_04164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08002_ (.A1_N(_05179_),
    .A2_N(_05207_),
    .B1(\design_top.MEM[5][9] ),
    .B2(_05210_),
    .X(_04163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08003_ (.A1_N(_05180_),
    .A2_N(_05207_),
    .B1(\design_top.MEM[5][8] ),
    .B2(_05210_),
    .X(_04162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08004_ (.A(_05157_),
    .B(_05206_),
    .X(_05212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08005_ (.A(_05212_),
    .X(_05213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _08006_ (.A(_05209_),
    .B_N(_05212_),
    .Y(_05214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08007_ (.A(_05214_),
    .X(_05215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08008_ (.A1_N(_05181_),
    .A2_N(_05213_),
    .B1(\design_top.MEM[5][23] ),
    .B2(_05215_),
    .X(_04161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08009_ (.A1_N(_05186_),
    .A2_N(_05213_),
    .B1(\design_top.MEM[5][22] ),
    .B2(_05215_),
    .X(_04160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08010_ (.A1_N(_05187_),
    .A2_N(_05213_),
    .B1(\design_top.MEM[5][21] ),
    .B2(_05215_),
    .X(_04159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08011_ (.A1_N(_05188_),
    .A2_N(_05213_),
    .B1(\design_top.MEM[5][20] ),
    .B2(_05215_),
    .X(_04158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08012_ (.A1_N(_05189_),
    .A2_N(_05213_),
    .B1(\design_top.MEM[5][19] ),
    .B2(_05215_),
    .X(_04157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08013_ (.A1_N(_05190_),
    .A2_N(_05212_),
    .B1(\design_top.MEM[5][18] ),
    .B2(_05214_),
    .X(_04156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08014_ (.A1_N(_05191_),
    .A2_N(_05212_),
    .B1(\design_top.MEM[5][17] ),
    .B2(_05214_),
    .X(_04155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08015_ (.A1_N(_05192_),
    .A2_N(_05212_),
    .B1(\design_top.MEM[5][16] ),
    .B2(_05214_),
    .X(_04154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08016_ (.A(_05194_),
    .B(_05206_),
    .X(_05216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08017_ (.A(_05216_),
    .X(_05217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _08018_ (.A(_05209_),
    .B_N(_05216_),
    .Y(_05218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08019_ (.A(_05218_),
    .X(_05219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08020_ (.A1_N(_05193_),
    .A2_N(_05217_),
    .B1(\design_top.MEM[5][31] ),
    .B2(_05219_),
    .X(_04153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08021_ (.A1_N(_05199_),
    .A2_N(_05217_),
    .B1(\design_top.MEM[5][30] ),
    .B2(_05219_),
    .X(_04152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08022_ (.A1_N(_05200_),
    .A2_N(_05217_),
    .B1(\design_top.MEM[5][29] ),
    .B2(_05219_),
    .X(_04151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08023_ (.A1_N(_05201_),
    .A2_N(_05217_),
    .B1(\design_top.MEM[5][28] ),
    .B2(_05219_),
    .X(_04150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08024_ (.A1_N(_05202_),
    .A2_N(_05217_),
    .B1(\design_top.MEM[5][27] ),
    .B2(_05219_),
    .X(_04149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08025_ (.A1_N(_05203_),
    .A2_N(_05216_),
    .B1(\design_top.MEM[5][26] ),
    .B2(_05218_),
    .X(_04148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08026_ (.A1_N(_05204_),
    .A2_N(_05216_),
    .B1(\design_top.MEM[5][25] ),
    .B2(_05218_),
    .X(_04147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08027_ (.A1_N(_05205_),
    .A2_N(_05216_),
    .B1(\design_top.MEM[5][24] ),
    .B2(_05218_),
    .X(_04146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08028_ (.A(_04906_),
    .B(_05167_),
    .X(_05220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08029_ (.A(_05150_),
    .B(_05220_),
    .X(_05221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08030_ (.A(_05221_),
    .X(_05222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _08031_ (.A(_04912_),
    .B(wbs_adr_i[1]),
    .C(_04914_),
    .Y(_05223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _08032_ (.A(_05223_),
    .B_N(_05221_),
    .Y(_05224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08033_ (.A(_05224_),
    .X(_05225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08034_ (.A1_N(_05166_),
    .A2_N(_05222_),
    .B1(\design_top.MEM[6][15] ),
    .B2(_05225_),
    .X(_04145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08035_ (.A1_N(_05174_),
    .A2_N(_05222_),
    .B1(\design_top.MEM[6][14] ),
    .B2(_05225_),
    .X(_04144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08036_ (.A1_N(_05175_),
    .A2_N(_05222_),
    .B1(\design_top.MEM[6][13] ),
    .B2(_05225_),
    .X(_04143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08037_ (.A1_N(_05176_),
    .A2_N(_05222_),
    .B1(\design_top.MEM[6][12] ),
    .B2(_05225_),
    .X(_04142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08038_ (.A1_N(_05177_),
    .A2_N(_05222_),
    .B1(\design_top.MEM[6][11] ),
    .B2(_05225_),
    .X(_04141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08039_ (.A1_N(_05178_),
    .A2_N(_05221_),
    .B1(\design_top.MEM[6][10] ),
    .B2(_05224_),
    .X(_04140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08040_ (.A1_N(_05179_),
    .A2_N(_05221_),
    .B1(\design_top.MEM[6][9] ),
    .B2(_05224_),
    .X(_04139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08041_ (.A1_N(_05180_),
    .A2_N(_05221_),
    .B1(\design_top.MEM[6][8] ),
    .B2(_05224_),
    .X(_04138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08042_ (.A(_05157_),
    .B(_05220_),
    .X(_05226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08043_ (.A(_05226_),
    .X(_05227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _08044_ (.A(_05223_),
    .B_N(_05226_),
    .Y(_05228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08045_ (.A(_05228_),
    .X(_05229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08046_ (.A1_N(_05181_),
    .A2_N(_05227_),
    .B1(\design_top.MEM[6][23] ),
    .B2(_05229_),
    .X(_04137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08047_ (.A1_N(_05186_),
    .A2_N(_05227_),
    .B1(\design_top.MEM[6][22] ),
    .B2(_05229_),
    .X(_04136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08048_ (.A1_N(_05187_),
    .A2_N(_05227_),
    .B1(\design_top.MEM[6][21] ),
    .B2(_05229_),
    .X(_04135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08049_ (.A1_N(_05188_),
    .A2_N(_05227_),
    .B1(\design_top.MEM[6][20] ),
    .B2(_05229_),
    .X(_04134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08050_ (.A1_N(_05189_),
    .A2_N(_05227_),
    .B1(\design_top.MEM[6][19] ),
    .B2(_05229_),
    .X(_04133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08051_ (.A1_N(_05190_),
    .A2_N(_05226_),
    .B1(\design_top.MEM[6][18] ),
    .B2(_05228_),
    .X(_04132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08052_ (.A1_N(_05191_),
    .A2_N(_05226_),
    .B1(\design_top.MEM[6][17] ),
    .B2(_05228_),
    .X(_04131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08053_ (.A1_N(_05192_),
    .A2_N(_05226_),
    .B1(\design_top.MEM[6][16] ),
    .B2(_05228_),
    .X(_04130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08054_ (.A(_05194_),
    .B(_05220_),
    .X(_05230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08055_ (.A(_05230_),
    .X(_05231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _08056_ (.A(_05223_),
    .B_N(_05230_),
    .Y(_05232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08057_ (.A(_05232_),
    .X(_05233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08058_ (.A1_N(_05193_),
    .A2_N(_05231_),
    .B1(\design_top.MEM[6][31] ),
    .B2(_05233_),
    .X(_04129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08059_ (.A1_N(_05199_),
    .A2_N(_05231_),
    .B1(\design_top.MEM[6][30] ),
    .B2(_05233_),
    .X(_04128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08060_ (.A1_N(_05200_),
    .A2_N(_05231_),
    .B1(\design_top.MEM[6][29] ),
    .B2(_05233_),
    .X(_04127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08061_ (.A1_N(_05201_),
    .A2_N(_05231_),
    .B1(\design_top.MEM[6][28] ),
    .B2(_05233_),
    .X(_04126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08062_ (.A1_N(_05202_),
    .A2_N(_05231_),
    .B1(\design_top.MEM[6][27] ),
    .B2(_05233_),
    .X(_04125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08063_ (.A1_N(_05203_),
    .A2_N(_05230_),
    .B1(\design_top.MEM[6][26] ),
    .B2(_05232_),
    .X(_04124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08064_ (.A1_N(_05204_),
    .A2_N(_05230_),
    .B1(\design_top.MEM[6][25] ),
    .B2(_05232_),
    .X(_04123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08065_ (.A1_N(_05205_),
    .A2_N(_05230_),
    .B1(\design_top.MEM[6][24] ),
    .B2(_05232_),
    .X(_04122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08066_ (.A(_04990_),
    .B(_05167_),
    .X(_05234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08067_ (.A(_05150_),
    .B(_05234_),
    .X(_05235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08068_ (.A(_05235_),
    .X(_05236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _08069_ (.A(_04912_),
    .B(wbs_adr_i[1]),
    .C(_04994_),
    .Y(_05237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _08070_ (.A(_05237_),
    .B_N(_05235_),
    .Y(_05238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08071_ (.A(_05238_),
    .X(_05239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08072_ (.A1_N(_05166_),
    .A2_N(_05236_),
    .B1(\design_top.MEM[7][15] ),
    .B2(_05239_),
    .X(_04121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08073_ (.A1_N(_05174_),
    .A2_N(_05236_),
    .B1(\design_top.MEM[7][14] ),
    .B2(_05239_),
    .X(_04120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08074_ (.A1_N(_05175_),
    .A2_N(_05236_),
    .B1(\design_top.MEM[7][13] ),
    .B2(_05239_),
    .X(_04119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08075_ (.A1_N(_05176_),
    .A2_N(_05236_),
    .B1(\design_top.MEM[7][12] ),
    .B2(_05239_),
    .X(_04118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08076_ (.A1_N(_05177_),
    .A2_N(_05236_),
    .B1(\design_top.MEM[7][11] ),
    .B2(_05239_),
    .X(_04117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08077_ (.A1_N(_05178_),
    .A2_N(_05235_),
    .B1(\design_top.MEM[7][10] ),
    .B2(_05238_),
    .X(_04116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08078_ (.A1_N(_05179_),
    .A2_N(_05235_),
    .B1(\design_top.MEM[7][9] ),
    .B2(_05238_),
    .X(_04115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08079_ (.A1_N(_05180_),
    .A2_N(_05235_),
    .B1(\design_top.MEM[7][8] ),
    .B2(_05238_),
    .X(_04114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08080_ (.A(_05157_),
    .B(_05234_),
    .X(_05240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08081_ (.A(_05240_),
    .X(_05241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _08082_ (.A(_05237_),
    .B_N(_05240_),
    .Y(_05242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08083_ (.A(_05242_),
    .X(_05243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08084_ (.A1_N(_05181_),
    .A2_N(_05241_),
    .B1(\design_top.MEM[7][23] ),
    .B2(_05243_),
    .X(_04113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08085_ (.A1_N(_05186_),
    .A2_N(_05241_),
    .B1(\design_top.MEM[7][22] ),
    .B2(_05243_),
    .X(_04112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08086_ (.A1_N(_05187_),
    .A2_N(_05241_),
    .B1(\design_top.MEM[7][21] ),
    .B2(_05243_),
    .X(_04111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08087_ (.A1_N(_05188_),
    .A2_N(_05241_),
    .B1(\design_top.MEM[7][20] ),
    .B2(_05243_),
    .X(_04110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08088_ (.A1_N(_05189_),
    .A2_N(_05241_),
    .B1(\design_top.MEM[7][19] ),
    .B2(_05243_),
    .X(_04109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08089_ (.A1_N(_05190_),
    .A2_N(_05240_),
    .B1(\design_top.MEM[7][18] ),
    .B2(_05242_),
    .X(_04108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08090_ (.A1_N(_05191_),
    .A2_N(_05240_),
    .B1(\design_top.MEM[7][17] ),
    .B2(_05242_),
    .X(_04107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08091_ (.A1_N(_05192_),
    .A2_N(_05240_),
    .B1(\design_top.MEM[7][16] ),
    .B2(_05242_),
    .X(_04106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08092_ (.A(_05194_),
    .B(_05234_),
    .X(_05244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08093_ (.A(_05244_),
    .X(_05245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _08094_ (.A(_05237_),
    .B_N(_05244_),
    .Y(_05246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08095_ (.A(_05246_),
    .X(_05247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08096_ (.A1_N(_05193_),
    .A2_N(_05245_),
    .B1(\design_top.MEM[7][31] ),
    .B2(_05247_),
    .X(_04105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08097_ (.A1_N(_05199_),
    .A2_N(_05245_),
    .B1(\design_top.MEM[7][30] ),
    .B2(_05247_),
    .X(_04104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08098_ (.A1_N(_05200_),
    .A2_N(_05245_),
    .B1(\design_top.MEM[7][29] ),
    .B2(_05247_),
    .X(_04103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08099_ (.A1_N(_05201_),
    .A2_N(_05245_),
    .B1(\design_top.MEM[7][28] ),
    .B2(_05247_),
    .X(_04102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08100_ (.A1_N(_05202_),
    .A2_N(_05245_),
    .B1(\design_top.MEM[7][27] ),
    .B2(_05247_),
    .X(_04101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08101_ (.A1_N(_05203_),
    .A2_N(_05244_),
    .B1(\design_top.MEM[7][26] ),
    .B2(_05246_),
    .X(_04100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08102_ (.A1_N(_05204_),
    .A2_N(_05244_),
    .B1(\design_top.MEM[7][25] ),
    .B2(_05246_),
    .X(_04099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08103_ (.A1_N(_05205_),
    .A2_N(_05244_),
    .B1(\design_top.MEM[7][24] ),
    .B2(_05246_),
    .X(_04098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08104_ (.A(_04875_),
    .B(_04958_),
    .X(_05248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08105_ (.A(_04908_),
    .B(_05248_),
    .X(_05249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08106_ (.A(_05249_),
    .X(_05250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _08107_ (.A(wbs_adr_i[0]),
    .B(_04880_),
    .C(_04964_),
    .Y(_05251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _08108_ (.A(_05251_),
    .B_N(_05249_),
    .Y(_05252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08109_ (.A(_05252_),
    .X(_05253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08110_ (.A1_N(_05166_),
    .A2_N(_05250_),
    .B1(\design_top.MEM[8][15] ),
    .B2(_05253_),
    .X(_04097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08111_ (.A1_N(_05174_),
    .A2_N(_05250_),
    .B1(\design_top.MEM[8][14] ),
    .B2(_05253_),
    .X(_04096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08112_ (.A1_N(_05175_),
    .A2_N(_05250_),
    .B1(\design_top.MEM[8][13] ),
    .B2(_05253_),
    .X(_04095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08113_ (.A1_N(_05176_),
    .A2_N(_05250_),
    .B1(\design_top.MEM[8][12] ),
    .B2(_05253_),
    .X(_04094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08114_ (.A1_N(_05177_),
    .A2_N(_05250_),
    .B1(\design_top.MEM[8][11] ),
    .B2(_05253_),
    .X(_04093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08115_ (.A1_N(_05178_),
    .A2_N(_05249_),
    .B1(\design_top.MEM[8][10] ),
    .B2(_05252_),
    .X(_04092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08116_ (.A1_N(_05179_),
    .A2_N(_05249_),
    .B1(\design_top.MEM[8][9] ),
    .B2(_05252_),
    .X(_04091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08117_ (.A1_N(_05180_),
    .A2_N(_05249_),
    .B1(\design_top.MEM[8][8] ),
    .B2(_05252_),
    .X(_04090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08118_ (.A(_04938_),
    .B(_05248_),
    .X(_05254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08119_ (.A(_05254_),
    .X(_05255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _08120_ (.A(_05251_),
    .B_N(_05254_),
    .Y(_05256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08121_ (.A(_05256_),
    .X(_05257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08122_ (.A1_N(_05181_),
    .A2_N(_05255_),
    .B1(\design_top.MEM[8][23] ),
    .B2(_05257_),
    .X(_04089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08123_ (.A1_N(_05186_),
    .A2_N(_05255_),
    .B1(\design_top.MEM[8][22] ),
    .B2(_05257_),
    .X(_04088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08124_ (.A1_N(_05187_),
    .A2_N(_05255_),
    .B1(\design_top.MEM[8][21] ),
    .B2(_05257_),
    .X(_04087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08125_ (.A1_N(_05188_),
    .A2_N(_05255_),
    .B1(\design_top.MEM[8][20] ),
    .B2(_05257_),
    .X(_04086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08126_ (.A1_N(_05189_),
    .A2_N(_05255_),
    .B1(\design_top.MEM[8][19] ),
    .B2(_05257_),
    .X(_04085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08127_ (.A1_N(_05190_),
    .A2_N(_05254_),
    .B1(\design_top.MEM[8][18] ),
    .B2(_05256_),
    .X(_04084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08128_ (.A1_N(_05191_),
    .A2_N(_05254_),
    .B1(\design_top.MEM[8][17] ),
    .B2(_05256_),
    .X(_04083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08129_ (.A1_N(_05192_),
    .A2_N(_05254_),
    .B1(\design_top.MEM[8][16] ),
    .B2(_05256_),
    .X(_04082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08130_ (.A(_05194_),
    .B(_05248_),
    .X(_05258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08131_ (.A(_05258_),
    .X(_05259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _08132_ (.A(_05251_),
    .B_N(_05258_),
    .Y(_05260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08133_ (.A(_05260_),
    .X(_05261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08134_ (.A1_N(_05193_),
    .A2_N(_05259_),
    .B1(\design_top.MEM[8][31] ),
    .B2(_05261_),
    .X(_04081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08135_ (.A1_N(_05199_),
    .A2_N(_05259_),
    .B1(\design_top.MEM[8][30] ),
    .B2(_05261_),
    .X(_04080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08136_ (.A1_N(_05200_),
    .A2_N(_05259_),
    .B1(\design_top.MEM[8][29] ),
    .B2(_05261_),
    .X(_04079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08137_ (.A1_N(_05201_),
    .A2_N(_05259_),
    .B1(\design_top.MEM[8][28] ),
    .B2(_05261_),
    .X(_04078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08138_ (.A1_N(_05202_),
    .A2_N(_05259_),
    .B1(\design_top.MEM[8][27] ),
    .B2(_05261_),
    .X(_04077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08139_ (.A1_N(_05203_),
    .A2_N(_05258_),
    .B1(\design_top.MEM[8][26] ),
    .B2(_05260_),
    .X(_04076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08140_ (.A1_N(_05204_),
    .A2_N(_05258_),
    .B1(\design_top.MEM[8][25] ),
    .B2(_05260_),
    .X(_04075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08141_ (.A1_N(_05205_),
    .A2_N(_05258_),
    .B1(\design_top.MEM[8][24] ),
    .B2(_05260_),
    .X(_04074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08142_ (.A(_04876_),
    .B(_04909_),
    .X(_05262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08143_ (.A(_05262_),
    .X(_05263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _08144_ (.A(_04886_),
    .B_N(_05262_),
    .Y(_05264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08145_ (.A(_05264_),
    .X(_05265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08146_ (.A1_N(_04903_),
    .A2_N(_05263_),
    .B1(\design_top.MEM[9][15] ),
    .B2(_05265_),
    .X(_04073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08147_ (.A1_N(_04918_),
    .A2_N(_05263_),
    .B1(\design_top.MEM[9][14] ),
    .B2(_05265_),
    .X(_04072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08148_ (.A1_N(_04920_),
    .A2_N(_05263_),
    .B1(\design_top.MEM[9][13] ),
    .B2(_05265_),
    .X(_04071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08149_ (.A1_N(_04922_),
    .A2_N(_05263_),
    .B1(\design_top.MEM[9][12] ),
    .B2(_05265_),
    .X(_04070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08150_ (.A1_N(_04924_),
    .A2_N(_05263_),
    .B1(\design_top.MEM[9][11] ),
    .B2(_05265_),
    .X(_04069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08151_ (.A1_N(_04926_),
    .A2_N(_05262_),
    .B1(\design_top.MEM[9][10] ),
    .B2(_05264_),
    .X(_04068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08152_ (.A1_N(_04928_),
    .A2_N(_05262_),
    .B1(\design_top.MEM[9][9] ),
    .B2(_05264_),
    .X(_04067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08153_ (.A1_N(_04930_),
    .A2_N(_05262_),
    .B1(\design_top.MEM[9][8] ),
    .B2(_05264_),
    .X(_04066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08154_ (.A(_04876_),
    .B(_04939_),
    .X(_05266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08155_ (.A(_05266_),
    .X(_05267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _08156_ (.A(_04886_),
    .B_N(_05266_),
    .Y(_05268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08157_ (.A(_05268_),
    .X(_05269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08158_ (.A1_N(_04936_),
    .A2_N(_05267_),
    .B1(\design_top.MEM[9][23] ),
    .B2(_05269_),
    .X(_04065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08159_ (.A1_N(_04944_),
    .A2_N(_05267_),
    .B1(\design_top.MEM[9][22] ),
    .B2(_05269_),
    .X(_04064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08160_ (.A1_N(_04946_),
    .A2_N(_05267_),
    .B1(\design_top.MEM[9][21] ),
    .B2(_05269_),
    .X(_04063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08161_ (.A1_N(_04948_),
    .A2_N(_05267_),
    .B1(\design_top.MEM[9][20] ),
    .B2(_05269_),
    .X(_04062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08162_ (.A1_N(_04950_),
    .A2_N(_05267_),
    .B1(\design_top.MEM[9][19] ),
    .B2(_05269_),
    .X(_04061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08163_ (.A1_N(_04952_),
    .A2_N(_05266_),
    .B1(\design_top.MEM[9][18] ),
    .B2(_05268_),
    .X(_04060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08164_ (.A1_N(_04954_),
    .A2_N(_05266_),
    .B1(\design_top.MEM[9][17] ),
    .B2(_05268_),
    .X(_04059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08165_ (.A1_N(_04956_),
    .A2_N(_05266_),
    .B1(\design_top.MEM[9][16] ),
    .B2(_05268_),
    .X(_04058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08166_ (.A(_04870_),
    .B(_05083_),
    .X(_05270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08167_ (.A(_05270_),
    .X(_05271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2b_2 _08168_ (.A(_05086_),
    .B_N(_05270_),
    .Y(_05272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08169_ (.A(_05272_),
    .X(_05273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08170_ (.A1_N(_04718_),
    .A2_N(_05271_),
    .B1(\design_top.MEM[13][31] ),
    .B2(_05273_),
    .X(_04057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08171_ (.A1_N(_04889_),
    .A2_N(_05271_),
    .B1(\design_top.MEM[13][30] ),
    .B2(_05273_),
    .X(_04056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08172_ (.A1_N(_04891_),
    .A2_N(_05271_),
    .B1(\design_top.MEM[13][29] ),
    .B2(_05273_),
    .X(_04055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08173_ (.A1_N(_04893_),
    .A2_N(_05271_),
    .B1(\design_top.MEM[13][28] ),
    .B2(_05273_),
    .X(_04054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08174_ (.A1_N(_04895_),
    .A2_N(_05271_),
    .B1(\design_top.MEM[13][27] ),
    .B2(_05273_),
    .X(_04053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08175_ (.A1_N(_04897_),
    .A2_N(_05270_),
    .B1(\design_top.MEM[13][26] ),
    .B2(_05272_),
    .X(_04052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08176_ (.A1_N(_04899_),
    .A2_N(_05270_),
    .B1(\design_top.MEM[13][25] ),
    .B2(_05272_),
    .X(_04051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08177_ (.A1_N(_04901_),
    .A2_N(_05270_),
    .B1(\design_top.MEM[13][24] ),
    .B2(_05272_),
    .X(_04050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _08178_ (.A1(_00326_),
    .A2(_04819_),
    .A3(_05013_),
    .B1(_04820_),
    .B2(_04822_),
    .X(_05274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08179_ (.A(_05014_),
    .B(_05274_),
    .X(_00548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _08180_ (.A(_04990_),
    .B(_00548_),
    .C(_05018_),
    .X(_05275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08181_ (.A(_05275_),
    .Y(_05276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08182_ (.A(_05276_),
    .X(_05277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08183_ (.A(_05277_),
    .X(_05278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08184_ (.A(_05275_),
    .X(_05279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08185_ (.A1(\design_top.IOMUX[3][31] ),
    .A2(_05278_),
    .B1(\design_top.DATAO[31] ),
    .B2(_05279_),
    .C1(_05063_),
    .X(_04049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08186_ (.A(_05277_),
    .X(_05280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08187_ (.A(_05275_),
    .X(_05281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08188_ (.A(_05281_),
    .X(_05282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08189_ (.A1(\design_top.IOMUX[3][30] ),
    .A2(_05280_),
    .B1(\design_top.DATAO[30] ),
    .B2(_05282_),
    .C1(_05063_),
    .X(_04048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08190_ (.A1(\design_top.IOMUX[3][29] ),
    .A2(_05280_),
    .B1(\design_top.DATAO[29] ),
    .B2(_05282_),
    .C1(_05063_),
    .X(_04047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08191_ (.A1(\design_top.IOMUX[3][28] ),
    .A2(_05280_),
    .B1(\design_top.DATAO[28] ),
    .B2(_05282_),
    .C1(_05063_),
    .X(_04046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08192_ (.A(_05062_),
    .X(_05283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08193_ (.A1(\design_top.IOMUX[3][27] ),
    .A2(_05280_),
    .B1(\design_top.DATAO[27] ),
    .B2(_05282_),
    .C1(_05283_),
    .X(_04045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08194_ (.A1(\design_top.IOMUX[3][26] ),
    .A2(_05280_),
    .B1(\design_top.DATAO[26] ),
    .B2(_05282_),
    .C1(_05283_),
    .X(_04044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08195_ (.A(_05277_),
    .X(_05284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08196_ (.A(_05281_),
    .X(_05285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08197_ (.A1(\design_top.IOMUX[3][25] ),
    .A2(_05284_),
    .B1(\design_top.DATAO[25] ),
    .B2(_05285_),
    .C1(_05283_),
    .X(_04043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08198_ (.A1(\design_top.IOMUX[3][24] ),
    .A2(_05284_),
    .B1(\design_top.DATAO[24] ),
    .B2(_05285_),
    .C1(_05283_),
    .X(_04042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08199_ (.A1(\design_top.IOMUX[3][23] ),
    .A2(_05284_),
    .B1(\design_top.DATAO[23] ),
    .B2(_05285_),
    .C1(_05283_),
    .X(_04041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08200_ (.A(_05062_),
    .X(_05286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08201_ (.A1(\design_top.IOMUX[3][22] ),
    .A2(_05284_),
    .B1(\design_top.DATAO[22] ),
    .B2(_05285_),
    .C1(_05286_),
    .X(_04040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08202_ (.A1(\design_top.IOMUX[3][21] ),
    .A2(_05284_),
    .B1(\design_top.DATAO[21] ),
    .B2(_05285_),
    .C1(_05286_),
    .X(_04039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08203_ (.A(_05276_),
    .X(_05287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08204_ (.A(_05281_),
    .X(_05288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08205_ (.A1(\design_top.IOMUX[3][20] ),
    .A2(_05287_),
    .B1(\design_top.DATAO[20] ),
    .B2(_05288_),
    .C1(_05286_),
    .X(_04038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08206_ (.A1(\design_top.IOMUX[3][19] ),
    .A2(_05287_),
    .B1(\design_top.DATAO[19] ),
    .B2(_05288_),
    .C1(_05286_),
    .X(_04037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08207_ (.A1(\design_top.IOMUX[3][18] ),
    .A2(_05287_),
    .B1(\design_top.DATAO[18] ),
    .B2(_05288_),
    .C1(_05286_),
    .X(_04036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08208_ (.A(_05022_),
    .X(_05289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08209_ (.A1(\design_top.IOMUX[3][17] ),
    .A2(_05287_),
    .B1(\design_top.DATAO[17] ),
    .B2(_05288_),
    .C1(_05289_),
    .X(_04035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08210_ (.A1(\design_top.IOMUX[3][16] ),
    .A2(_05287_),
    .B1(\design_top.DATAO[16] ),
    .B2(_05288_),
    .C1(_05289_),
    .X(_04034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08211_ (.A(_05276_),
    .X(_05290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08212_ (.A(_05275_),
    .X(_05291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08213_ (.A1(\design_top.IOMUX[3][15] ),
    .A2(_05290_),
    .B1(\design_top.DATAO[15] ),
    .B2(_05291_),
    .C1(_05289_),
    .X(_04033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08214_ (.A1(\design_top.IOMUX[3][14] ),
    .A2(_05290_),
    .B1(\design_top.DATAO[14] ),
    .B2(_05291_),
    .C1(_05289_),
    .X(_04032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08215_ (.A1(\design_top.IOMUX[3][13] ),
    .A2(_05290_),
    .B1(\design_top.DATAO[13] ),
    .B2(_05291_),
    .C1(_05289_),
    .X(_04031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08216_ (.A(_05022_),
    .X(_05292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08217_ (.A1(\design_top.IOMUX[3][12] ),
    .A2(_05290_),
    .B1(\design_top.DATAO[12] ),
    .B2(_05291_),
    .C1(_05292_),
    .X(_04030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08218_ (.A1(\design_top.IOMUX[3][11] ),
    .A2(_05290_),
    .B1(\design_top.DATAO[11] ),
    .B2(_05291_),
    .C1(_05292_),
    .X(_04029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08219_ (.A(_05276_),
    .X(_05293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08220_ (.A(_05275_),
    .X(_05294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08221_ (.A1(\design_top.IOMUX[3][10] ),
    .A2(_05293_),
    .B1(\design_top.DATAO[10] ),
    .B2(_05294_),
    .C1(_05292_),
    .X(_04028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08222_ (.A1(\design_top.IOMUX[3][9] ),
    .A2(_05293_),
    .B1(\design_top.DATAO[9] ),
    .B2(_05294_),
    .C1(_05292_),
    .X(_04027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08223_ (.A1(\design_top.IOMUX[3][8] ),
    .A2(_05293_),
    .B1(\design_top.DATAO[8] ),
    .B2(_05294_),
    .C1(_05292_),
    .X(_04026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08224_ (.A(_05022_),
    .X(_05295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08225_ (.A1(\design_top.IOMUX[3][7] ),
    .A2(_05293_),
    .B1(\design_top.DATAO[7] ),
    .B2(_05294_),
    .C1(_05295_),
    .X(_04025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08226_ (.A(\design_top.IRES[7] ),
    .X(_05296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08227_ (.A(_05296_),
    .X(_05297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a221o_2 _08228_ (.A1(\design_top.DATAO[6] ),
    .A2(_05278_),
    .B1(\design_top.IOMUX[3][6] ),
    .B2(_05279_),
    .C1(_05297_),
    .X(_04024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a221o_2 _08229_ (.A1(\design_top.DATAO[5] ),
    .A2(_05278_),
    .B1(\design_top.IOMUX[3][5] ),
    .B2(_05279_),
    .C1(_05297_),
    .X(_04023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08230_ (.A1(\design_top.IOMUX[3][4] ),
    .A2(_05293_),
    .B1(\design_top.DATAO[4] ),
    .B2(_05294_),
    .C1(_05295_),
    .X(_04022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08231_ (.A1(\design_top.IOMUX[3][3] ),
    .A2(_05277_),
    .B1(\design_top.DATAO[3] ),
    .B2(_05281_),
    .C1(_05295_),
    .X(_04021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08232_ (.A1(\design_top.IOMUX[3][2] ),
    .A2(_05277_),
    .B1(\design_top.DATAO[2] ),
    .B2(_05281_),
    .C1(_05295_),
    .X(_04020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a221o_2 _08233_ (.A1(\design_top.DATAO[1] ),
    .A2(_05278_),
    .B1(\design_top.IOMUX[3][1] ),
    .B2(_05279_),
    .C1(_05296_),
    .X(_04019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a221o_2 _08234_ (.A1(\design_top.DATAO[0] ),
    .A2(_05278_),
    .B1(\design_top.IOMUX[3][0] ),
    .B2(_05279_),
    .C1(_05296_),
    .X(_04018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08235_ (.A(\design_top.core0.XRES ),
    .X(_05298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08236_ (.A(_05298_),
    .X(_05299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08237_ (.A(\design_top.IDATA[31] ),
    .Y(_05300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08238_ (.A(_04619_),
    .X(_05301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08239_ (.A(_05301_),
    .X(_05302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08240_ (.A(_00904_),
    .Y(_05303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _08241_ (.A(_00905_),
    .B(_05303_),
    .C(_00906_),
    .X(_05304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _08242_ (.A(io_out[21]),
    .B(io_out[20]),
    .Y(_05305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _08243_ (.A(io_out[23]),
    .B(_05305_),
    .C_N(io_out[22]),
    .X(_05306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08244_ (.A(_05304_),
    .B(_05306_),
    .Y(_05307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08245_ (.A(_00905_),
    .Y(_05308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _08246_ (.A(_05308_),
    .B(_05303_),
    .C(_00906_),
    .X(_05309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08247_ (.A(_05306_),
    .B(_05309_),
    .Y(_05310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08248_ (.A(_05307_),
    .B(_05310_),
    .X(_05311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08249_ (.A(_05311_),
    .Y(_05312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08250_ (.A(_05312_),
    .X(_01240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08251_ (.A(\design_top.core0.UIMM[31] ),
    .Y(_05313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08252_ (.A(_04618_),
    .X(_05314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08253_ (.A(_05314_),
    .X(_05315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08254_ (.A(_05315_),
    .X(_05316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _08255_ (.A1(_05300_),
    .A2(_05302_),
    .A3(_01240_),
    .B1(_05313_),
    .B2(_05316_),
    .X(_05317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08256_ (.A(_05299_),
    .B(_05317_),
    .Y(_04017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08257_ (.A(_04620_),
    .X(_05318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08258_ (.A(_05318_),
    .X(_05319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08259_ (.A(_05319_),
    .X(\design_top.HLT ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08260_ (.A(\design_top.IDATA[30] ),
    .Y(_05320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08261_ (.A(\design_top.core0.UIMM[30] ),
    .Y(_05321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08262_ (.A(_05315_),
    .X(_05322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _08263_ (.A1(_05320_),
    .A2(_05302_),
    .A3(_01240_),
    .B1(_05321_),
    .B2(_05322_),
    .X(_05323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08264_ (.A(_05299_),
    .B(_05323_),
    .Y(_04016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08265_ (.A(_05318_),
    .X(_05324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08266_ (.A(_01298_),
    .Y(_05325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08267_ (.A(_04619_),
    .B(_05312_),
    .X(_05326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08268_ (.A(_05326_),
    .X(_05327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _08269_ (.A1_N(\design_top.core0.UIMM[29] ),
    .A2_N(_05324_),
    .B1(_05325_),
    .B2(_05327_),
    .X(_05328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08270_ (.A(_05299_),
    .B(_05328_),
    .Y(_04015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08271_ (.A(_01294_),
    .Y(_05329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _08272_ (.A1_N(\design_top.core0.UIMM[28] ),
    .A2_N(_05324_),
    .B1(_05329_),
    .B2(_05327_),
    .X(_05330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08273_ (.A(_05299_),
    .B(_05330_),
    .Y(_04014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08274_ (.A(_01290_),
    .Y(_05331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _08275_ (.A1_N(\design_top.core0.UIMM[27] ),
    .A2_N(_05324_),
    .B1(_05331_),
    .B2(_05327_),
    .X(_05332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08276_ (.A(_05299_),
    .B(_05332_),
    .Y(_04013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08277_ (.A(_05298_),
    .X(_05333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08278_ (.A(_04620_),
    .X(_05334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08279_ (.A(_05334_),
    .X(_05335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08280_ (.A(_01286_),
    .Y(_05336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _08281_ (.A1_N(\design_top.core0.UIMM[26] ),
    .A2_N(_05335_),
    .B1(_05336_),
    .B2(_05327_),
    .X(_05337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08282_ (.A(_05333_),
    .B(_05337_),
    .Y(_04012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08283_ (.A(_01282_),
    .Y(_05338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _08284_ (.A1_N(\design_top.core0.UIMM[25] ),
    .A2_N(_05335_),
    .B1(_05338_),
    .B2(_05327_),
    .X(_05339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08285_ (.A(_05333_),
    .B(_05339_),
    .Y(_04011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08286_ (.A(_01278_),
    .Y(_05340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _08287_ (.A1_N(\design_top.core0.UIMM[24] ),
    .A2_N(_05335_),
    .B1(_05340_),
    .B2(_05326_),
    .X(_05341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08288_ (.A(_05333_),
    .B(_05341_),
    .Y(_04010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08289_ (.A(\design_top.IDATA[23] ),
    .Y(_05342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08290_ (.A(\design_top.core0.UIMM[23] ),
    .Y(_05343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _08291_ (.A1(_05342_),
    .A2(_05302_),
    .A3(_01240_),
    .B1(_05343_),
    .B2(_05322_),
    .X(_05344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08292_ (.A(_05333_),
    .B(_05344_),
    .Y(_04009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08293_ (.A(\design_top.IDATA[22] ),
    .Y(_05345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08294_ (.A(_05301_),
    .X(_05346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08295_ (.A(\design_top.core0.UIMM[22] ),
    .Y(_05347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _08296_ (.A1(_05345_),
    .A2(_05346_),
    .A3(_05312_),
    .B1(_05347_),
    .B2(_05322_),
    .X(_05348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08297_ (.A(_05333_),
    .B(_05348_),
    .Y(_04008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08298_ (.A(_05298_),
    .X(_05349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08299_ (.A(\design_top.IDATA[21] ),
    .Y(_05350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08300_ (.A(\design_top.core0.UIMM[21] ),
    .Y(_05351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _08301_ (.A1(_05350_),
    .A2(_05346_),
    .A3(_05312_),
    .B1(_05351_),
    .B2(_05322_),
    .X(_05352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08302_ (.A(_05349_),
    .B(_05352_),
    .Y(_04007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08303_ (.A(_01358_),
    .Y(_05353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _08304_ (.A(io_out[23]),
    .B(io_out[22]),
    .C(_05305_),
    .X(_05354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31ai_2 _08305_ (.A1(_05308_),
    .A2(_00904_),
    .A3(_05354_),
    .B1(_05314_),
    .Y(_05355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08306_ (.A(_05355_),
    .X(_05356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _08307_ (.A1_N(\design_top.core0.UIMM[20] ),
    .A2_N(_05335_),
    .B1(_05353_),
    .B2(_05356_),
    .X(_05357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08308_ (.A(_05349_),
    .B(_05357_),
    .Y(_04006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08309_ (.A(_01356_),
    .Y(_05358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _08310_ (.A1_N(\design_top.core0.UIMM[19] ),
    .A2_N(_05335_),
    .B1(_05358_),
    .B2(_05356_),
    .X(_05359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08311_ (.A(_05349_),
    .B(_05359_),
    .Y(_04005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08312_ (.A(_05334_),
    .X(_05360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08313_ (.A(_01354_),
    .Y(_05361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _08314_ (.A1_N(\design_top.core0.UIMM[18] ),
    .A2_N(_05360_),
    .B1(_05361_),
    .B2(_05356_),
    .X(_05362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08315_ (.A(_05349_),
    .B(_05362_),
    .Y(_04004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08316_ (.A(_01352_),
    .Y(_05363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _08317_ (.A1_N(\design_top.core0.UIMM[17] ),
    .A2_N(_05360_),
    .B1(_05363_),
    .B2(_05356_),
    .X(_05364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08318_ (.A(_05349_),
    .B(_05364_),
    .Y(_04003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08319_ (.A(_05298_),
    .X(_05365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08320_ (.A(_01350_),
    .Y(_05366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _08321_ (.A1_N(\design_top.core0.UIMM[16] ),
    .A2_N(_05360_),
    .B1(_05366_),
    .B2(_05356_),
    .X(_05367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08322_ (.A(_05365_),
    .B(_05367_),
    .Y(_04002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08323_ (.A(_01348_),
    .Y(_05368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _08324_ (.A1_N(\design_top.core0.UIMM[15] ),
    .A2_N(_05360_),
    .B1(_05368_),
    .B2(_05355_),
    .X(_05369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08325_ (.A(_05365_),
    .B(_05369_),
    .Y(_04001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08326_ (.A(_01346_),
    .Y(_05370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _08327_ (.A1_N(\design_top.core0.UIMM[14] ),
    .A2_N(_05360_),
    .B1(_05370_),
    .B2(_05355_),
    .X(_05371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08328_ (.A(_05365_),
    .B(_05371_),
    .Y(_04000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08329_ (.A(_01344_),
    .Y(_05372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _08330_ (.A1_N(\design_top.core0.UIMM[13] ),
    .A2_N(_05319_),
    .B1(_05372_),
    .B2(_05355_),
    .X(_05373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08331_ (.A(_05365_),
    .B(_05373_),
    .Y(_03999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08332_ (.A(_01342_),
    .Y(_05374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08333_ (.A(_00906_),
    .Y(_05375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and4b_2 _08334_ (.A_N(_05354_),
    .B(_05303_),
    .C(_05375_),
    .D(_00905_),
    .X(_00010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08335_ (.A(_04620_),
    .B(_00010_),
    .X(_05376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _08336_ (.A1_N(\design_top.core0.UIMM[12] ),
    .A2_N(_05319_),
    .B1(_05374_),
    .B2(_05376_),
    .X(_05377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08337_ (.A(_05365_),
    .B(_05377_),
    .Y(_03998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08338_ (.A(_05346_),
    .X(_05378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08339_ (.A(_05315_),
    .X(_05379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08340_ (.A(_04716_),
    .X(_05380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08341_ (.A(_05380_),
    .X(_05381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08342_ (.A1(_00049_),
    .A2(_05378_),
    .B1(_04799_),
    .B2(_05379_),
    .C1(_05381_),
    .X(_03997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08343_ (.A1(_00048_),
    .A2(_05378_),
    .B1(\design_top.core0.SIMM[10] ),
    .B2(_05379_),
    .C1(_05381_),
    .X(_03996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08344_ (.A(\design_top.core0.SIMM[9] ),
    .X(_05382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08345_ (.A(_05314_),
    .X(_05383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08346_ (.A(_05383_),
    .X(_05384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08347_ (.A(_05384_),
    .X(_05385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08348_ (.A1(_00077_),
    .A2(_05378_),
    .B1(_05382_),
    .B2(_05385_),
    .C1(_05381_),
    .X(_03995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08349_ (.A(\design_top.core0.SIMM[8] ),
    .X(_05386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08350_ (.A1(_00076_),
    .A2(_05378_),
    .B1(_05386_),
    .B2(_05385_),
    .C1(_05381_),
    .X(_03994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08351_ (.A(_05346_),
    .X(_05387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08352_ (.A(\design_top.core0.SIMM[7] ),
    .X(_05388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08353_ (.A1(_00075_),
    .A2(_05387_),
    .B1(_05388_),
    .B2(_05385_),
    .C1(_05381_),
    .X(_03993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08354_ (.A(\design_top.core0.SIMM[6] ),
    .X(_05389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08355_ (.A(_05380_),
    .X(_05390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08356_ (.A1(_00074_),
    .A2(_05387_),
    .B1(_05389_),
    .B2(_05385_),
    .C1(_05390_),
    .X(_03992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08357_ (.A(\design_top.core0.SIMM[5] ),
    .X(_05391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08358_ (.A1(_00073_),
    .A2(_05387_),
    .B1(_05391_),
    .B2(_05385_),
    .C1(_05390_),
    .X(_03991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08359_ (.A(\design_top.core0.SIMM[4] ),
    .X(_05392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08360_ (.A(_05384_),
    .X(_05393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08361_ (.A1(_00072_),
    .A2(_05387_),
    .B1(_05392_),
    .B2(_05393_),
    .C1(_05390_),
    .X(_03990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08362_ (.A1(_00071_),
    .A2(_05387_),
    .B1(_04811_),
    .B2(_05393_),
    .C1(_05390_),
    .X(_03989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08363_ (.A(_05301_),
    .X(_05394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08364_ (.A(_05394_),
    .X(_05395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08365_ (.A1(_00069_),
    .A2(_05395_),
    .B1(_04814_),
    .B2(_05393_),
    .C1(_05390_),
    .X(_03988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08366_ (.A(_05380_),
    .X(_05396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08367_ (.A1(_00058_),
    .A2(_05395_),
    .B1(_04817_),
    .B2(_05393_),
    .C1(_05396_),
    .X(_03987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08368_ (.A1(_00047_),
    .A2(_05395_),
    .B1(\design_top.core0.SIMM[0] ),
    .B2(_05393_),
    .C1(_05396_),
    .X(_03986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08369_ (.A(_05298_),
    .X(_05397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08370_ (.A1(_05300_),
    .A2(_05319_),
    .B1(_01360_),
    .B2(_05316_),
    .X(_05398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08371_ (.A(_05397_),
    .B(_05398_),
    .Y(_03985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08372_ (.A(_05384_),
    .X(_05399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08373_ (.A1(_00070_),
    .A2(_05395_),
    .B1(\design_top.core0.SIMM[30] ),
    .B2(_05399_),
    .C1(_05396_),
    .X(_03984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08374_ (.A1(_00068_),
    .A2(_05395_),
    .B1(_04724_),
    .B2(_05399_),
    .C1(_05396_),
    .X(_03983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08375_ (.A(_05394_),
    .X(_05400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08376_ (.A1(_00067_),
    .A2(_05400_),
    .B1(_04729_),
    .B2(_05399_),
    .C1(_05396_),
    .X(_03982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08377_ (.A(_05380_),
    .X(_05401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08378_ (.A1(_00066_),
    .A2(_05400_),
    .B1(\design_top.core0.SIMM[27] ),
    .B2(_05399_),
    .C1(_05401_),
    .X(_03981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08379_ (.A1(_00065_),
    .A2(_05400_),
    .B1(\design_top.core0.SIMM[26] ),
    .B2(_05399_),
    .C1(_05401_),
    .X(_03980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08380_ (.A(\design_top.core0.SIMM[25] ),
    .X(_05402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08381_ (.A(_05314_),
    .X(_05403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08382_ (.A(_05403_),
    .X(_05404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08383_ (.A1(_00064_),
    .A2(_05400_),
    .B1(_05402_),
    .B2(_05404_),
    .C1(_05401_),
    .X(_03979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08384_ (.A(\design_top.core0.SIMM[24] ),
    .X(_05405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08385_ (.A1(_00063_),
    .A2(_05400_),
    .B1(_05405_),
    .B2(_05404_),
    .C1(_05401_),
    .X(_03978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08386_ (.A(_05394_),
    .X(_05406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08387_ (.A1(_00062_),
    .A2(_05406_),
    .B1(_04846_),
    .B2(_05404_),
    .C1(_05401_),
    .X(_03977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08388_ (.A(_05380_),
    .X(_05407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08389_ (.A1(_00061_),
    .A2(_05406_),
    .B1(_04769_),
    .B2(_05404_),
    .C1(_05407_),
    .X(_03976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08390_ (.A(\design_top.core0.SIMM[21] ),
    .X(_05408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08391_ (.A1(_00060_),
    .A2(_05406_),
    .B1(_05408_),
    .B2(_05404_),
    .C1(_05407_),
    .X(_03975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08392_ (.A(_05403_),
    .X(_05409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08393_ (.A1(_00059_),
    .A2(_05406_),
    .B1(_04765_),
    .B2(_05409_),
    .C1(_05407_),
    .X(_03974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08394_ (.A1(_00057_),
    .A2(_05406_),
    .B1(_04753_),
    .B2(_05409_),
    .C1(_05407_),
    .X(_03973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08395_ (.A(_05394_),
    .X(_05410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08396_ (.A1(_00056_),
    .A2(_05410_),
    .B1(_04751_),
    .B2(_05409_),
    .C1(_05407_),
    .X(_03972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08397_ (.A(\design_top.core0.SIMM[17] ),
    .X(_05411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08398_ (.A(_04716_),
    .X(_05412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08399_ (.A(_05412_),
    .X(_05413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08400_ (.A1(_00055_),
    .A2(_05410_),
    .B1(_05411_),
    .B2(_05409_),
    .C1(_05413_),
    .X(_03971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08401_ (.A(\design_top.core0.SIMM[16] ),
    .X(_05414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08402_ (.A1(_00054_),
    .A2(_05410_),
    .B1(_05414_),
    .B2(_05409_),
    .C1(_05413_),
    .X(_03970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08403_ (.A(_05403_),
    .X(_05415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08404_ (.A1(_00053_),
    .A2(_05410_),
    .B1(_04841_),
    .B2(_05415_),
    .C1(_05413_),
    .X(_03969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08405_ (.A1(_00052_),
    .A2(_05410_),
    .B1(_04776_),
    .B2(_05415_),
    .C1(_05413_),
    .X(_03968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08406_ (.A(_05394_),
    .X(_05416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08407_ (.A(\design_top.core0.SIMM[13] ),
    .X(_05417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08408_ (.A1(_00051_),
    .A2(_05416_),
    .B1(_05417_),
    .B2(_05415_),
    .C1(_05413_),
    .X(_03967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08409_ (.A(_05412_),
    .X(_05418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08410_ (.A1(_00050_),
    .A2(_05416_),
    .B1(_04786_),
    .B2(_05415_),
    .C1(_05418_),
    .X(_03966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08411_ (.A(_05301_),
    .X(_05419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08412_ (.A(_05354_),
    .X(_05420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08413_ (.A(\design_top.core0.XRCC ),
    .Y(_05421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _08414_ (.A1(_05419_),
    .A2(_05420_),
    .A3(_05309_),
    .B1(_05421_),
    .B2(_05322_),
    .X(_05422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08415_ (.A(_05397_),
    .B(_05422_),
    .Y(_03965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08416_ (.A(\design_top.core0.XMCC ),
    .Y(_05423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08417_ (.A(_05383_),
    .X(_05424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _08418_ (.A1(_05419_),
    .A2(_05420_),
    .A3(_05304_),
    .B1(_05423_),
    .B2(_05424_),
    .X(_05425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08419_ (.A(_05397_),
    .B(_05425_),
    .Y(_03964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08420_ (.A(_04716_),
    .X(_05426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _08421_ (.A1(\design_top.core0.XSCC ),
    .A2(_05379_),
    .B1(_05426_),
    .C1(_05376_),
    .X(_03963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and4b_2 _08422_ (.A_N(_05420_),
    .B(_05375_),
    .C(_05308_),
    .D(_05303_),
    .X(_05427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08423_ (.A(_05426_),
    .X(_05428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _08424_ (.A1(\design_top.HLT ),
    .A2(_05427_),
    .B1(_05428_),
    .X(_03962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _08425_ (.A(_05308_),
    .B(_00904_),
    .C(_05375_),
    .X(_05429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08426_ (.A(\design_top.core0.XBCC ),
    .Y(_05430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _08427_ (.A1(_05419_),
    .A2(_05420_),
    .A3(_05429_),
    .B1(_05430_),
    .B2(_05424_),
    .X(_05431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08428_ (.A(_05397_),
    .B(_05431_),
    .Y(_03961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08429_ (.A(_05420_),
    .B(_05429_),
    .Y(_00009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _08430_ (.A1(_05419_),
    .A2(_05429_),
    .A3(_05306_),
    .B1(_04621_),
    .B2(_05424_),
    .X(_05432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08431_ (.A(_05397_),
    .B(_05432_),
    .Y(_03960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08432_ (.A(_05315_),
    .X(_05433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08433_ (.A(_05346_),
    .X(_05434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and4bb_2 _08434_ (.A_N(_05429_),
    .B_N(_05305_),
    .C(io_out[23]),
    .D(io_out[22]),
    .X(_00008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08435_ (.A1(\design_top.core0.XJAL ),
    .A2(_05433_),
    .B1(_05434_),
    .B2(_00008_),
    .C1(_05418_),
    .X(_03959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08436_ (.A1(\design_top.core0.XAUIPC ),
    .A2(_05433_),
    .B1(_05434_),
    .B2(_05307_),
    .C1(_05418_),
    .X(_03958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08437_ (.A1(\design_top.core0.XLUI ),
    .A2(_05433_),
    .B1(_05378_),
    .B2(_05310_),
    .C1(_05418_),
    .X(_03957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08438_ (.A(\design_top.core0.XRES ),
    .X(_05435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08439_ (.A(\design_top.core0.FCT7[5] ),
    .Y(_05436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08440_ (.A1(_05320_),
    .A2(_05319_),
    .B1(_05436_),
    .B2(_05316_),
    .X(_05437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08441_ (.A(_05435_),
    .B(_05437_),
    .Y(_03956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08442_ (.A(_05334_),
    .X(_05438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22oi_2 _08443_ (.A1(\design_top.IDATA[23] ),
    .A2(_05433_),
    .B1(\design_top.core0.S2PTR[3] ),
    .B2(_05438_),
    .Y(_05439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08444_ (.A(_05435_),
    .B(_05439_),
    .Y(_03955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22oi_2 _08445_ (.A1(\design_top.IDATA[22] ),
    .A2(_05316_),
    .B1(\design_top.core0.S2PTR[2] ),
    .B2(_05324_),
    .Y(_05440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08446_ (.A(_05435_),
    .B(_05440_),
    .Y(_03954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22oi_2 _08447_ (.A1(\design_top.IDATA[21] ),
    .A2(_05316_),
    .B1(\design_top.core0.S2PTR[1] ),
    .B2(_05324_),
    .Y(_05441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08448_ (.A(_05435_),
    .B(_05441_),
    .Y(_03953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08449_ (.A1(\design_top.IDATA[20] ),
    .A2(_05416_),
    .B1(\design_top.core0.S2PTR[0] ),
    .B2(_05415_),
    .C1(_05418_),
    .X(_03952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08450_ (.A(_05403_),
    .X(_05442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08451_ (.A(_05412_),
    .X(_05443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08452_ (.A1(\design_top.IDATA[18] ),
    .A2(_05416_),
    .B1(\design_top.core0.S1PTR[3] ),
    .B2(_05442_),
    .C1(_05443_),
    .X(_03951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08453_ (.A1(\design_top.IDATA[17] ),
    .A2(_05416_),
    .B1(\design_top.core0.S1PTR[2] ),
    .B2(_05442_),
    .C1(_05443_),
    .X(_03950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08454_ (.A(_05301_),
    .X(_05444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08455_ (.A(_05444_),
    .X(_05445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08456_ (.A1(\design_top.IDATA[16] ),
    .A2(_05445_),
    .B1(\design_top.core0.S1PTR[1] ),
    .B2(_05442_),
    .C1(_05443_),
    .X(_03949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08457_ (.A1(\design_top.IDATA[15] ),
    .A2(_05445_),
    .B1(\design_top.core0.S1PTR[0] ),
    .B2(_05442_),
    .C1(_05443_),
    .X(_03948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08458_ (.A1(\design_top.IDATA[14] ),
    .A2(_05445_),
    .B1(\design_top.core0.FCT3[2] ),
    .B2(_05442_),
    .C1(_05443_),
    .X(_03947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08459_ (.A(\design_top.core0.FCT3[1] ),
    .X(_05446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08460_ (.A(_05403_),
    .X(_05447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08461_ (.A(_05412_),
    .X(_05448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08462_ (.A1(\design_top.IDATA[13] ),
    .A2(_05445_),
    .B1(_05446_),
    .B2(_05447_),
    .C1(_05448_),
    .X(_03946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08463_ (.A1(\design_top.IDATA[12] ),
    .A2(_05445_),
    .B1(\design_top.core0.FCT3[0] ),
    .B2(_05447_),
    .C1(_05448_),
    .X(_03945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08464_ (.A(_05444_),
    .X(_05449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08465_ (.A1(\design_top.IDATA[10] ),
    .A2(_05449_),
    .B1(\design_top.core0.XIDATA[10] ),
    .B2(_05447_),
    .C1(_05448_),
    .X(_03944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08466_ (.A1(\design_top.IDATA[9] ),
    .A2(_05449_),
    .B1(\design_top.core0.XIDATA[9] ),
    .B2(_05447_),
    .C1(_05448_),
    .X(_03943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08467_ (.A1(\design_top.IDATA[8] ),
    .A2(_05449_),
    .B1(\design_top.core0.XIDATA[8] ),
    .B2(_05447_),
    .C1(_05448_),
    .X(_03942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08468_ (.A(_05314_),
    .X(_05450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08469_ (.A(_05450_),
    .X(_05451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08470_ (.A(_05412_),
    .X(_05452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08471_ (.A1(\design_top.IDATA[7] ),
    .A2(_05449_),
    .B1(\design_top.core0.XIDATA[7] ),
    .B2(_05451_),
    .C1(_05452_),
    .X(_03941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08472_ (.A1(_00101_),
    .A2(_05449_),
    .B1(\design_top.IADDR[31] ),
    .B2(_05451_),
    .C1(_05452_),
    .X(_03940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08473_ (.A(_05444_),
    .X(_05453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08474_ (.A1(_00100_),
    .A2(_05453_),
    .B1(\design_top.IADDR[30] ),
    .B2(_05451_),
    .C1(_05452_),
    .X(_03939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08475_ (.A1(_00098_),
    .A2(_05453_),
    .B1(\design_top.IADDR[29] ),
    .B2(_05451_),
    .C1(_05452_),
    .X(_03938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08476_ (.A1(_00097_),
    .A2(_05453_),
    .B1(\design_top.IADDR[28] ),
    .B2(_05451_),
    .C1(_05452_),
    .X(_03937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08477_ (.A(_05450_),
    .X(_05454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08478_ (.A(_04716_),
    .X(_05455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08479_ (.A(_05455_),
    .X(_05456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08480_ (.A1(_00096_),
    .A2(_05453_),
    .B1(\design_top.IADDR[27] ),
    .B2(_05454_),
    .C1(_05456_),
    .X(_03936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08481_ (.A1(_00095_),
    .A2(_05453_),
    .B1(\design_top.IADDR[26] ),
    .B2(_05454_),
    .C1(_05456_),
    .X(_03935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08482_ (.A(_05444_),
    .X(_05457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08483_ (.A1(_00094_),
    .A2(_05457_),
    .B1(\design_top.IADDR[25] ),
    .B2(_05454_),
    .C1(_05456_),
    .X(_03934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08484_ (.A1(_00093_),
    .A2(_05457_),
    .B1(\design_top.IADDR[24] ),
    .B2(_05454_),
    .C1(_05456_),
    .X(_03933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08485_ (.A1(_00092_),
    .A2(_05457_),
    .B1(\design_top.IADDR[23] ),
    .B2(_05454_),
    .C1(_05456_),
    .X(_03932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08486_ (.A(_05450_),
    .X(_05458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08487_ (.A(_05455_),
    .X(_05459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08488_ (.A1(_00091_),
    .A2(_05457_),
    .B1(\design_top.IADDR[22] ),
    .B2(_05458_),
    .C1(_05459_),
    .X(_03931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08489_ (.A1(_00090_),
    .A2(_05457_),
    .B1(\design_top.IADDR[21] ),
    .B2(_05458_),
    .C1(_05459_),
    .X(_03930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08490_ (.A(_05444_),
    .X(_05460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08491_ (.A1(_00089_),
    .A2(_05460_),
    .B1(\design_top.IADDR[20] ),
    .B2(_05458_),
    .C1(_05459_),
    .X(_03929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08492_ (.A1(_00088_),
    .A2(_05460_),
    .B1(\design_top.IADDR[19] ),
    .B2(_05458_),
    .C1(_05459_),
    .X(_03928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08493_ (.A1(_00087_),
    .A2(_05460_),
    .B1(\design_top.IADDR[18] ),
    .B2(_05458_),
    .C1(_05459_),
    .X(_03927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08494_ (.A(_05450_),
    .X(_05461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08495_ (.A(_05455_),
    .X(_05462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08496_ (.A1(_00086_),
    .A2(_05460_),
    .B1(\design_top.IADDR[17] ),
    .B2(_05461_),
    .C1(_05462_),
    .X(_03926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08497_ (.A1(_00085_),
    .A2(_05460_),
    .B1(\design_top.IADDR[16] ),
    .B2(_05461_),
    .C1(_05462_),
    .X(_03925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08498_ (.A(_05334_),
    .X(_05463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08499_ (.A1(_00084_),
    .A2(_05463_),
    .B1(\design_top.IADDR[15] ),
    .B2(_05461_),
    .C1(_05462_),
    .X(_03924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08500_ (.A1(_00083_),
    .A2(_05463_),
    .B1(\design_top.IADDR[14] ),
    .B2(_05461_),
    .C1(_05462_),
    .X(_03923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08501_ (.A1(_00082_),
    .A2(_05463_),
    .B1(\design_top.IADDR[13] ),
    .B2(_05461_),
    .C1(_05462_),
    .X(_03922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08502_ (.A(_05450_),
    .X(_05464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08503_ (.A(_05455_),
    .X(_05465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08504_ (.A1(_00081_),
    .A2(_05463_),
    .B1(\design_top.IADDR[12] ),
    .B2(_05464_),
    .C1(_05465_),
    .X(_03921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08505_ (.A1(_00080_),
    .A2(_05463_),
    .B1(\design_top.IADDR[11] ),
    .B2(_05464_),
    .C1(_05465_),
    .X(_03920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08506_ (.A(_05334_),
    .X(_05466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08507_ (.A1(_00079_),
    .A2(_05466_),
    .B1(\design_top.IADDR[10] ),
    .B2(_05464_),
    .C1(_05465_),
    .X(_03919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08508_ (.A1(_00108_),
    .A2(_05466_),
    .B1(\design_top.IADDR[9] ),
    .B2(_05464_),
    .C1(_05465_),
    .X(_03918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08509_ (.A1(_00107_),
    .A2(_05466_),
    .B1(\design_top.IADDR[8] ),
    .B2(_05464_),
    .C1(_05465_),
    .X(_03917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08510_ (.A(_05315_),
    .X(_05467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08511_ (.A(_05455_),
    .X(_05468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08512_ (.A1(_00106_),
    .A2(_05466_),
    .B1(\design_top.IADDR[7] ),
    .B2(_05467_),
    .C1(_05468_),
    .X(_03916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08513_ (.A1(_00105_),
    .A2(_05466_),
    .B1(\design_top.IADDR[6] ),
    .B2(_05467_),
    .C1(_05468_),
    .X(_03915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08514_ (.A1(_00104_),
    .A2(_05438_),
    .B1(\design_top.IADDR[5] ),
    .B2(_05467_),
    .C1(_05468_),
    .X(_03914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08515_ (.A(\design_top.IADDR[4] ),
    .X(_05469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08516_ (.A1(_00103_),
    .A2(_05438_),
    .B1(_05469_),
    .B2(_05467_),
    .C1(_05468_),
    .X(_03913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08517_ (.A1(_00102_),
    .A2(_05438_),
    .B1(io_out[19]),
    .B2(_05467_),
    .C1(_05468_),
    .X(_03912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08518_ (.A1(_00099_),
    .A2(_05438_),
    .B1(io_out[18]),
    .B2(_05433_),
    .C1(_05426_),
    .X(_03911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08519_ (.A(_05424_),
    .X(_05470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _08520_ (.A1(_00011_),
    .A2(_05470_),
    .B1(_05435_),
    .X(_03910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _08521_ (.A(_05426_),
    .B(\design_top.core0.FLUSH[1] ),
    .C(_04616_),
    .X(_03909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _08522_ (.A(_05428_),
    .B(_00007_),
    .X(_03908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _08523_ (.A(_05428_),
    .B(_00006_),
    .X(_03907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _08524_ (.A(_05428_),
    .B(_00005_),
    .X(_03906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _08525_ (.A(_05428_),
    .B(_00004_),
    .X(_03905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08526_ (.A(\design_top.uart0.UART_RBAUD[1] ),
    .B(\design_top.uart0.UART_RBAUD[0] ),
    .X(_05471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _08527_ (.A(\design_top.uart0.UART_RBAUD[2] ),
    .B(_05471_),
    .C(\design_top.uart0.UART_RBAUD[3] ),
    .X(_05472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08528_ (.A(\design_top.uart0.UART_RBAUD[4] ),
    .B(_05472_),
    .X(_05473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08529_ (.A(\design_top.uart0.UART_RBAUD[5] ),
    .B(_05473_),
    .X(_05474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08530_ (.A(\design_top.uart0.UART_RBAUD[6] ),
    .B(_05474_),
    .X(_05475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08531_ (.A(\design_top.uart0.UART_RBAUD[7] ),
    .B(_05475_),
    .X(_05476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08532_ (.A(\design_top.uart0.UART_RBAUD[8] ),
    .B(_05476_),
    .X(_05477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08533_ (.A(\design_top.uart0.UART_RBAUD[9] ),
    .B(_05477_),
    .X(_05478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08534_ (.A(\design_top.uart0.UART_RBAUD[10] ),
    .B(_05478_),
    .X(_05479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08535_ (.A(\design_top.uart0.UART_RBAUD[11] ),
    .B(_05479_),
    .X(_05480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08536_ (.A(\design_top.uart0.UART_RBAUD[12] ),
    .B(_05480_),
    .X(_05481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08537_ (.A(\design_top.uart0.UART_RBAUD[13] ),
    .B(_05481_),
    .X(_05482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _08538_ (.A(\design_top.uart0.UART_RBAUD[14] ),
    .B(_05482_),
    .C(\design_top.uart0.UART_RBAUD[15] ),
    .X(_00926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08539_ (.A(_00926_),
    .Y(_05483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08540_ (.A(\design_top.uart0.UART_RSTATE[1] ),
    .Y(_05484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08541_ (.A(\design_top.uart0.UART_RSTATE[2] ),
    .Y(_05485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08542_ (.A(_05484_),
    .B(\design_top.uart0.UART_RSTATE[0] ),
    .C(\design_top.uart0.UART_RSTATE[3] ),
    .D(_05485_),
    .X(_05486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08543_ (.A(_05486_),
    .Y(_00344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08544_ (.A(_05483_),
    .B(_00344_),
    .X(_05487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08545_ (.A(_05487_),
    .Y(_05488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _08546_ (.A1(\design_top.uart0.UART_RBAUD[14] ),
    .A2(_05482_),
    .B1(\design_top.uart0.UART_RBAUD[15] ),
    .C1(_05488_),
    .X(_03904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08547_ (.A(_05487_),
    .X(_05489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _08548_ (.A1_N(\design_top.uart0.UART_RBAUD[14] ),
    .A2_N(_05482_),
    .B1(\design_top.uart0.UART_RBAUD[14] ),
    .B2(_05482_),
    .Y(_05490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08549_ (.A(_05489_),
    .B(_05490_),
    .Y(_03903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _08550_ (.A(\design_top.uart0.UART_RBAUD[13] ),
    .B(_05481_),
    .Y(_05491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _08551_ (.A1(_05482_),
    .A2(_05491_),
    .B1(_05489_),
    .Y(_03902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _08552_ (.A(\design_top.uart0.UART_RBAUD[12] ),
    .B(_05480_),
    .Y(_05492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _08553_ (.A1(_05481_),
    .A2(_05492_),
    .B1(_05489_),
    .Y(_03901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _08554_ (.A(\design_top.uart0.UART_RBAUD[11] ),
    .B(_05479_),
    .Y(_05493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _08555_ (.A1(_05480_),
    .A2(_05493_),
    .B1(_05489_),
    .Y(_03900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _08556_ (.A(\design_top.uart0.UART_RBAUD[10] ),
    .B(_05478_),
    .Y(_05494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _08557_ (.A1(_05479_),
    .A2(_05494_),
    .B1(_05487_),
    .Y(_03899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08558_ (.A(_05477_),
    .Y(_05495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _08559_ (.A1(\design_top.uart0.UART_RBAUD[8] ),
    .A2(_05476_),
    .B1(_05495_),
    .C1(_05487_),
    .X(_03898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08560_ (.A(_05474_),
    .Y(_05496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _08561_ (.A1(\design_top.uart0.UART_RBAUD[5] ),
    .A2(_05473_),
    .B1(_05496_),
    .C1(_05487_),
    .X(_03897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08562_ (.A(_05472_),
    .Y(_05497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _08563_ (.A1(\design_top.uart0.UART_RBAUD[2] ),
    .A2(_05471_),
    .B1(\design_top.uart0.UART_RBAUD[3] ),
    .X(_05498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _08564_ (.A1(_05497_),
    .A2(_05498_),
    .B1(_05488_),
    .X(_03896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08565_ (.A(\design_top.uart0.UART_RBAUD[0] ),
    .B(_05489_),
    .Y(_03895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08566_ (.A(\design_top.uart0.UART_XBAUD[1] ),
    .B(\design_top.uart0.UART_XBAUD[0] ),
    .C(\design_top.uart0.UART_XBAUD[2] ),
    .D(\design_top.uart0.UART_XBAUD[3] ),
    .X(_05499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08567_ (.A(\design_top.uart0.UART_XBAUD[4] ),
    .B(_05499_),
    .X(_05500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08568_ (.A(\design_top.uart0.UART_XBAUD[5] ),
    .B(_05500_),
    .X(_05501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08569_ (.A(\design_top.uart0.UART_XBAUD[6] ),
    .B(_05501_),
    .X(_05502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08570_ (.A(\design_top.uart0.UART_XBAUD[7] ),
    .B(_05502_),
    .X(_05503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08571_ (.A(\design_top.uart0.UART_XBAUD[8] ),
    .B(_05503_),
    .X(_05504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08572_ (.A(\design_top.uart0.UART_XBAUD[9] ),
    .B(_05504_),
    .X(_05505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08573_ (.A(\design_top.uart0.UART_XBAUD[10] ),
    .B(_05505_),
    .X(_05506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08574_ (.A(\design_top.uart0.UART_XBAUD[11] ),
    .B(_05506_),
    .X(_05507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08575_ (.A(\design_top.uart0.UART_XBAUD[12] ),
    .B(_05507_),
    .X(_05508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08576_ (.A(\design_top.uart0.UART_XBAUD[13] ),
    .B(_05508_),
    .X(_05509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08577_ (.A(\design_top.uart0.UART_XSTATE[1] ),
    .Y(_05510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08578_ (.A(\design_top.uart0.UART_XSTATE[2] ),
    .Y(_05511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _08579_ (.A(_05510_),
    .B(\design_top.uart0.UART_XSTATE[3] ),
    .C(_05511_),
    .X(_05512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _08580_ (.A(\design_top.uart0.UART_XBAUD[14] ),
    .B(_05509_),
    .C(\design_top.uart0.UART_XBAUD[15] ),
    .X(_05513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08581_ (.A(_05513_),
    .X(_02510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08582_ (.A1(\design_top.uart0.UART_XSTATE[0] ),
    .A2(_05512_),
    .B1(_02510_),
    .Y(_05514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08583_ (.A(_05514_),
    .Y(_05515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _08584_ (.A1(\design_top.uart0.UART_XBAUD[14] ),
    .A2(_05509_),
    .B1(\design_top.uart0.UART_XBAUD[15] ),
    .C1(_05515_),
    .X(_03894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08585_ (.A(_05514_),
    .X(_05516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08586_ (.A(_05516_),
    .X(_05517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _08587_ (.A1_N(\design_top.uart0.UART_XBAUD[14] ),
    .A2_N(_05509_),
    .B1(\design_top.uart0.UART_XBAUD[14] ),
    .B2(_05509_),
    .Y(_05518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08588_ (.A(_05517_),
    .B(_05518_),
    .Y(_03893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _08589_ (.A(\design_top.uart0.UART_XBAUD[13] ),
    .B(_05508_),
    .Y(_05519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _08590_ (.A1(_05509_),
    .A2(_05519_),
    .B1(_05517_),
    .Y(_03892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _08591_ (.A(\design_top.uart0.UART_XBAUD[12] ),
    .B(_05507_),
    .Y(_05520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _08592_ (.A1(_05508_),
    .A2(_05520_),
    .B1(_05517_),
    .Y(_03891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _08593_ (.A(\design_top.uart0.UART_XBAUD[11] ),
    .B(_05506_),
    .Y(_05521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08594_ (.A(_05516_),
    .X(_05522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _08595_ (.A1(_05507_),
    .A2(_05521_),
    .B1(_05522_),
    .Y(_03890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _08596_ (.A(\design_top.uart0.UART_XBAUD[10] ),
    .B(_05505_),
    .Y(_05523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _08597_ (.A1(_05506_),
    .A2(_05523_),
    .B1(_05522_),
    .Y(_03889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08598_ (.A(_05505_),
    .Y(_05524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _08599_ (.A1(\design_top.uart0.UART_XBAUD[9] ),
    .A2(_05504_),
    .B1(_05524_),
    .C1(_05522_),
    .X(_03888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08600_ (.A(_05504_),
    .Y(_05525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _08601_ (.A1(\design_top.uart0.UART_XBAUD[8] ),
    .A2(_05503_),
    .B1(_05525_),
    .C1(_05516_),
    .X(_03887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _08602_ (.A(\design_top.uart0.UART_XBAUD[7] ),
    .B(_05502_),
    .Y(_05526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _08603_ (.A1(_05503_),
    .A2(_05526_),
    .B1(_05522_),
    .Y(_03886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08604_ (.A(_05502_),
    .Y(_05527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _08605_ (.A1(\design_top.uart0.UART_XBAUD[6] ),
    .A2(_05501_),
    .B1(_05527_),
    .C1(_05516_),
    .X(_03885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08606_ (.A(_05501_),
    .Y(_05528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _08607_ (.A1(\design_top.uart0.UART_XBAUD[5] ),
    .A2(_05500_),
    .B1(_05528_),
    .C1(_05516_),
    .X(_03884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _08608_ (.A(\design_top.uart0.UART_XBAUD[4] ),
    .B(_05499_),
    .Y(_05529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _08609_ (.A1(_05500_),
    .A2(_05529_),
    .B1(_05522_),
    .Y(_03883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08610_ (.A(_05499_),
    .Y(_05530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08611_ (.A(\design_top.uart0.UART_XBAUD[1] ),
    .X(_05531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08612_ (.A(\design_top.uart0.UART_XBAUD[0] ),
    .X(_05532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _08613_ (.A1(_05531_),
    .A2(_05532_),
    .A3(\design_top.uart0.UART_XBAUD[2] ),
    .B1(\design_top.uart0.UART_XBAUD[3] ),
    .X(_05533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _08614_ (.A1(_05530_),
    .A2(_05533_),
    .B1(_05515_),
    .X(_03882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08615_ (.A1(_05531_),
    .A2(\design_top.uart0.UART_XBAUD[0] ),
    .B1(\design_top.uart0.UART_XBAUD[2] ),
    .Y(_05534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o311a_2 _08616_ (.A1(_05531_),
    .A2(_05532_),
    .A3(\design_top.uart0.UART_XBAUD[2] ),
    .B1(_05534_),
    .C1(_05515_),
    .X(_05535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08617_ (.A(_05535_),
    .Y(_03881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _08618_ (.A1_N(_05531_),
    .A2_N(_05532_),
    .B1(_05531_),
    .B2(_05532_),
    .Y(_05536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08619_ (.A(_05517_),
    .B(_05536_),
    .Y(_03880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08620_ (.A(_05532_),
    .B(_05517_),
    .Y(_03879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _08621_ (.A(_04717_),
    .B(_00003_),
    .X(_03878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _08622_ (.A(_04717_),
    .B(_00002_),
    .X(_03877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _08623_ (.A(_04717_),
    .B(_00001_),
    .X(_03876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _08624_ (.A(_04717_),
    .B(_00000_),
    .X(_03875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _08625_ (.A(_05295_),
    .B(\design_top.DACK[0] ),
    .C(\design_top.DACK[1] ),
    .X(_03874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _08626_ (.A(_05023_),
    .B(_00012_),
    .X(_03873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08627_ (.A(\design_top.uart0.UART_XSTATE[3] ),
    .Y(_05537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a41o_2 _08628_ (.A1(\design_top.uart0.UART_XSTATE[0] ),
    .A2(_05510_),
    .A3(_05537_),
    .A4(_05511_),
    .B1(_05296_),
    .X(_05538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08629_ (.A(\design_top.uart0.UART_XSTATE[0] ),
    .Y(_05539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _08630_ (.A(_05539_),
    .B(_02511_),
    .C(_05510_),
    .X(_05540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08631_ (.A(_05511_),
    .B(_05540_),
    .Y(_05541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _08632_ (.A1(_05539_),
    .A2(_02511_),
    .A3(_05512_),
    .B1(_05537_),
    .B2(_05541_),
    .X(_05542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08633_ (.A(_05538_),
    .B(_05542_),
    .Y(_03872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _08634_ (.A1(_05511_),
    .A2(_05540_),
    .B1(_05541_),
    .Y(_05543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08635_ (.A(_05538_),
    .B(_05543_),
    .X(_03871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08636_ (.A(_05540_),
    .Y(_05544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _08637_ (.A1(_05539_),
    .A2(_02511_),
    .B1(_05510_),
    .X(_05545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08638_ (.A(_05538_),
    .Y(_05546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08639_ (.A1(_05544_),
    .A2(_05545_),
    .B1(_05546_),
    .Y(_03870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08640_ (.A(_02511_),
    .Y(_05547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08641_ (.A1(_05539_),
    .A2(_02511_),
    .B1(\design_top.uart0.UART_XSTATE[0] ),
    .B2(_05547_),
    .C1(_05546_),
    .X(_03869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08642_ (.A(_05485_),
    .X(_05548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08643_ (.A(\design_top.uart0.UART_RSTATE[0] ),
    .Y(_05549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _08644_ (.A(_05549_),
    .B(_02513_),
    .C(_05484_),
    .X(_05550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08645_ (.A(\design_top.uart0.UART_RSTATE[3] ),
    .Y(_05551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08646_ (.A(_05551_),
    .X(_05552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08647_ (.A(\design_top.uart0.UART_RSTATE[1] ),
    .X(_05553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08648_ (.A(_05553_),
    .B(_05549_),
    .C(\design_top.uart0.UART_RSTATE[3] ),
    .D(\design_top.uart0.UART_RSTATE[2] ),
    .X(_05554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _08649_ (.A(_05022_),
    .B(_05554_),
    .Y(_05555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08650_ (.A(_05555_),
    .Y(_05556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08651_ (.A1(_05548_),
    .A2(_05550_),
    .B1(_05552_),
    .Y(_05557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o311a_2 _08652_ (.A1(_05548_),
    .A2(_05550_),
    .A3(_05552_),
    .B1(_05556_),
    .C1(_05557_),
    .X(_03868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08653_ (.A(\design_top.uart0.UART_RSTATE[2] ),
    .X(_05558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08654_ (.A(_05550_),
    .Y(_05559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08655_ (.A1(_05548_),
    .A2(_05550_),
    .B1(_05558_),
    .B2(_05559_),
    .X(_05560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08656_ (.A(_05555_),
    .B(_05560_),
    .X(_03867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08657_ (.A(_05549_),
    .X(_05561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08658_ (.A(_05484_),
    .X(_05562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _08659_ (.A1(_05561_),
    .A2(_02513_),
    .B1(_05562_),
    .X(_05563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08660_ (.A1(_05559_),
    .A2(_05563_),
    .B1(_05556_),
    .Y(_03866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08661_ (.A(\design_top.uart0.UART_RSTATE[0] ),
    .X(_05564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08662_ (.A(_02513_),
    .Y(_05565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08663_ (.A1(_05561_),
    .A2(_02513_),
    .B1(_05564_),
    .B2(_05565_),
    .C1(_05556_),
    .X(_03865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08664_ (.A(_05478_),
    .Y(_05566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _08665_ (.A(\design_top.uart0.UART_RBAUD[9] ),
    .B(_05477_),
    .X(_05567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08666_ (.A(_05486_),
    .X(_05568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _08667_ (.A1(_05566_),
    .A2(_05567_),
    .B1(_05568_),
    .X(_03864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _08668_ (.A1(\design_top.uart0.UART_RBAUD[7] ),
    .A2(_05475_),
    .B1_N(_05476_),
    .Y(_05569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08669_ (.A1(_05483_),
    .A2(_05569_),
    .B1(_05568_),
    .Y(_03863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08670_ (.A(_05475_),
    .Y(_05570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _08671_ (.A(\design_top.uart0.UART_RBAUD[6] ),
    .B(_05474_),
    .X(_05571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _08672_ (.A1(_05570_),
    .A2(_05571_),
    .B1(_05568_),
    .X(_03862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _08673_ (.A1(\design_top.uart0.UART_RBAUD[4] ),
    .A2(_05472_),
    .B1_N(_05473_),
    .Y(_05572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08674_ (.A1(_05483_),
    .A2(_05572_),
    .B1(_05568_),
    .Y(_03861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _08675_ (.A1_N(\design_top.uart0.UART_RBAUD[2] ),
    .A2_N(_05471_),
    .B1(\design_top.uart0.UART_RBAUD[2] ),
    .B2(_05471_),
    .Y(_05573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08676_ (.A(_00344_),
    .B(_05573_),
    .Y(_03860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _08677_ (.A1(\design_top.uart0.UART_RBAUD[1] ),
    .A2(\design_top.uart0.UART_RBAUD[0] ),
    .B1_N(_05471_),
    .Y(_05574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08678_ (.A1(_05483_),
    .A2(_05574_),
    .B1(_05568_),
    .Y(_03859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08679_ (.A(\design_top.core0.RESMODE[2] ),
    .Y(_05575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08680_ (.A(\design_top.core0.RESMODE[0] ),
    .B(\design_top.core0.RESMODE[1] ),
    .Y(_00902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _08681_ (.A(_05575_),
    .B(_00902_),
    .Y(_05576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _08682_ (.A1(\design_top.core0.RESMODE[3] ),
    .A2(_05576_),
    .B1(_05297_),
    .X(_03858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08683_ (.A1(_05575_),
    .A2(_00902_),
    .B1(_05062_),
    .Y(_05577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _08684_ (.A1(_05575_),
    .A2(_00902_),
    .A3(\design_top.core0.RESMODE[3] ),
    .B1(_05577_),
    .X(_03857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08685_ (.A(_05297_),
    .B(_00078_),
    .X(_03856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08686_ (.A(\design_top.core0.RESMODE[0] ),
    .Y(_05578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08687_ (.A(\design_top.core0.RESMODE[2] ),
    .B(\design_top.core0.RESMODE[3] ),
    .X(_05579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08688_ (.A(_05579_),
    .X(_00903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _08689_ (.A(\design_top.core0.RESMODE[0] ),
    .B(\design_top.core0.RESMODE[1] ),
    .C(_00903_),
    .X(_00046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _08690_ (.A1(_05578_),
    .A2(_00046_),
    .B1(_05297_),
    .X(_03855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08691_ (.A(_05062_),
    .X(_05580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08692_ (.A(\design_top.IRES[0] ),
    .B(\design_top.IRES[1] ),
    .X(_05581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _08693_ (.A(\design_top.IRES[2] ),
    .B(_05581_),
    .C(\design_top.IRES[3] ),
    .X(_05582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08694_ (.A(\design_top.IRES[4] ),
    .B(_05582_),
    .X(_05583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08695_ (.A(\design_top.IRES[5] ),
    .B(_05583_),
    .X(_05584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08696_ (.A(\design_top.IRES[6] ),
    .B(_05584_),
    .Y(_05585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08697_ (.A(_04883_),
    .X(_05586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08698_ (.A1(_05580_),
    .A2(_05585_),
    .B1(_05586_),
    .Y(_03854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _08699_ (.A1(\design_top.IRES[6] ),
    .A2(_05584_),
    .B1(_05585_),
    .Y(_05587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08700_ (.A1(_05580_),
    .A2(_05587_),
    .B1(_05586_),
    .Y(_03853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _08701_ (.A1(\design_top.IRES[5] ),
    .A2(_05583_),
    .B1_N(_05584_),
    .Y(_05588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08702_ (.A1(_05580_),
    .A2(_05588_),
    .B1(_05586_),
    .Y(_03852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _08703_ (.A1(\design_top.IRES[4] ),
    .A2(_05582_),
    .B1_N(_05583_),
    .Y(_05589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08704_ (.A1(_05580_),
    .A2(_05589_),
    .B1(_05586_),
    .Y(_03851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _08705_ (.A1(\design_top.IRES[2] ),
    .A2(_05581_),
    .B1(\design_top.IRES[3] ),
    .X(_05590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2b_2 _08706_ (.A_N(_05590_),
    .B(_05582_),
    .X(_05591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08707_ (.A1(_05580_),
    .A2(_05591_),
    .B1(_05586_),
    .Y(_03850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _08708_ (.A1_N(\design_top.IRES[2] ),
    .A2_N(_05581_),
    .B1(\design_top.IRES[2] ),
    .B2(_05581_),
    .Y(_05592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08709_ (.A1(_05023_),
    .A2(_05592_),
    .B1(_04883_),
    .Y(_03849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _08710_ (.A1(\design_top.IRES[0] ),
    .A2(\design_top.IRES[1] ),
    .B1_N(_05581_),
    .Y(_05593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08711_ (.A1(_05023_),
    .A2(_05593_),
    .B1(_04883_),
    .Y(_03848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08712_ (.A1(_05023_),
    .A2(\design_top.IRES[0] ),
    .B1(_04883_),
    .Y(_03847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08713_ (.A(_01440_),
    .X(_05594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08714_ (.A(_01439_),
    .Y(_05595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08715_ (.A(_05595_),
    .X(_05596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08716_ (.A(_01442_),
    .Y(_05597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08717_ (.A(_05594_),
    .B(_05596_),
    .C(_05597_),
    .D(_01441_),
    .X(_05598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08718_ (.A(_05598_),
    .X(_05599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08719_ (.A(_05599_),
    .X(_05600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08720_ (.A(_05599_),
    .Y(_05601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08721_ (.A(_05601_),
    .X(_05602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08722_ (.A(_01440_),
    .B(_01439_),
    .C(_01442_),
    .D(_01441_),
    .X(_05603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08723_ (.A(_05603_),
    .Y(_05604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08724_ (.A(\design_top.core0.XRES ),
    .B(_05604_),
    .X(_05605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08725_ (.A(_05605_),
    .X(_05606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08726_ (.A(_05606_),
    .X(_05607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08727_ (.A(_01438_),
    .B(_05607_),
    .Y(_05608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08728_ (.A(_05608_),
    .X(_05609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08729_ (.A1(\design_top.core0.REG2[9][31] ),
    .A2(_05600_),
    .B1(_05602_),
    .B2(_05609_),
    .X(_03846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08730_ (.A(_05600_),
    .X(_05610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08731_ (.A(_02402_),
    .B(_05607_),
    .Y(_05611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08732_ (.A(_05611_),
    .X(_05612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08733_ (.A(_05602_),
    .X(_05613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08734_ (.A1(_05610_),
    .A2(_05612_),
    .B1(\design_top.core0.REG2[9][30] ),
    .B2(_05613_),
    .X(_03845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08735_ (.A(_02382_),
    .B(_05607_),
    .Y(_05614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08736_ (.A(_05614_),
    .X(_05615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08737_ (.A1(_05610_),
    .A2(_05615_),
    .B1(\design_top.core0.REG2[9][29] ),
    .B2(_05613_),
    .X(_03844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08738_ (.A(_02363_),
    .B(_05607_),
    .Y(_05616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08739_ (.A(_05616_),
    .X(_05617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08740_ (.A1(_05610_),
    .A2(_05617_),
    .B1(\design_top.core0.REG2[9][28] ),
    .B2(_05613_),
    .X(_03843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08741_ (.A(_02341_),
    .B(_05607_),
    .Y(_05618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08742_ (.A(_05618_),
    .X(_05619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08743_ (.A1(_05610_),
    .A2(_05619_),
    .B1(\design_top.core0.REG2[9][27] ),
    .B2(_05613_),
    .X(_03842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08744_ (.A(_05606_),
    .X(_05620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08745_ (.A(_02322_),
    .B(_05620_),
    .Y(_05621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08746_ (.A(_05621_),
    .X(_05622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08747_ (.A1(_05610_),
    .A2(_05622_),
    .B1(\design_top.core0.REG2[9][26] ),
    .B2(_05613_),
    .X(_03841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08748_ (.A(_05600_),
    .X(_05623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08749_ (.A(_02300_),
    .B(_05620_),
    .Y(_05624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08750_ (.A(_05624_),
    .X(_05625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08751_ (.A(_05602_),
    .X(_05626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08752_ (.A1(_05623_),
    .A2(_05625_),
    .B1(\design_top.core0.REG2[9][25] ),
    .B2(_05626_),
    .X(_03840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08753_ (.A(_02280_),
    .B(_05620_),
    .Y(_05627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08754_ (.A(_05627_),
    .X(_05628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08755_ (.A1(_05623_),
    .A2(_05628_),
    .B1(\design_top.core0.REG2[9][24] ),
    .B2(_05626_),
    .X(_03839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08756_ (.A(_02258_),
    .B(_05620_),
    .Y(_05629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08757_ (.A(_05629_),
    .X(_05630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08758_ (.A1(_05623_),
    .A2(_05630_),
    .B1(\design_top.core0.REG2[9][23] ),
    .B2(_05626_),
    .X(_03838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08759_ (.A(_02240_),
    .B(_05620_),
    .Y(_05631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08760_ (.A(_05631_),
    .X(_05632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08761_ (.A1(_05623_),
    .A2(_05632_),
    .B1(\design_top.core0.REG2[9][22] ),
    .B2(_05626_),
    .X(_03837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08762_ (.A(_05606_),
    .X(_05633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08763_ (.A(_02218_),
    .B(_05633_),
    .Y(_05634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08764_ (.A(_05634_),
    .X(_05635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08765_ (.A1(_05623_),
    .A2(_05635_),
    .B1(\design_top.core0.REG2[9][21] ),
    .B2(_05626_),
    .X(_03836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08766_ (.A(_05600_),
    .X(_05636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08767_ (.A(_02198_),
    .B(_05633_),
    .Y(_05637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08768_ (.A(_05637_),
    .X(_05638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08769_ (.A(_05602_),
    .X(_05639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08770_ (.A1(_05636_),
    .A2(_05638_),
    .B1(\design_top.core0.REG2[9][20] ),
    .B2(_05639_),
    .X(_03835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08771_ (.A(_02176_),
    .B(_05633_),
    .Y(_05640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08772_ (.A(_05640_),
    .X(_05641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08773_ (.A1(_05636_),
    .A2(_05641_),
    .B1(\design_top.core0.REG2[9][19] ),
    .B2(_05639_),
    .X(_03834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08774_ (.A(_02157_),
    .B(_05633_),
    .Y(_05642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08775_ (.A(_05642_),
    .X(_05643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08776_ (.A1(_05636_),
    .A2(_05643_),
    .B1(\design_top.core0.REG2[9][18] ),
    .B2(_05639_),
    .X(_03833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08777_ (.A(_02134_),
    .B(_05633_),
    .Y(_05644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08778_ (.A(_05644_),
    .X(_05645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08779_ (.A1(_05636_),
    .A2(_05645_),
    .B1(\design_top.core0.REG2[9][17] ),
    .B2(_05639_),
    .X(_03832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08780_ (.A(_05606_),
    .X(_05646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08781_ (.A(_02114_),
    .B(_05646_),
    .Y(_05647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08782_ (.A(_05647_),
    .X(_05648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08783_ (.A1(_05636_),
    .A2(_05648_),
    .B1(\design_top.core0.REG2[9][16] ),
    .B2(_05639_),
    .X(_03831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08784_ (.A(_05599_),
    .X(_05649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08785_ (.A(_02092_),
    .B(_05646_),
    .Y(_05650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08786_ (.A(_05650_),
    .X(_05651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08787_ (.A(_05601_),
    .X(_05652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08788_ (.A1(_05649_),
    .A2(_05651_),
    .B1(\design_top.core0.REG2[9][15] ),
    .B2(_05652_),
    .X(_03830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08789_ (.A(_02076_),
    .B(_05646_),
    .Y(_05653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08790_ (.A(_05653_),
    .X(_05654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08791_ (.A1(_05649_),
    .A2(_05654_),
    .B1(\design_top.core0.REG2[9][14] ),
    .B2(_05652_),
    .X(_03829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08792_ (.A(_00045_),
    .X(_05655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08793_ (.A(_05655_),
    .X(_05656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08794_ (.A1(\design_top.core0.REG2[9][13] ),
    .A2(_05600_),
    .B1(_05656_),
    .B2(_05602_),
    .X(_03828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08795_ (.A(_02027_),
    .B(_05646_),
    .Y(_05657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08796_ (.A(_05657_),
    .X(_05658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08797_ (.A1(_05649_),
    .A2(_05658_),
    .B1(\design_top.core0.REG2[9][12] ),
    .B2(_05652_),
    .X(_03827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08798_ (.A(_02003_),
    .B(_05646_),
    .Y(_05659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08799_ (.A(_05659_),
    .X(_05660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08800_ (.A1(_05649_),
    .A2(_05660_),
    .B1(\design_top.core0.REG2[9][11] ),
    .B2(_05652_),
    .X(_03826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08801_ (.A(_05605_),
    .X(_05661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08802_ (.A(_01982_),
    .B(_05661_),
    .Y(_05662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08803_ (.A(_05662_),
    .X(_05663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08804_ (.A1(_05649_),
    .A2(_05663_),
    .B1(\design_top.core0.REG2[9][10] ),
    .B2(_05652_),
    .X(_03825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08805_ (.A(_05599_),
    .X(_05664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08806_ (.A(_01958_),
    .B(_05661_),
    .Y(_05665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08807_ (.A(_05665_),
    .X(_05666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08808_ (.A(_05601_),
    .X(_05667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08809_ (.A1(_05664_),
    .A2(_05666_),
    .B1(\design_top.core0.REG2[9][9] ),
    .B2(_05667_),
    .X(_03824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08810_ (.A(_01936_),
    .B(_05661_),
    .Y(_05668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08811_ (.A(_05668_),
    .X(_05669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08812_ (.A1(_05664_),
    .A2(_05669_),
    .B1(\design_top.core0.REG2[9][8] ),
    .B2(_05667_),
    .X(_03823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08813_ (.A(_01912_),
    .B(_05661_),
    .Y(_05670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08814_ (.A(_05670_),
    .X(_05671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08815_ (.A1(_05664_),
    .A2(_05671_),
    .B1(\design_top.core0.REG2[9][7] ),
    .B2(_05667_),
    .X(_03822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08816_ (.A(_01889_),
    .B(_05661_),
    .Y(_05672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08817_ (.A(_05672_),
    .X(_05673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08818_ (.A1(_05664_),
    .A2(_05673_),
    .B1(\design_top.core0.REG2[9][6] ),
    .B2(_05667_),
    .X(_03821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08819_ (.A(_05605_),
    .X(_05674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08820_ (.A(_01843_),
    .B(_05674_),
    .Y(_05675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08821_ (.A(_05675_),
    .X(_05676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08822_ (.A1(_05664_),
    .A2(_05676_),
    .B1(\design_top.core0.REG2[9][5] ),
    .B2(_05667_),
    .X(_03820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08823_ (.A(_05599_),
    .X(_05677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08824_ (.A(_01800_),
    .B(_05674_),
    .Y(_05678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08825_ (.A(_05678_),
    .X(_05679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08826_ (.A(_05601_),
    .X(_05680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08827_ (.A1(_05677_),
    .A2(_05679_),
    .B1(\design_top.core0.REG2[9][4] ),
    .B2(_05680_),
    .X(_03819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08828_ (.A(_01756_),
    .B(_05674_),
    .Y(_05681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08829_ (.A(_05681_),
    .X(_05682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08830_ (.A1(_05677_),
    .A2(_05682_),
    .B1(\design_top.core0.REG2[9][3] ),
    .B2(_05680_),
    .X(_03818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08831_ (.A(_01708_),
    .B(_05674_),
    .Y(_05683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08832_ (.A(_05683_),
    .X(_05684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08833_ (.A1(_05677_),
    .A2(_05684_),
    .B1(\design_top.core0.REG2[9][2] ),
    .B2(_05680_),
    .X(_03817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08834_ (.A(_01653_),
    .B(_05674_),
    .Y(_05685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08835_ (.A(_05685_),
    .X(_05686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08836_ (.A1(_05677_),
    .A2(_05686_),
    .B1(\design_top.core0.REG2[9][1] ),
    .B2(_05680_),
    .X(_03816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08837_ (.A(_01585_),
    .B(_05606_),
    .Y(_05687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08838_ (.A(_05687_),
    .X(_05688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08839_ (.A1(_05677_),
    .A2(_05688_),
    .B1(\design_top.core0.REG2[9][0] ),
    .B2(_05680_),
    .X(_03815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08840_ (.A(_00549_),
    .B(_04869_),
    .X(_05689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08841_ (.A(_05689_),
    .X(_05690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08842_ (.A(_04907_),
    .B(_05690_),
    .Y(_00587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08843_ (.A(_04915_),
    .B(_00587_),
    .X(_05691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08844_ (.A(_05691_),
    .X(_05692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08845_ (.A(_05691_),
    .Y(_05693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08846_ (.A(_05693_),
    .X(_05694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08847_ (.A1(_00220_),
    .A2(_05692_),
    .B1(\design_top.MEM[14][7] ),
    .B2(_05694_),
    .X(_03814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08848_ (.A1(_00219_),
    .A2(_05692_),
    .B1(\design_top.MEM[14][6] ),
    .B2(_05694_),
    .X(_03813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08849_ (.A1(_00218_),
    .A2(_05692_),
    .B1(\design_top.MEM[14][5] ),
    .B2(_05694_),
    .X(_03812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08850_ (.A1(_00217_),
    .A2(_05692_),
    .B1(\design_top.MEM[14][4] ),
    .B2(_05694_),
    .X(_03811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08851_ (.A1(_00216_),
    .A2(_05692_),
    .B1(\design_top.MEM[14][3] ),
    .B2(_05694_),
    .X(_03810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08852_ (.A1(_00215_),
    .A2(_05691_),
    .B1(\design_top.MEM[14][2] ),
    .B2(_05693_),
    .X(_03809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08853_ (.A1(_00214_),
    .A2(_05691_),
    .B1(\design_top.MEM[14][1] ),
    .B2(_05693_),
    .X(_03808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08854_ (.A1(_00213_),
    .A2(_05691_),
    .B1(\design_top.MEM[14][0] ),
    .B2(_05693_),
    .X(_03807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _08855_ (.A(_01111_),
    .B(\design_top.DACK[1] ),
    .C(_00547_),
    .Y(_05695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08856_ (.A(_05017_),
    .B(_04873_),
    .X(_05696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08857_ (.A(_05696_),
    .Y(_05697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _08858_ (.A1(io_out[12]),
    .A2(_05695_),
    .A3(_05697_),
    .B1(_05296_),
    .X(_05698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _08859_ (.A0(\design_top.uart0.UART_RACK ),
    .A1(\design_top.uart0.UART_RREQ ),
    .S(_05698_),
    .X(_03806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08860_ (.A(\design_top.uart0.UART_XACK ),
    .Y(_05699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08861_ (.A(_04620_),
    .B(_04720_),
    .C(_00547_),
    .D(_05696_),
    .X(_05700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08862_ (.A(_05700_),
    .X(_05701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _08863_ (.A0(_05699_),
    .A1(\design_top.uart0.UART_XREQ ),
    .S(_05701_),
    .X(_03805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _08864_ (.A0(\design_top.DATAO[15] ),
    .A1(\design_top.uart0.UART_XFIFO[7] ),
    .S(_05701_),
    .X(_03804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _08865_ (.A0(\design_top.DATAO[14] ),
    .A1(\design_top.uart0.UART_XFIFO[6] ),
    .S(_05701_),
    .X(_03803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _08866_ (.A0(\design_top.DATAO[13] ),
    .A1(\design_top.uart0.UART_XFIFO[5] ),
    .S(_05701_),
    .X(_03802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _08867_ (.A0(\design_top.DATAO[12] ),
    .A1(\design_top.uart0.UART_XFIFO[4] ),
    .S(_05701_),
    .X(_03801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _08868_ (.A0(\design_top.DATAO[11] ),
    .A1(\design_top.uart0.UART_XFIFO[3] ),
    .S(_05700_),
    .X(_03800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _08869_ (.A0(\design_top.DATAO[10] ),
    .A1(\design_top.uart0.UART_XFIFO[2] ),
    .S(_05700_),
    .X(_03799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _08870_ (.A0(\design_top.DATAO[9] ),
    .A1(\design_top.uart0.UART_XFIFO[1] ),
    .S(_05700_),
    .X(_03798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _08871_ (.A0(\design_top.DATAO[8] ),
    .A1(\design_top.uart0.UART_XFIFO[0] ),
    .S(_05700_),
    .X(_03797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08872_ (.A(_04960_),
    .B(_05690_),
    .Y(_00585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08873_ (.A(_04965_),
    .B(_00585_),
    .X(_05702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08874_ (.A(_05702_),
    .X(_05703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08875_ (.A(_05702_),
    .Y(_05704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08876_ (.A(_05704_),
    .X(_05705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08877_ (.A1(_00180_),
    .A2(_05703_),
    .B1(\design_top.MEM[0][7] ),
    .B2(_05705_),
    .X(_03796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08878_ (.A1(_00179_),
    .A2(_05703_),
    .B1(\design_top.MEM[0][6] ),
    .B2(_05705_),
    .X(_03795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08879_ (.A1(_00178_),
    .A2(_05703_),
    .B1(\design_top.MEM[0][5] ),
    .B2(_05705_),
    .X(_03794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08880_ (.A1(_00177_),
    .A2(_05703_),
    .B1(\design_top.MEM[0][4] ),
    .B2(_05705_),
    .X(_03793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08881_ (.A1(_00176_),
    .A2(_05703_),
    .B1(\design_top.MEM[0][3] ),
    .B2(_05705_),
    .X(_03792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08882_ (.A1(_00175_),
    .A2(_05702_),
    .B1(\design_top.MEM[0][2] ),
    .B2(_05704_),
    .X(_03791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08883_ (.A1(_00174_),
    .A2(_05702_),
    .B1(\design_top.MEM[0][1] ),
    .B2(_05704_),
    .X(_03790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08884_ (.A1(_00173_),
    .A2(_05702_),
    .B1(\design_top.MEM[0][0] ),
    .B2(_05704_),
    .X(_03789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08885_ (.A(_04976_),
    .B(_05690_),
    .Y(_00584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08886_ (.A(_04979_),
    .B(_00584_),
    .X(_05706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08887_ (.A(_05706_),
    .X(_05707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08888_ (.A(_05706_),
    .Y(_05708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08889_ (.A(_05708_),
    .X(_05709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08890_ (.A1(_00188_),
    .A2(_05707_),
    .B1(\design_top.MEM[10][7] ),
    .B2(_05709_),
    .X(_03788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08891_ (.A1(_00187_),
    .A2(_05707_),
    .B1(\design_top.MEM[10][6] ),
    .B2(_05709_),
    .X(_03787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08892_ (.A1(_00186_),
    .A2(_05707_),
    .B1(\design_top.MEM[10][5] ),
    .B2(_05709_),
    .X(_03786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08893_ (.A1(_00185_),
    .A2(_05707_),
    .B1(\design_top.MEM[10][4] ),
    .B2(_05709_),
    .X(_03785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08894_ (.A1(_00184_),
    .A2(_05707_),
    .B1(\design_top.MEM[10][3] ),
    .B2(_05709_),
    .X(_03784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08895_ (.A1(_00183_),
    .A2(_05706_),
    .B1(\design_top.MEM[10][2] ),
    .B2(_05708_),
    .X(_03783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08896_ (.A1(_00182_),
    .A2(_05706_),
    .B1(\design_top.MEM[10][1] ),
    .B2(_05708_),
    .X(_03782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08897_ (.A1(_00181_),
    .A2(_05706_),
    .B1(\design_top.MEM[10][0] ),
    .B2(_05708_),
    .X(_03781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08898_ (.A(_04991_),
    .B(_05690_),
    .Y(_00565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08899_ (.A(_04995_),
    .B(_00565_),
    .X(_05710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08900_ (.A(_05710_),
    .X(_05711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08901_ (.A(_05710_),
    .Y(_05712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08902_ (.A(_05712_),
    .X(_05713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08903_ (.A1(_00196_),
    .A2(_05711_),
    .B1(\design_top.MEM[11][7] ),
    .B2(_05713_),
    .X(_03780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08904_ (.A1(_00195_),
    .A2(_05711_),
    .B1(\design_top.MEM[11][6] ),
    .B2(_05713_),
    .X(_03779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08905_ (.A1(_00194_),
    .A2(_05711_),
    .B1(\design_top.MEM[11][5] ),
    .B2(_05713_),
    .X(_03778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08906_ (.A1(_00193_),
    .A2(_05711_),
    .B1(\design_top.MEM[11][4] ),
    .B2(_05713_),
    .X(_03777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08907_ (.A1(_00192_),
    .A2(_05711_),
    .B1(\design_top.MEM[11][3] ),
    .B2(_05713_),
    .X(_03776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08908_ (.A1(_00191_),
    .A2(_05710_),
    .B1(\design_top.MEM[11][2] ),
    .B2(_05712_),
    .X(_03775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08909_ (.A1(_00190_),
    .A2(_05710_),
    .B1(\design_top.MEM[11][1] ),
    .B2(_05712_),
    .X(_03774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08910_ (.A1(_00189_),
    .A2(_05710_),
    .B1(\design_top.MEM[11][0] ),
    .B2(_05712_),
    .X(_03773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08911_ (.A(_05007_),
    .B(_05690_),
    .Y(_00564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08912_ (.A(_05010_),
    .B(_00564_),
    .X(_05714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08913_ (.A(_05714_),
    .X(_05715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08914_ (.A(_05714_),
    .Y(_05716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08915_ (.A(_05716_),
    .X(_05717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08916_ (.A1(_00204_),
    .A2(_05715_),
    .B1(\design_top.MEM[12][7] ),
    .B2(_05717_),
    .X(_03772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08917_ (.A1(_00203_),
    .A2(_05715_),
    .B1(\design_top.MEM[12][6] ),
    .B2(_05717_),
    .X(_03771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08918_ (.A1(_00202_),
    .A2(_05715_),
    .B1(\design_top.MEM[12][5] ),
    .B2(_05717_),
    .X(_03770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08919_ (.A1(_00201_),
    .A2(_05715_),
    .B1(\design_top.MEM[12][4] ),
    .B2(_05717_),
    .X(_03769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08920_ (.A1(_00200_),
    .A2(_05715_),
    .B1(\design_top.MEM[12][3] ),
    .B2(_05717_),
    .X(_03768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08921_ (.A1(_00199_),
    .A2(_05714_),
    .B1(\design_top.MEM[12][2] ),
    .B2(_05716_),
    .X(_03767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08922_ (.A1(_00198_),
    .A2(_05714_),
    .B1(\design_top.MEM[12][1] ),
    .B2(_05716_),
    .X(_03766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08923_ (.A1(_00197_),
    .A2(_05714_),
    .B1(\design_top.MEM[12][0] ),
    .B2(_05716_),
    .X(_03765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08924_ (.A(\design_top.IRES[7] ),
    .B(_05034_),
    .X(_05718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08925_ (.A(_05718_),
    .X(_05719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08926_ (.A(_05719_),
    .X(_05720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08927_ (.A(_05720_),
    .X(_05721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08928_ (.A(_05718_),
    .Y(_05722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08929_ (.A(_05722_),
    .X(_05723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08930_ (.A1(\design_top.TIMER[31] ),
    .A2(_05721_),
    .B1(_00037_),
    .B2(_05723_),
    .X(_03764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08931_ (.A1(\design_top.TIMER[30] ),
    .A2(_05721_),
    .B1(_00036_),
    .B2(_05723_),
    .X(_03763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08932_ (.A1(\design_top.TIMER[29] ),
    .A2(_05721_),
    .B1(_00034_),
    .B2(_05723_),
    .X(_03762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08933_ (.A1(\design_top.TIMER[28] ),
    .A2(_05721_),
    .B1(_00033_),
    .B2(_05723_),
    .X(_03761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08934_ (.A(_05722_),
    .X(_05724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08935_ (.A(_05724_),
    .X(_05725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08936_ (.A1(\design_top.TIMER[27] ),
    .A2(_05721_),
    .B1(_00032_),
    .B2(_05725_),
    .X(_03760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08937_ (.A(_05720_),
    .X(_05726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08938_ (.A1(\design_top.TIMER[26] ),
    .A2(_05726_),
    .B1(_00031_),
    .B2(_05725_),
    .X(_03759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08939_ (.A1(\design_top.TIMER[25] ),
    .A2(_05726_),
    .B1(_00030_),
    .B2(_05725_),
    .X(_03758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08940_ (.A1(\design_top.TIMER[24] ),
    .A2(_05726_),
    .B1(_00029_),
    .B2(_05725_),
    .X(_03757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08941_ (.A1(\design_top.TIMER[23] ),
    .A2(_05726_),
    .B1(_00028_),
    .B2(_05725_),
    .X(_03756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08942_ (.A(_05724_),
    .X(_05727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08943_ (.A1(\design_top.TIMER[22] ),
    .A2(_05726_),
    .B1(_00027_),
    .B2(_05727_),
    .X(_03755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08944_ (.A(_05719_),
    .X(_05728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08945_ (.A1(\design_top.TIMER[21] ),
    .A2(_05728_),
    .B1(_00026_),
    .B2(_05727_),
    .X(_03754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08946_ (.A1(\design_top.TIMER[20] ),
    .A2(_05728_),
    .B1(_00025_),
    .B2(_05727_),
    .X(_03753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08947_ (.A1(\design_top.TIMER[19] ),
    .A2(_05728_),
    .B1(_00023_),
    .B2(_05727_),
    .X(_03752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08948_ (.A1(\design_top.TIMER[18] ),
    .A2(_05728_),
    .B1(_00022_),
    .B2(_05727_),
    .X(_03751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08949_ (.A(_05722_),
    .X(_05729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08950_ (.A1(\design_top.TIMER[17] ),
    .A2(_05728_),
    .B1(_00021_),
    .B2(_05729_),
    .X(_03750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08951_ (.A(_05719_),
    .X(_05730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08952_ (.A1(\design_top.TIMER[16] ),
    .A2(_05730_),
    .B1(_00020_),
    .B2(_05729_),
    .X(_03749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08953_ (.A1(\design_top.TIMER[15] ),
    .A2(_05730_),
    .B1(_00019_),
    .B2(_05729_),
    .X(_03748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08954_ (.A1(\design_top.TIMER[14] ),
    .A2(_05730_),
    .B1(_00018_),
    .B2(_05729_),
    .X(_03747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08955_ (.A1(\design_top.TIMER[13] ),
    .A2(_05730_),
    .B1(_00017_),
    .B2(_05729_),
    .X(_03746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08956_ (.A(_05722_),
    .X(_05731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08957_ (.A1(\design_top.TIMER[12] ),
    .A2(_05730_),
    .B1(_00016_),
    .B2(_05731_),
    .X(_03745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08958_ (.A(_05719_),
    .X(_05732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08959_ (.A1(\design_top.TIMER[11] ),
    .A2(_05732_),
    .B1(_00015_),
    .B2(_05731_),
    .X(_03744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08960_ (.A1(\design_top.TIMER[10] ),
    .A2(_05732_),
    .B1(_00014_),
    .B2(_05731_),
    .X(_03743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08961_ (.A1(\design_top.TIMER[9] ),
    .A2(_05732_),
    .B1(_00044_),
    .B2(_05731_),
    .X(_03742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08962_ (.A1(\design_top.TIMER[8] ),
    .A2(_05732_),
    .B1(_00043_),
    .B2(_05731_),
    .X(_03741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08963_ (.A(_05722_),
    .X(_05733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08964_ (.A1(\design_top.TIMER[7] ),
    .A2(_05732_),
    .B1(_00042_),
    .B2(_05733_),
    .X(_03740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08965_ (.A(_05719_),
    .X(_05734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08966_ (.A1(\design_top.TIMER[6] ),
    .A2(_05734_),
    .B1(_00041_),
    .B2(_05733_),
    .X(_03739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08967_ (.A1(\design_top.TIMER[5] ),
    .A2(_05734_),
    .B1(_00040_),
    .B2(_05733_),
    .X(_03738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08968_ (.A1(\design_top.TIMER[4] ),
    .A2(_05734_),
    .B1(_00039_),
    .B2(_05733_),
    .X(_03737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08969_ (.A1(\design_top.TIMER[3] ),
    .A2(_05734_),
    .B1(_00038_),
    .B2(_05733_),
    .X(_03736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08970_ (.A1(\design_top.TIMER[2] ),
    .A2(_05734_),
    .B1(_00035_),
    .B2(_05724_),
    .X(_03735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08971_ (.A1(\design_top.TIMER[1] ),
    .A2(_05720_),
    .B1(_00024_),
    .B2(_05724_),
    .X(_03734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08972_ (.A1(\design_top.TIMER[0] ),
    .A2(_05720_),
    .B1(_00013_),
    .B2(_05724_),
    .X(_03733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08973_ (.A(_05058_),
    .Y(_00345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08974_ (.A(io_out[14]),
    .Y(_05735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _08975_ (.A1(_05058_),
    .A2(_05720_),
    .B1(io_out[14]),
    .X(_05736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _08976_ (.A1(_00345_),
    .A2(_05723_),
    .A3(_05735_),
    .B1(_05736_),
    .X(_03732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08977_ (.A(_05689_),
    .X(_05737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08978_ (.A(_05083_),
    .B(_05737_),
    .Y(_00563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08979_ (.A(_05086_),
    .B(_00563_),
    .X(_05738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08980_ (.A(_05738_),
    .X(_05739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08981_ (.A(_05738_),
    .Y(_05740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08982_ (.A(_05740_),
    .X(_05741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08983_ (.A1(_00212_),
    .A2(_05739_),
    .B1(\design_top.MEM[13][7] ),
    .B2(_05741_),
    .X(_03731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08984_ (.A1(_00211_),
    .A2(_05739_),
    .B1(\design_top.MEM[13][6] ),
    .B2(_05741_),
    .X(_03730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08985_ (.A1(_00210_),
    .A2(_05739_),
    .B1(\design_top.MEM[13][5] ),
    .B2(_05741_),
    .X(_03729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08986_ (.A1(_00209_),
    .A2(_05739_),
    .B1(\design_top.MEM[13][4] ),
    .B2(_05741_),
    .X(_03728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08987_ (.A1(_00208_),
    .A2(_05739_),
    .B1(\design_top.MEM[13][3] ),
    .B2(_05741_),
    .X(_03727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08988_ (.A1(_00207_),
    .A2(_05738_),
    .B1(\design_top.MEM[13][2] ),
    .B2(_05740_),
    .X(_03726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08989_ (.A1(_00206_),
    .A2(_05738_),
    .B1(\design_top.MEM[13][1] ),
    .B2(_05740_),
    .X(_03725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08990_ (.A1(_00205_),
    .A2(_05738_),
    .B1(\design_top.MEM[13][0] ),
    .B2(_05740_),
    .X(_03724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08991_ (.A(\design_top.core0.XJALR ),
    .B(\design_top.core0.XJAL ),
    .C(\design_top.core0.XRCC ),
    .D(\design_top.core0.XMCC ),
    .X(_05742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08992_ (.A(\design_top.core0.XLCC ),
    .B(\design_top.core0.XAUIPC ),
    .C(\design_top.core0.XLUI ),
    .D(_05742_),
    .X(_05743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _08993_ (.A1(_00309_),
    .A2(_05743_),
    .B1(_05604_),
    .Y(_05744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _08994_ (.A1(_04619_),
    .A2(_05744_),
    .B1(_04715_),
    .X(_05745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08995_ (.A(_05745_),
    .X(_05746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08996_ (.A(_05598_),
    .B(_05746_),
    .X(_05747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08997_ (.A(_05747_),
    .X(_05748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08998_ (.A(_05608_),
    .X(_05749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08999_ (.A(_05749_),
    .X(_05750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09000_ (.A(_05747_),
    .Y(_05751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09001_ (.A(_05751_),
    .X(_05752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09002_ (.A1(\design_top.core0.REG1[9][31] ),
    .A2(_05748_),
    .B1(_05750_),
    .B2(_05752_),
    .X(_03723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09003_ (.A(_05611_),
    .X(_05753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09004_ (.A(_05753_),
    .X(_05754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09005_ (.A(_05748_),
    .X(_05755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09006_ (.A(_05752_),
    .X(_05756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09007_ (.A1(_05754_),
    .A2(_05755_),
    .B1(\design_top.core0.REG1[9][30] ),
    .B2(_05756_),
    .X(_03722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09008_ (.A(_05614_),
    .X(_05757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09009_ (.A(_05757_),
    .X(_05758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09010_ (.A1(_05758_),
    .A2(_05755_),
    .B1(\design_top.core0.REG1[9][29] ),
    .B2(_05756_),
    .X(_03721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09011_ (.A(_05616_),
    .X(_05759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09012_ (.A(_05759_),
    .X(_05760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09013_ (.A1(_05760_),
    .A2(_05755_),
    .B1(\design_top.core0.REG1[9][28] ),
    .B2(_05756_),
    .X(_03720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09014_ (.A(_05618_),
    .X(_05761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09015_ (.A(_05761_),
    .X(_05762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09016_ (.A1(_05762_),
    .A2(_05755_),
    .B1(\design_top.core0.REG1[9][27] ),
    .B2(_05756_),
    .X(_03719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09017_ (.A(_05621_),
    .X(_05763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09018_ (.A(_05763_),
    .X(_05764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09019_ (.A1(_05764_),
    .A2(_05755_),
    .B1(\design_top.core0.REG1[9][26] ),
    .B2(_05756_),
    .X(_03718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09020_ (.A(_05624_),
    .X(_05765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09021_ (.A(_05765_),
    .X(_05766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09022_ (.A(_05748_),
    .X(_05767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09023_ (.A(_05752_),
    .X(_05768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09024_ (.A1(_05766_),
    .A2(_05767_),
    .B1(\design_top.core0.REG1[9][25] ),
    .B2(_05768_),
    .X(_03717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09025_ (.A(_05627_),
    .X(_05769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09026_ (.A(_05769_),
    .X(_05770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09027_ (.A1(_05770_),
    .A2(_05767_),
    .B1(\design_top.core0.REG1[9][24] ),
    .B2(_05768_),
    .X(_03716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09028_ (.A(_05629_),
    .X(_05771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09029_ (.A(_05771_),
    .X(_05772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09030_ (.A1(_05772_),
    .A2(_05767_),
    .B1(\design_top.core0.REG1[9][23] ),
    .B2(_05768_),
    .X(_03715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09031_ (.A(_05631_),
    .X(_05773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09032_ (.A(_05773_),
    .X(_05774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09033_ (.A1(_05774_),
    .A2(_05767_),
    .B1(\design_top.core0.REG1[9][22] ),
    .B2(_05768_),
    .X(_03714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09034_ (.A(_05634_),
    .X(_05775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09035_ (.A(_05775_),
    .X(_05776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09036_ (.A1(_05776_),
    .A2(_05767_),
    .B1(\design_top.core0.REG1[9][21] ),
    .B2(_05768_),
    .X(_03713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09037_ (.A(_05637_),
    .X(_05777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09038_ (.A(_05777_),
    .X(_05778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09039_ (.A(_05748_),
    .X(_05779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09040_ (.A(_05752_),
    .X(_05780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09041_ (.A1(_05778_),
    .A2(_05779_),
    .B1(\design_top.core0.REG1[9][20] ),
    .B2(_05780_),
    .X(_03712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09042_ (.A(_05640_),
    .X(_05781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09043_ (.A(_05781_),
    .X(_05782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09044_ (.A1(_05782_),
    .A2(_05779_),
    .B1(\design_top.core0.REG1[9][19] ),
    .B2(_05780_),
    .X(_03711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09045_ (.A(_05642_),
    .X(_05783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09046_ (.A(_05783_),
    .X(_05784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09047_ (.A1(_05784_),
    .A2(_05779_),
    .B1(\design_top.core0.REG1[9][18] ),
    .B2(_05780_),
    .X(_03710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09048_ (.A(_05644_),
    .X(_05785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09049_ (.A(_05785_),
    .X(_05786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09050_ (.A1(_05786_),
    .A2(_05779_),
    .B1(\design_top.core0.REG1[9][17] ),
    .B2(_05780_),
    .X(_03709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09051_ (.A(_05647_),
    .X(_05787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09052_ (.A(_05787_),
    .X(_05788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09053_ (.A1(_05788_),
    .A2(_05779_),
    .B1(\design_top.core0.REG1[9][16] ),
    .B2(_05780_),
    .X(_03708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09054_ (.A(_05650_),
    .X(_05789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09055_ (.A(_05789_),
    .X(_05790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09056_ (.A(_05747_),
    .X(_05791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09057_ (.A(_05751_),
    .X(_05792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09058_ (.A1(_05790_),
    .A2(_05791_),
    .B1(\design_top.core0.REG1[9][15] ),
    .B2(_05792_),
    .X(_03707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09059_ (.A(_05653_),
    .X(_05793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09060_ (.A(_05793_),
    .X(_05794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09061_ (.A1(_05794_),
    .A2(_05791_),
    .B1(\design_top.core0.REG1[9][14] ),
    .B2(_05792_),
    .X(_03706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09062_ (.A1(\design_top.core0.REG1[9][13] ),
    .A2(_05748_),
    .B1(_05656_),
    .B2(_05752_),
    .X(_03705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09063_ (.A(_05657_),
    .X(_05795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09064_ (.A(_05795_),
    .X(_05796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09065_ (.A1(_05796_),
    .A2(_05791_),
    .B1(\design_top.core0.REG1[9][12] ),
    .B2(_05792_),
    .X(_03704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09066_ (.A(_05659_),
    .X(_05797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09067_ (.A(_05797_),
    .X(_05798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09068_ (.A1(_05798_),
    .A2(_05791_),
    .B1(\design_top.core0.REG1[9][11] ),
    .B2(_05792_),
    .X(_03703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09069_ (.A(_05662_),
    .X(_05799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09070_ (.A(_05799_),
    .X(_05800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09071_ (.A1(_05800_),
    .A2(_05791_),
    .B1(\design_top.core0.REG1[9][10] ),
    .B2(_05792_),
    .X(_03702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09072_ (.A(_05665_),
    .X(_05801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09073_ (.A(_05801_),
    .X(_05802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09074_ (.A(_05747_),
    .X(_05803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09075_ (.A(_05751_),
    .X(_05804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09076_ (.A1(_05802_),
    .A2(_05803_),
    .B1(\design_top.core0.REG1[9][9] ),
    .B2(_05804_),
    .X(_03701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09077_ (.A(_05668_),
    .X(_05805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09078_ (.A(_05805_),
    .X(_05806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09079_ (.A1(_05806_),
    .A2(_05803_),
    .B1(\design_top.core0.REG1[9][8] ),
    .B2(_05804_),
    .X(_03700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09080_ (.A(_05670_),
    .X(_05807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09081_ (.A(_05807_),
    .X(_05808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09082_ (.A1(_05808_),
    .A2(_05803_),
    .B1(\design_top.core0.REG1[9][7] ),
    .B2(_05804_),
    .X(_03699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09083_ (.A(_05672_),
    .X(_05809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09084_ (.A(_05809_),
    .X(_05810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09085_ (.A1(_05810_),
    .A2(_05803_),
    .B1(\design_top.core0.REG1[9][6] ),
    .B2(_05804_),
    .X(_03698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09086_ (.A(_05675_),
    .X(_05811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09087_ (.A(_05811_),
    .X(_05812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09088_ (.A1(_05812_),
    .A2(_05803_),
    .B1(\design_top.core0.REG1[9][5] ),
    .B2(_05804_),
    .X(_03697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09089_ (.A(_05678_),
    .X(_05813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09090_ (.A(_05813_),
    .X(_05814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09091_ (.A(_05747_),
    .X(_05815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09092_ (.A(_05751_),
    .X(_05816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09093_ (.A1(_05814_),
    .A2(_05815_),
    .B1(\design_top.core0.REG1[9][4] ),
    .B2(_05816_),
    .X(_03696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09094_ (.A(_05681_),
    .X(_05817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09095_ (.A(_05817_),
    .X(_05818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09096_ (.A1(_05818_),
    .A2(_05815_),
    .B1(\design_top.core0.REG1[9][3] ),
    .B2(_05816_),
    .X(_03695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09097_ (.A(_05683_),
    .X(_05819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09098_ (.A(_05819_),
    .X(_05820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09099_ (.A1(_05820_),
    .A2(_05815_),
    .B1(\design_top.core0.REG1[9][2] ),
    .B2(_05816_),
    .X(_03694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09100_ (.A(_05685_),
    .X(_05821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09101_ (.A(_05821_),
    .X(_05822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09102_ (.A1(_05822_),
    .A2(_05815_),
    .B1(\design_top.core0.REG1[9][1] ),
    .B2(_05816_),
    .X(_03693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09103_ (.A(_05687_),
    .X(_05823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09104_ (.A(_05823_),
    .X(_05824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09105_ (.A1(_05824_),
    .A2(_05815_),
    .B1(\design_top.core0.REG1[9][0] ),
    .B2(_05816_),
    .X(_03692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _09106_ (.A(_05108_),
    .B(_05737_),
    .Y(_00562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09107_ (.A(_05111_),
    .B(_00562_),
    .X(_05825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09108_ (.A(_05825_),
    .X(_05826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09109_ (.A(_05825_),
    .Y(_05827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09110_ (.A(_05827_),
    .X(_05828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09111_ (.A1(_00228_),
    .A2(_05826_),
    .B1(\design_top.MEM[15][7] ),
    .B2(_05828_),
    .X(_03691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09112_ (.A1(_00227_),
    .A2(_05826_),
    .B1(\design_top.MEM[15][6] ),
    .B2(_05828_),
    .X(_03690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09113_ (.A1(_00226_),
    .A2(_05826_),
    .B1(\design_top.MEM[15][5] ),
    .B2(_05828_),
    .X(_03689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09114_ (.A1(_00225_),
    .A2(_05826_),
    .B1(\design_top.MEM[15][4] ),
    .B2(_05828_),
    .X(_03688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09115_ (.A1(_00224_),
    .A2(_05826_),
    .B1(\design_top.MEM[15][3] ),
    .B2(_05828_),
    .X(_03687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09116_ (.A1(_00223_),
    .A2(_05825_),
    .B1(\design_top.MEM[15][2] ),
    .B2(_05827_),
    .X(_03686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09117_ (.A1(_00222_),
    .A2(_05825_),
    .B1(\design_top.MEM[15][1] ),
    .B2(_05827_),
    .X(_03685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09118_ (.A1(_00221_),
    .A2(_05825_),
    .B1(\design_top.MEM[15][0] ),
    .B2(_05827_),
    .X(_03684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _09119_ (.A(_05122_),
    .B(_05737_),
    .Y(_00561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09120_ (.A(_05125_),
    .B(_00561_),
    .X(_05829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09121_ (.A(_05829_),
    .X(_05830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09122_ (.A(_05829_),
    .Y(_05831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09123_ (.A(_05831_),
    .X(_05832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09124_ (.A1(_00236_),
    .A2(_05830_),
    .B1(\design_top.MEM[1][7] ),
    .B2(_05832_),
    .X(_03683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09125_ (.A1(_00235_),
    .A2(_05830_),
    .B1(\design_top.MEM[1][6] ),
    .B2(_05832_),
    .X(_03682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09126_ (.A1(_00234_),
    .A2(_05830_),
    .B1(\design_top.MEM[1][5] ),
    .B2(_05832_),
    .X(_03681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09127_ (.A1(_00233_),
    .A2(_05830_),
    .B1(\design_top.MEM[1][4] ),
    .B2(_05832_),
    .X(_03680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09128_ (.A1(_00232_),
    .A2(_05830_),
    .B1(\design_top.MEM[1][3] ),
    .B2(_05832_),
    .X(_03679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09129_ (.A1(_00231_),
    .A2(_05829_),
    .B1(\design_top.MEM[1][2] ),
    .B2(_05831_),
    .X(_03678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09130_ (.A1(_00230_),
    .A2(_05829_),
    .B1(\design_top.MEM[1][1] ),
    .B2(_05831_),
    .X(_03677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09131_ (.A1(_00229_),
    .A2(_05829_),
    .B1(\design_top.MEM[1][0] ),
    .B2(_05831_),
    .X(_03676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _09132_ (.A(_05136_),
    .B(_05737_),
    .Y(_00560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09133_ (.A(_05139_),
    .B(_00560_),
    .X(_05833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09134_ (.A(_05833_),
    .X(_05834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09135_ (.A(_05833_),
    .Y(_05835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09136_ (.A(_05835_),
    .X(_05836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09137_ (.A1(_00244_),
    .A2(_05834_),
    .B1(\design_top.MEM[2][7] ),
    .B2(_05836_),
    .X(_03675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09138_ (.A1(_00243_),
    .A2(_05834_),
    .B1(\design_top.MEM[2][6] ),
    .B2(_05836_),
    .X(_03674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09139_ (.A1(_00242_),
    .A2(_05834_),
    .B1(\design_top.MEM[2][5] ),
    .B2(_05836_),
    .X(_03673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09140_ (.A1(_00241_),
    .A2(_05834_),
    .B1(\design_top.MEM[2][4] ),
    .B2(_05836_),
    .X(_03672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09141_ (.A1(_00240_),
    .A2(_05834_),
    .B1(\design_top.MEM[2][3] ),
    .B2(_05836_),
    .X(_03671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09142_ (.A1(_00239_),
    .A2(_05833_),
    .B1(\design_top.MEM[2][2] ),
    .B2(_05835_),
    .X(_03670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09143_ (.A1(_00238_),
    .A2(_05833_),
    .B1(\design_top.MEM[2][1] ),
    .B2(_05835_),
    .X(_03669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09144_ (.A1(_00237_),
    .A2(_05833_),
    .B1(\design_top.MEM[2][0] ),
    .B2(_05835_),
    .X(_03668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _09145_ (.A(_05151_),
    .B(_05737_),
    .Y(_00559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09146_ (.A(_05154_),
    .B(_00559_),
    .X(_05837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09147_ (.A(_05837_),
    .X(_05838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09148_ (.A(_05837_),
    .Y(_05839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09149_ (.A(_05839_),
    .X(_05840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09150_ (.A1(_00252_),
    .A2(_05838_),
    .B1(\design_top.MEM[3][7] ),
    .B2(_05840_),
    .X(_03667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09151_ (.A1(_00251_),
    .A2(_05838_),
    .B1(\design_top.MEM[3][6] ),
    .B2(_05840_),
    .X(_03666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09152_ (.A1(_00250_),
    .A2(_05838_),
    .B1(\design_top.MEM[3][5] ),
    .B2(_05840_),
    .X(_03665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09153_ (.A1(_00249_),
    .A2(_05838_),
    .B1(\design_top.MEM[3][4] ),
    .B2(_05840_),
    .X(_03664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09154_ (.A1(_00248_),
    .A2(_05838_),
    .B1(\design_top.MEM[3][3] ),
    .B2(_05840_),
    .X(_03663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09155_ (.A1(_00247_),
    .A2(_05837_),
    .B1(\design_top.MEM[3][2] ),
    .B2(_05839_),
    .X(_03662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09156_ (.A1(_00246_),
    .A2(_05837_),
    .B1(\design_top.MEM[3][1] ),
    .B2(_05839_),
    .X(_03661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09157_ (.A1(_00245_),
    .A2(_05837_),
    .B1(\design_top.MEM[3][0] ),
    .B2(_05839_),
    .X(_03660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09158_ (.A(_05597_),
    .X(_05841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09159_ (.A(_01441_),
    .Y(_05842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09160_ (.A(_05842_),
    .X(_05843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09161_ (.A(_01440_),
    .Y(_05844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09162_ (.A(_05844_),
    .X(_05845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _09163_ (.A(_05841_),
    .B(_05843_),
    .C(_05845_),
    .D(_05595_),
    .X(_05846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09164_ (.A(_05746_),
    .B(_05846_),
    .X(_05847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09165_ (.A(_05847_),
    .X(_05848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09166_ (.A(_05848_),
    .X(_05849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09167_ (.A(_05847_),
    .Y(_05850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09168_ (.A(_05850_),
    .X(_05851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09169_ (.A(_05851_),
    .X(_05852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09170_ (.A1(\design_top.core0.REG1[15][31] ),
    .A2(_05849_),
    .B1(_05750_),
    .B2(_05852_),
    .X(_03659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09171_ (.A(_05753_),
    .X(_05853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09172_ (.A1(\design_top.core0.REG1[15][30] ),
    .A2(_05849_),
    .B1(_05853_),
    .B2(_05852_),
    .X(_03658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09173_ (.A(_05757_),
    .X(_05854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09174_ (.A1(\design_top.core0.REG1[15][29] ),
    .A2(_05849_),
    .B1(_05854_),
    .B2(_05852_),
    .X(_03657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09175_ (.A(_05759_),
    .X(_05855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09176_ (.A1(\design_top.core0.REG1[15][28] ),
    .A2(_05849_),
    .B1(_05855_),
    .B2(_05852_),
    .X(_03656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09177_ (.A(_05848_),
    .X(_05856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09178_ (.A(_05761_),
    .X(_05857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09179_ (.A1(\design_top.core0.REG1[15][27] ),
    .A2(_05856_),
    .B1(_05857_),
    .B2(_05852_),
    .X(_03655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09180_ (.A(_05763_),
    .X(_05858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09181_ (.A(_05851_),
    .X(_05859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09182_ (.A1(\design_top.core0.REG1[15][26] ),
    .A2(_05856_),
    .B1(_05858_),
    .B2(_05859_),
    .X(_03654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09183_ (.A(_05765_),
    .X(_05860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09184_ (.A1(\design_top.core0.REG1[15][25] ),
    .A2(_05856_),
    .B1(_05860_),
    .B2(_05859_),
    .X(_03653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09185_ (.A(_05769_),
    .X(_05861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09186_ (.A1(\design_top.core0.REG1[15][24] ),
    .A2(_05856_),
    .B1(_05861_),
    .B2(_05859_),
    .X(_03652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09187_ (.A(_05771_),
    .X(_05862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09188_ (.A1(\design_top.core0.REG1[15][23] ),
    .A2(_05856_),
    .B1(_05862_),
    .B2(_05859_),
    .X(_03651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09189_ (.A(_05848_),
    .X(_05863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09190_ (.A(_05773_),
    .X(_05864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09191_ (.A1(\design_top.core0.REG1[15][22] ),
    .A2(_05863_),
    .B1(_05864_),
    .B2(_05859_),
    .X(_03650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09192_ (.A(_05775_),
    .X(_05865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09193_ (.A(_05851_),
    .X(_05866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09194_ (.A1(\design_top.core0.REG1[15][21] ),
    .A2(_05863_),
    .B1(_05865_),
    .B2(_05866_),
    .X(_03649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09195_ (.A(_05777_),
    .X(_05867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09196_ (.A1(\design_top.core0.REG1[15][20] ),
    .A2(_05863_),
    .B1(_05867_),
    .B2(_05866_),
    .X(_03648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09197_ (.A(_05781_),
    .X(_05868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09198_ (.A1(\design_top.core0.REG1[15][19] ),
    .A2(_05863_),
    .B1(_05868_),
    .B2(_05866_),
    .X(_03647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09199_ (.A(_05783_),
    .X(_05869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09200_ (.A1(\design_top.core0.REG1[15][18] ),
    .A2(_05863_),
    .B1(_05869_),
    .B2(_05866_),
    .X(_03646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09201_ (.A(_05847_),
    .X(_05870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09202_ (.A(_05785_),
    .X(_05871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09203_ (.A1(\design_top.core0.REG1[15][17] ),
    .A2(_05870_),
    .B1(_05871_),
    .B2(_05866_),
    .X(_03645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09204_ (.A(_05787_),
    .X(_05872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09205_ (.A(_05850_),
    .X(_05873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09206_ (.A1(\design_top.core0.REG1[15][16] ),
    .A2(_05870_),
    .B1(_05872_),
    .B2(_05873_),
    .X(_03644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09207_ (.A(_05789_),
    .X(_05874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09208_ (.A1(\design_top.core0.REG1[15][15] ),
    .A2(_05870_),
    .B1(_05874_),
    .B2(_05873_),
    .X(_03643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09209_ (.A(_05793_),
    .X(_05875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09210_ (.A1(\design_top.core0.REG1[15][14] ),
    .A2(_05870_),
    .B1(_05875_),
    .B2(_05873_),
    .X(_03642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09211_ (.A(_00045_),
    .X(_05876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09212_ (.A1(\design_top.core0.REG1[15][13] ),
    .A2(_05851_),
    .B1(_05876_),
    .B2(_05849_),
    .X(_03641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09213_ (.A(_05795_),
    .X(_05877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09214_ (.A1(\design_top.core0.REG1[15][12] ),
    .A2(_05870_),
    .B1(_05877_),
    .B2(_05873_),
    .X(_03640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09215_ (.A(_05847_),
    .X(_05878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09216_ (.A(_05797_),
    .X(_05879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09217_ (.A1(\design_top.core0.REG1[15][11] ),
    .A2(_05878_),
    .B1(_05879_),
    .B2(_05873_),
    .X(_03639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09218_ (.A(_05799_),
    .X(_05880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09219_ (.A(_05850_),
    .X(_05881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09220_ (.A1(\design_top.core0.REG1[15][10] ),
    .A2(_05878_),
    .B1(_05880_),
    .B2(_05881_),
    .X(_03638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09221_ (.A(_05801_),
    .X(_05882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09222_ (.A1(\design_top.core0.REG1[15][9] ),
    .A2(_05878_),
    .B1(_05882_),
    .B2(_05881_),
    .X(_03637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09223_ (.A(_05805_),
    .X(_05883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09224_ (.A1(\design_top.core0.REG1[15][8] ),
    .A2(_05878_),
    .B1(_05883_),
    .B2(_05881_),
    .X(_03636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09225_ (.A(_05807_),
    .X(_05884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09226_ (.A1(\design_top.core0.REG1[15][7] ),
    .A2(_05878_),
    .B1(_05884_),
    .B2(_05881_),
    .X(_03635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09227_ (.A(_05847_),
    .X(_05885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09228_ (.A(_05809_),
    .X(_05886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09229_ (.A1(\design_top.core0.REG1[15][6] ),
    .A2(_05885_),
    .B1(_05886_),
    .B2(_05881_),
    .X(_03634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09230_ (.A(_05811_),
    .X(_05887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09231_ (.A(_05850_),
    .X(_05888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09232_ (.A1(\design_top.core0.REG1[15][5] ),
    .A2(_05885_),
    .B1(_05887_),
    .B2(_05888_),
    .X(_03633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09233_ (.A(_05813_),
    .X(_05889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09234_ (.A1(\design_top.core0.REG1[15][4] ),
    .A2(_05885_),
    .B1(_05889_),
    .B2(_05888_),
    .X(_03632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09235_ (.A(_05817_),
    .X(_05890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09236_ (.A1(\design_top.core0.REG1[15][3] ),
    .A2(_05885_),
    .B1(_05890_),
    .B2(_05888_),
    .X(_03631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09237_ (.A(_05819_),
    .X(_05891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09238_ (.A1(\design_top.core0.REG1[15][2] ),
    .A2(_05885_),
    .B1(_05891_),
    .B2(_05888_),
    .X(_03630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09239_ (.A(_05821_),
    .X(_05892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09240_ (.A1(\design_top.core0.REG1[15][1] ),
    .A2(_05848_),
    .B1(_05892_),
    .B2(_05888_),
    .X(_03629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09241_ (.A(_05823_),
    .X(_05893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09242_ (.A1(\design_top.core0.REG1[15][0] ),
    .A2(_05848_),
    .B1(_05893_),
    .B2(_05851_),
    .X(_03628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09243_ (.A(_01442_),
    .X(_05894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _09244_ (.A(_05594_),
    .B(_05596_),
    .C(_05894_),
    .D(_01441_),
    .X(_05895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09245_ (.A(_05746_),
    .B(_05895_),
    .X(_05896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09246_ (.A(_05896_),
    .X(_05897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09247_ (.A(_05897_),
    .X(_05898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09248_ (.A(_05896_),
    .Y(_05899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09249_ (.A(_05899_),
    .X(_05900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09250_ (.A(_05900_),
    .X(_05901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09251_ (.A1(\design_top.core0.REG1[1][31] ),
    .A2(_05898_),
    .B1(_05750_),
    .B2(_05901_),
    .X(_03627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09252_ (.A1(\design_top.core0.REG1[1][30] ),
    .A2(_05898_),
    .B1(_05853_),
    .B2(_05901_),
    .X(_03626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09253_ (.A1(\design_top.core0.REG1[1][29] ),
    .A2(_05898_),
    .B1(_05854_),
    .B2(_05901_),
    .X(_03625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09254_ (.A1(\design_top.core0.REG1[1][28] ),
    .A2(_05898_),
    .B1(_05855_),
    .B2(_05901_),
    .X(_03624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09255_ (.A(_05897_),
    .X(_05902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09256_ (.A1(\design_top.core0.REG1[1][27] ),
    .A2(_05902_),
    .B1(_05857_),
    .B2(_05901_),
    .X(_03623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09257_ (.A(_05900_),
    .X(_05903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09258_ (.A1(\design_top.core0.REG1[1][26] ),
    .A2(_05902_),
    .B1(_05858_),
    .B2(_05903_),
    .X(_03622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09259_ (.A1(\design_top.core0.REG1[1][25] ),
    .A2(_05902_),
    .B1(_05860_),
    .B2(_05903_),
    .X(_03621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09260_ (.A1(\design_top.core0.REG1[1][24] ),
    .A2(_05902_),
    .B1(_05861_),
    .B2(_05903_),
    .X(_03620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09261_ (.A1(\design_top.core0.REG1[1][23] ),
    .A2(_05902_),
    .B1(_05862_),
    .B2(_05903_),
    .X(_03619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09262_ (.A(_05897_),
    .X(_05904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09263_ (.A1(\design_top.core0.REG1[1][22] ),
    .A2(_05904_),
    .B1(_05864_),
    .B2(_05903_),
    .X(_03618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09264_ (.A(_05900_),
    .X(_05905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09265_ (.A1(\design_top.core0.REG1[1][21] ),
    .A2(_05904_),
    .B1(_05865_),
    .B2(_05905_),
    .X(_03617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09266_ (.A1(\design_top.core0.REG1[1][20] ),
    .A2(_05904_),
    .B1(_05867_),
    .B2(_05905_),
    .X(_03616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09267_ (.A1(\design_top.core0.REG1[1][19] ),
    .A2(_05904_),
    .B1(_05868_),
    .B2(_05905_),
    .X(_03615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09268_ (.A1(\design_top.core0.REG1[1][18] ),
    .A2(_05904_),
    .B1(_05869_),
    .B2(_05905_),
    .X(_03614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09269_ (.A(_05896_),
    .X(_05906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09270_ (.A1(\design_top.core0.REG1[1][17] ),
    .A2(_05906_),
    .B1(_05871_),
    .B2(_05905_),
    .X(_03613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09271_ (.A(_05899_),
    .X(_05907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09272_ (.A1(\design_top.core0.REG1[1][16] ),
    .A2(_05906_),
    .B1(_05872_),
    .B2(_05907_),
    .X(_03612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09273_ (.A1(\design_top.core0.REG1[1][15] ),
    .A2(_05906_),
    .B1(_05874_),
    .B2(_05907_),
    .X(_03611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09274_ (.A1(\design_top.core0.REG1[1][14] ),
    .A2(_05906_),
    .B1(_05875_),
    .B2(_05907_),
    .X(_03610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09275_ (.A1(\design_top.core0.REG1[1][13] ),
    .A2(_05900_),
    .B1(_05876_),
    .B2(_05898_),
    .X(_03609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09276_ (.A1(\design_top.core0.REG1[1][12] ),
    .A2(_05906_),
    .B1(_05877_),
    .B2(_05907_),
    .X(_03608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09277_ (.A(_05896_),
    .X(_05908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09278_ (.A1(\design_top.core0.REG1[1][11] ),
    .A2(_05908_),
    .B1(_05879_),
    .B2(_05907_),
    .X(_03607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09279_ (.A(_05899_),
    .X(_05909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09280_ (.A1(\design_top.core0.REG1[1][10] ),
    .A2(_05908_),
    .B1(_05880_),
    .B2(_05909_),
    .X(_03606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09281_ (.A1(\design_top.core0.REG1[1][9] ),
    .A2(_05908_),
    .B1(_05882_),
    .B2(_05909_),
    .X(_03605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09282_ (.A1(\design_top.core0.REG1[1][8] ),
    .A2(_05908_),
    .B1(_05883_),
    .B2(_05909_),
    .X(_03604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09283_ (.A1(\design_top.core0.REG1[1][7] ),
    .A2(_05908_),
    .B1(_05884_),
    .B2(_05909_),
    .X(_03603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09284_ (.A(_05896_),
    .X(_05910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09285_ (.A1(\design_top.core0.REG1[1][6] ),
    .A2(_05910_),
    .B1(_05886_),
    .B2(_05909_),
    .X(_03602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09286_ (.A(_05899_),
    .X(_05911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09287_ (.A1(\design_top.core0.REG1[1][5] ),
    .A2(_05910_),
    .B1(_05887_),
    .B2(_05911_),
    .X(_03601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09288_ (.A1(\design_top.core0.REG1[1][4] ),
    .A2(_05910_),
    .B1(_05889_),
    .B2(_05911_),
    .X(_03600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09289_ (.A1(\design_top.core0.REG1[1][3] ),
    .A2(_05910_),
    .B1(_05890_),
    .B2(_05911_),
    .X(_03599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09290_ (.A1(\design_top.core0.REG1[1][2] ),
    .A2(_05910_),
    .B1(_05891_),
    .B2(_05911_),
    .X(_03598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09291_ (.A1(\design_top.core0.REG1[1][1] ),
    .A2(_05897_),
    .B1(_05892_),
    .B2(_05911_),
    .X(_03597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09292_ (.A1(\design_top.core0.REG1[1][0] ),
    .A2(_05897_),
    .B1(_05893_),
    .B2(_05900_),
    .X(_03596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09293_ (.A(_01441_),
    .X(_05912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09294_ (.A(_01439_),
    .X(_05913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _09295_ (.A(_05894_),
    .B(_05912_),
    .C(_05845_),
    .D(_05913_),
    .X(_05914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09296_ (.A(_05746_),
    .B(_05914_),
    .X(_05915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09297_ (.A(_05915_),
    .X(_05916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09298_ (.A(_05916_),
    .X(_05917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09299_ (.A(_05915_),
    .Y(_05918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09300_ (.A(_05918_),
    .X(_05919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09301_ (.A(_05919_),
    .X(_05920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09302_ (.A1(\design_top.core0.REG1[2][31] ),
    .A2(_05917_),
    .B1(_05750_),
    .B2(_05920_),
    .X(_03595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09303_ (.A1(\design_top.core0.REG1[2][30] ),
    .A2(_05917_),
    .B1(_05853_),
    .B2(_05920_),
    .X(_03594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09304_ (.A1(\design_top.core0.REG1[2][29] ),
    .A2(_05917_),
    .B1(_05854_),
    .B2(_05920_),
    .X(_03593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09305_ (.A1(\design_top.core0.REG1[2][28] ),
    .A2(_05917_),
    .B1(_05855_),
    .B2(_05920_),
    .X(_03592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09306_ (.A(_05916_),
    .X(_05921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09307_ (.A1(\design_top.core0.REG1[2][27] ),
    .A2(_05921_),
    .B1(_05857_),
    .B2(_05920_),
    .X(_03591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09308_ (.A(_05919_),
    .X(_05922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09309_ (.A1(\design_top.core0.REG1[2][26] ),
    .A2(_05921_),
    .B1(_05858_),
    .B2(_05922_),
    .X(_03590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09310_ (.A1(\design_top.core0.REG1[2][25] ),
    .A2(_05921_),
    .B1(_05860_),
    .B2(_05922_),
    .X(_03589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09311_ (.A1(\design_top.core0.REG1[2][24] ),
    .A2(_05921_),
    .B1(_05861_),
    .B2(_05922_),
    .X(_03588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09312_ (.A1(\design_top.core0.REG1[2][23] ),
    .A2(_05921_),
    .B1(_05862_),
    .B2(_05922_),
    .X(_03587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09313_ (.A(_05916_),
    .X(_05923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09314_ (.A1(\design_top.core0.REG1[2][22] ),
    .A2(_05923_),
    .B1(_05864_),
    .B2(_05922_),
    .X(_03586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09315_ (.A(_05919_),
    .X(_05924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09316_ (.A1(\design_top.core0.REG1[2][21] ),
    .A2(_05923_),
    .B1(_05865_),
    .B2(_05924_),
    .X(_03585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09317_ (.A1(\design_top.core0.REG1[2][20] ),
    .A2(_05923_),
    .B1(_05867_),
    .B2(_05924_),
    .X(_03584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09318_ (.A1(\design_top.core0.REG1[2][19] ),
    .A2(_05923_),
    .B1(_05868_),
    .B2(_05924_),
    .X(_03583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09319_ (.A1(\design_top.core0.REG1[2][18] ),
    .A2(_05923_),
    .B1(_05869_),
    .B2(_05924_),
    .X(_03582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09320_ (.A(_05915_),
    .X(_05925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09321_ (.A1(\design_top.core0.REG1[2][17] ),
    .A2(_05925_),
    .B1(_05871_),
    .B2(_05924_),
    .X(_03581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09322_ (.A(_05918_),
    .X(_05926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09323_ (.A1(\design_top.core0.REG1[2][16] ),
    .A2(_05925_),
    .B1(_05872_),
    .B2(_05926_),
    .X(_03580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09324_ (.A1(\design_top.core0.REG1[2][15] ),
    .A2(_05925_),
    .B1(_05874_),
    .B2(_05926_),
    .X(_03579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09325_ (.A1(\design_top.core0.REG1[2][14] ),
    .A2(_05925_),
    .B1(_05875_),
    .B2(_05926_),
    .X(_03578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09326_ (.A1(\design_top.core0.REG1[2][13] ),
    .A2(_05919_),
    .B1(_05876_),
    .B2(_05917_),
    .X(_03577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09327_ (.A1(\design_top.core0.REG1[2][12] ),
    .A2(_05925_),
    .B1(_05877_),
    .B2(_05926_),
    .X(_03576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09328_ (.A(_05915_),
    .X(_05927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09329_ (.A1(\design_top.core0.REG1[2][11] ),
    .A2(_05927_),
    .B1(_05879_),
    .B2(_05926_),
    .X(_03575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09330_ (.A(_05918_),
    .X(_05928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09331_ (.A1(\design_top.core0.REG1[2][10] ),
    .A2(_05927_),
    .B1(_05880_),
    .B2(_05928_),
    .X(_03574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09332_ (.A1(\design_top.core0.REG1[2][9] ),
    .A2(_05927_),
    .B1(_05882_),
    .B2(_05928_),
    .X(_03573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09333_ (.A1(\design_top.core0.REG1[2][8] ),
    .A2(_05927_),
    .B1(_05883_),
    .B2(_05928_),
    .X(_03572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09334_ (.A1(\design_top.core0.REG1[2][7] ),
    .A2(_05927_),
    .B1(_05884_),
    .B2(_05928_),
    .X(_03571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09335_ (.A(_05915_),
    .X(_05929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09336_ (.A1(\design_top.core0.REG1[2][6] ),
    .A2(_05929_),
    .B1(_05886_),
    .B2(_05928_),
    .X(_03570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09337_ (.A(_05918_),
    .X(_05930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09338_ (.A1(\design_top.core0.REG1[2][5] ),
    .A2(_05929_),
    .B1(_05887_),
    .B2(_05930_),
    .X(_03569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09339_ (.A1(\design_top.core0.REG1[2][4] ),
    .A2(_05929_),
    .B1(_05889_),
    .B2(_05930_),
    .X(_03568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09340_ (.A1(\design_top.core0.REG1[2][3] ),
    .A2(_05929_),
    .B1(_05890_),
    .B2(_05930_),
    .X(_03567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09341_ (.A1(\design_top.core0.REG1[2][2] ),
    .A2(_05929_),
    .B1(_05891_),
    .B2(_05930_),
    .X(_03566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09342_ (.A1(\design_top.core0.REG1[2][1] ),
    .A2(_05916_),
    .B1(_05892_),
    .B2(_05930_),
    .X(_03565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09343_ (.A1(\design_top.core0.REG1[2][0] ),
    .A2(_05916_),
    .B1(_05893_),
    .B2(_05919_),
    .X(_03564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09344_ (.A(_05745_),
    .X(_05931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _09345_ (.A(_05894_),
    .B(_05912_),
    .C(_05845_),
    .D(_05595_),
    .X(_05932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09346_ (.A(_05931_),
    .B(_05932_),
    .X(_05933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09347_ (.A(_05933_),
    .X(_05934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09348_ (.A(_05934_),
    .X(_05935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09349_ (.A(_05933_),
    .Y(_05936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09350_ (.A(_05936_),
    .X(_05937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09351_ (.A(_05937_),
    .X(_05938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09352_ (.A1(\design_top.core0.REG1[3][31] ),
    .A2(_05935_),
    .B1(_05750_),
    .B2(_05938_),
    .X(_03563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09353_ (.A1(\design_top.core0.REG1[3][30] ),
    .A2(_05935_),
    .B1(_05853_),
    .B2(_05938_),
    .X(_03562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09354_ (.A1(\design_top.core0.REG1[3][29] ),
    .A2(_05935_),
    .B1(_05854_),
    .B2(_05938_),
    .X(_03561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09355_ (.A1(\design_top.core0.REG1[3][28] ),
    .A2(_05935_),
    .B1(_05855_),
    .B2(_05938_),
    .X(_03560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09356_ (.A(_05934_),
    .X(_05939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09357_ (.A1(\design_top.core0.REG1[3][27] ),
    .A2(_05939_),
    .B1(_05857_),
    .B2(_05938_),
    .X(_03559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09358_ (.A(_05937_),
    .X(_05940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09359_ (.A1(\design_top.core0.REG1[3][26] ),
    .A2(_05939_),
    .B1(_05858_),
    .B2(_05940_),
    .X(_03558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09360_ (.A1(\design_top.core0.REG1[3][25] ),
    .A2(_05939_),
    .B1(_05860_),
    .B2(_05940_),
    .X(_03557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09361_ (.A1(\design_top.core0.REG1[3][24] ),
    .A2(_05939_),
    .B1(_05861_),
    .B2(_05940_),
    .X(_03556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09362_ (.A1(\design_top.core0.REG1[3][23] ),
    .A2(_05939_),
    .B1(_05862_),
    .B2(_05940_),
    .X(_03555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09363_ (.A(_05934_),
    .X(_05941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09364_ (.A1(\design_top.core0.REG1[3][22] ),
    .A2(_05941_),
    .B1(_05864_),
    .B2(_05940_),
    .X(_03554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09365_ (.A(_05937_),
    .X(_05942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09366_ (.A1(\design_top.core0.REG1[3][21] ),
    .A2(_05941_),
    .B1(_05865_),
    .B2(_05942_),
    .X(_03553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09367_ (.A1(\design_top.core0.REG1[3][20] ),
    .A2(_05941_),
    .B1(_05867_),
    .B2(_05942_),
    .X(_03552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09368_ (.A1(\design_top.core0.REG1[3][19] ),
    .A2(_05941_),
    .B1(_05868_),
    .B2(_05942_),
    .X(_03551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09369_ (.A1(\design_top.core0.REG1[3][18] ),
    .A2(_05941_),
    .B1(_05869_),
    .B2(_05942_),
    .X(_03550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09370_ (.A(_05933_),
    .X(_05943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09371_ (.A1(\design_top.core0.REG1[3][17] ),
    .A2(_05943_),
    .B1(_05871_),
    .B2(_05942_),
    .X(_03549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09372_ (.A(_05936_),
    .X(_05944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09373_ (.A1(\design_top.core0.REG1[3][16] ),
    .A2(_05943_),
    .B1(_05872_),
    .B2(_05944_),
    .X(_03548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09374_ (.A1(\design_top.core0.REG1[3][15] ),
    .A2(_05943_),
    .B1(_05874_),
    .B2(_05944_),
    .X(_03547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09375_ (.A1(\design_top.core0.REG1[3][14] ),
    .A2(_05943_),
    .B1(_05875_),
    .B2(_05944_),
    .X(_03546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09376_ (.A(_00045_),
    .X(_05945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09377_ (.A1(\design_top.core0.REG1[3][13] ),
    .A2(_05937_),
    .B1(_05945_),
    .B2(_05935_),
    .X(_03545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09378_ (.A1(\design_top.core0.REG1[3][12] ),
    .A2(_05943_),
    .B1(_05877_),
    .B2(_05944_),
    .X(_03544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09379_ (.A(_05933_),
    .X(_05946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09380_ (.A1(\design_top.core0.REG1[3][11] ),
    .A2(_05946_),
    .B1(_05879_),
    .B2(_05944_),
    .X(_03543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09381_ (.A(_05936_),
    .X(_05947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09382_ (.A1(\design_top.core0.REG1[3][10] ),
    .A2(_05946_),
    .B1(_05880_),
    .B2(_05947_),
    .X(_03542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09383_ (.A1(\design_top.core0.REG1[3][9] ),
    .A2(_05946_),
    .B1(_05882_),
    .B2(_05947_),
    .X(_03541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09384_ (.A1(\design_top.core0.REG1[3][8] ),
    .A2(_05946_),
    .B1(_05883_),
    .B2(_05947_),
    .X(_03540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09385_ (.A1(\design_top.core0.REG1[3][7] ),
    .A2(_05946_),
    .B1(_05884_),
    .B2(_05947_),
    .X(_03539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09386_ (.A(_05933_),
    .X(_05948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09387_ (.A1(\design_top.core0.REG1[3][6] ),
    .A2(_05948_),
    .B1(_05886_),
    .B2(_05947_),
    .X(_03538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09388_ (.A(_05936_),
    .X(_05949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09389_ (.A1(\design_top.core0.REG1[3][5] ),
    .A2(_05948_),
    .B1(_05887_),
    .B2(_05949_),
    .X(_03537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09390_ (.A1(\design_top.core0.REG1[3][4] ),
    .A2(_05948_),
    .B1(_05889_),
    .B2(_05949_),
    .X(_03536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09391_ (.A1(\design_top.core0.REG1[3][3] ),
    .A2(_05948_),
    .B1(_05890_),
    .B2(_05949_),
    .X(_03535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09392_ (.A1(\design_top.core0.REG1[3][2] ),
    .A2(_05948_),
    .B1(_05891_),
    .B2(_05949_),
    .X(_03534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09393_ (.A1(\design_top.core0.REG1[3][1] ),
    .A2(_05934_),
    .B1(_05892_),
    .B2(_05949_),
    .X(_03533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09394_ (.A1(\design_top.core0.REG1[3][0] ),
    .A2(_05934_),
    .B1(_05893_),
    .B2(_05937_),
    .X(_03532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _09395_ (.A(_05594_),
    .B(_05913_),
    .C(_05894_),
    .D(_05843_),
    .X(_05950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09396_ (.A(_05931_),
    .B(_05950_),
    .X(_05951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09397_ (.A(_05951_),
    .X(_05952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09398_ (.A(_05952_),
    .X(_05953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09399_ (.A(_05749_),
    .X(_05954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09400_ (.A(_05951_),
    .Y(_05955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09401_ (.A(_05955_),
    .X(_05956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09402_ (.A(_05956_),
    .X(_05957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09403_ (.A1(\design_top.core0.REG1[4][31] ),
    .A2(_05953_),
    .B1(_05954_),
    .B2(_05957_),
    .X(_03531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09404_ (.A1(\design_top.core0.REG1[4][30] ),
    .A2(_05953_),
    .B1(_05853_),
    .B2(_05957_),
    .X(_03530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09405_ (.A1(\design_top.core0.REG1[4][29] ),
    .A2(_05953_),
    .B1(_05854_),
    .B2(_05957_),
    .X(_03529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09406_ (.A1(\design_top.core0.REG1[4][28] ),
    .A2(_05953_),
    .B1(_05855_),
    .B2(_05957_),
    .X(_03528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09407_ (.A(_05952_),
    .X(_05958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09408_ (.A1(\design_top.core0.REG1[4][27] ),
    .A2(_05958_),
    .B1(_05857_),
    .B2(_05957_),
    .X(_03527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09409_ (.A(_05956_),
    .X(_05959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09410_ (.A1(\design_top.core0.REG1[4][26] ),
    .A2(_05958_),
    .B1(_05858_),
    .B2(_05959_),
    .X(_03526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09411_ (.A1(\design_top.core0.REG1[4][25] ),
    .A2(_05958_),
    .B1(_05860_),
    .B2(_05959_),
    .X(_03525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09412_ (.A1(\design_top.core0.REG1[4][24] ),
    .A2(_05958_),
    .B1(_05861_),
    .B2(_05959_),
    .X(_03524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09413_ (.A1(\design_top.core0.REG1[4][23] ),
    .A2(_05958_),
    .B1(_05862_),
    .B2(_05959_),
    .X(_03523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09414_ (.A(_05952_),
    .X(_05960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09415_ (.A1(\design_top.core0.REG1[4][22] ),
    .A2(_05960_),
    .B1(_05864_),
    .B2(_05959_),
    .X(_03522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09416_ (.A(_05956_),
    .X(_05961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09417_ (.A1(\design_top.core0.REG1[4][21] ),
    .A2(_05960_),
    .B1(_05865_),
    .B2(_05961_),
    .X(_03521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09418_ (.A1(\design_top.core0.REG1[4][20] ),
    .A2(_05960_),
    .B1(_05867_),
    .B2(_05961_),
    .X(_03520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09419_ (.A1(\design_top.core0.REG1[4][19] ),
    .A2(_05960_),
    .B1(_05868_),
    .B2(_05961_),
    .X(_03519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09420_ (.A1(\design_top.core0.REG1[4][18] ),
    .A2(_05960_),
    .B1(_05869_),
    .B2(_05961_),
    .X(_03518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09421_ (.A(_05951_),
    .X(_05962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09422_ (.A1(\design_top.core0.REG1[4][17] ),
    .A2(_05962_),
    .B1(_05871_),
    .B2(_05961_),
    .X(_03517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09423_ (.A(_05955_),
    .X(_05963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09424_ (.A1(\design_top.core0.REG1[4][16] ),
    .A2(_05962_),
    .B1(_05872_),
    .B2(_05963_),
    .X(_03516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09425_ (.A1(\design_top.core0.REG1[4][15] ),
    .A2(_05962_),
    .B1(_05874_),
    .B2(_05963_),
    .X(_03515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09426_ (.A1(\design_top.core0.REG1[4][14] ),
    .A2(_05962_),
    .B1(_05875_),
    .B2(_05963_),
    .X(_03514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09427_ (.A1(\design_top.core0.REG1[4][13] ),
    .A2(_05956_),
    .B1(_05945_),
    .B2(_05953_),
    .X(_03513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09428_ (.A1(\design_top.core0.REG1[4][12] ),
    .A2(_05962_),
    .B1(_05877_),
    .B2(_05963_),
    .X(_03512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09429_ (.A(_05951_),
    .X(_05964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09430_ (.A1(\design_top.core0.REG1[4][11] ),
    .A2(_05964_),
    .B1(_05879_),
    .B2(_05963_),
    .X(_03511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09431_ (.A(_05955_),
    .X(_05965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09432_ (.A1(\design_top.core0.REG1[4][10] ),
    .A2(_05964_),
    .B1(_05880_),
    .B2(_05965_),
    .X(_03510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09433_ (.A1(\design_top.core0.REG1[4][9] ),
    .A2(_05964_),
    .B1(_05882_),
    .B2(_05965_),
    .X(_03509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09434_ (.A1(\design_top.core0.REG1[4][8] ),
    .A2(_05964_),
    .B1(_05883_),
    .B2(_05965_),
    .X(_03508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09435_ (.A1(\design_top.core0.REG1[4][7] ),
    .A2(_05964_),
    .B1(_05884_),
    .B2(_05965_),
    .X(_03507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09436_ (.A(_05951_),
    .X(_05966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09437_ (.A1(\design_top.core0.REG1[4][6] ),
    .A2(_05966_),
    .B1(_05886_),
    .B2(_05965_),
    .X(_03506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09438_ (.A(_05955_),
    .X(_05967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09439_ (.A1(\design_top.core0.REG1[4][5] ),
    .A2(_05966_),
    .B1(_05887_),
    .B2(_05967_),
    .X(_03505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09440_ (.A1(\design_top.core0.REG1[4][4] ),
    .A2(_05966_),
    .B1(_05889_),
    .B2(_05967_),
    .X(_03504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09441_ (.A1(\design_top.core0.REG1[4][3] ),
    .A2(_05966_),
    .B1(_05890_),
    .B2(_05967_),
    .X(_03503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09442_ (.A1(\design_top.core0.REG1[4][2] ),
    .A2(_05966_),
    .B1(_05891_),
    .B2(_05967_),
    .X(_03502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09443_ (.A1(\design_top.core0.REG1[4][1] ),
    .A2(_05952_),
    .B1(_05892_),
    .B2(_05967_),
    .X(_03501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09444_ (.A1(\design_top.core0.REG1[4][0] ),
    .A2(_05952_),
    .B1(_05893_),
    .B2(_05956_),
    .X(_03500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _09445_ (.A(_05594_),
    .B(_05596_),
    .C(_05894_),
    .D(_05843_),
    .X(_05968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09446_ (.A(_05931_),
    .B(_05968_),
    .X(_05969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09447_ (.A(_05969_),
    .X(_05970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09448_ (.A(_05970_),
    .X(_05971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09449_ (.A(_05969_),
    .Y(_05972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09450_ (.A(_05972_),
    .X(_05973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09451_ (.A(_05973_),
    .X(_05974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09452_ (.A1(\design_top.core0.REG1[5][31] ),
    .A2(_05971_),
    .B1(_05954_),
    .B2(_05974_),
    .X(_03499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09453_ (.A(_05753_),
    .X(_05975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09454_ (.A1(\design_top.core0.REG1[5][30] ),
    .A2(_05971_),
    .B1(_05975_),
    .B2(_05974_),
    .X(_03498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09455_ (.A(_05757_),
    .X(_05976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09456_ (.A1(\design_top.core0.REG1[5][29] ),
    .A2(_05971_),
    .B1(_05976_),
    .B2(_05974_),
    .X(_03497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09457_ (.A(_05759_),
    .X(_05977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09458_ (.A1(\design_top.core0.REG1[5][28] ),
    .A2(_05971_),
    .B1(_05977_),
    .B2(_05974_),
    .X(_03496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09459_ (.A(_05970_),
    .X(_05978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09460_ (.A(_05761_),
    .X(_05979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09461_ (.A1(\design_top.core0.REG1[5][27] ),
    .A2(_05978_),
    .B1(_05979_),
    .B2(_05974_),
    .X(_03495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09462_ (.A(_05763_),
    .X(_05980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09463_ (.A(_05973_),
    .X(_05981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09464_ (.A1(\design_top.core0.REG1[5][26] ),
    .A2(_05978_),
    .B1(_05980_),
    .B2(_05981_),
    .X(_03494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09465_ (.A(_05765_),
    .X(_05982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09466_ (.A1(\design_top.core0.REG1[5][25] ),
    .A2(_05978_),
    .B1(_05982_),
    .B2(_05981_),
    .X(_03493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09467_ (.A(_05769_),
    .X(_05983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09468_ (.A1(\design_top.core0.REG1[5][24] ),
    .A2(_05978_),
    .B1(_05983_),
    .B2(_05981_),
    .X(_03492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09469_ (.A(_05771_),
    .X(_05984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09470_ (.A1(\design_top.core0.REG1[5][23] ),
    .A2(_05978_),
    .B1(_05984_),
    .B2(_05981_),
    .X(_03491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09471_ (.A(_05970_),
    .X(_05985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09472_ (.A(_05773_),
    .X(_05986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09473_ (.A1(\design_top.core0.REG1[5][22] ),
    .A2(_05985_),
    .B1(_05986_),
    .B2(_05981_),
    .X(_03490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09474_ (.A(_05775_),
    .X(_05987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09475_ (.A(_05973_),
    .X(_05988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09476_ (.A1(\design_top.core0.REG1[5][21] ),
    .A2(_05985_),
    .B1(_05987_),
    .B2(_05988_),
    .X(_03489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09477_ (.A(_05777_),
    .X(_05989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09478_ (.A1(\design_top.core0.REG1[5][20] ),
    .A2(_05985_),
    .B1(_05989_),
    .B2(_05988_),
    .X(_03488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09479_ (.A(_05781_),
    .X(_05990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09480_ (.A1(\design_top.core0.REG1[5][19] ),
    .A2(_05985_),
    .B1(_05990_),
    .B2(_05988_),
    .X(_03487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09481_ (.A(_05783_),
    .X(_05991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09482_ (.A1(\design_top.core0.REG1[5][18] ),
    .A2(_05985_),
    .B1(_05991_),
    .B2(_05988_),
    .X(_03486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09483_ (.A(_05969_),
    .X(_05992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09484_ (.A(_05785_),
    .X(_05993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09485_ (.A1(\design_top.core0.REG1[5][17] ),
    .A2(_05992_),
    .B1(_05993_),
    .B2(_05988_),
    .X(_03485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09486_ (.A(_05787_),
    .X(_05994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09487_ (.A(_05972_),
    .X(_05995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09488_ (.A1(\design_top.core0.REG1[5][16] ),
    .A2(_05992_),
    .B1(_05994_),
    .B2(_05995_),
    .X(_03484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09489_ (.A(_05789_),
    .X(_05996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09490_ (.A1(\design_top.core0.REG1[5][15] ),
    .A2(_05992_),
    .B1(_05996_),
    .B2(_05995_),
    .X(_03483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09491_ (.A(_05793_),
    .X(_05997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09492_ (.A1(\design_top.core0.REG1[5][14] ),
    .A2(_05992_),
    .B1(_05997_),
    .B2(_05995_),
    .X(_03482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09493_ (.A1(\design_top.core0.REG1[5][13] ),
    .A2(_05973_),
    .B1(_05945_),
    .B2(_05971_),
    .X(_03481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09494_ (.A(_05795_),
    .X(_05998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09495_ (.A1(\design_top.core0.REG1[5][12] ),
    .A2(_05992_),
    .B1(_05998_),
    .B2(_05995_),
    .X(_03480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09496_ (.A(_05969_),
    .X(_05999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09497_ (.A(_05797_),
    .X(_06000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09498_ (.A1(\design_top.core0.REG1[5][11] ),
    .A2(_05999_),
    .B1(_06000_),
    .B2(_05995_),
    .X(_03479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09499_ (.A(_05799_),
    .X(_06001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09500_ (.A(_05972_),
    .X(_06002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09501_ (.A1(\design_top.core0.REG1[5][10] ),
    .A2(_05999_),
    .B1(_06001_),
    .B2(_06002_),
    .X(_03478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09502_ (.A(_05801_),
    .X(_06003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09503_ (.A1(\design_top.core0.REG1[5][9] ),
    .A2(_05999_),
    .B1(_06003_),
    .B2(_06002_),
    .X(_03477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09504_ (.A(_05805_),
    .X(_06004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09505_ (.A1(\design_top.core0.REG1[5][8] ),
    .A2(_05999_),
    .B1(_06004_),
    .B2(_06002_),
    .X(_03476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09506_ (.A(_05807_),
    .X(_06005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09507_ (.A1(\design_top.core0.REG1[5][7] ),
    .A2(_05999_),
    .B1(_06005_),
    .B2(_06002_),
    .X(_03475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09508_ (.A(_05969_),
    .X(_06006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09509_ (.A(_05809_),
    .X(_06007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09510_ (.A1(\design_top.core0.REG1[5][6] ),
    .A2(_06006_),
    .B1(_06007_),
    .B2(_06002_),
    .X(_03474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09511_ (.A(_05811_),
    .X(_06008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09512_ (.A(_05972_),
    .X(_06009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09513_ (.A1(\design_top.core0.REG1[5][5] ),
    .A2(_06006_),
    .B1(_06008_),
    .B2(_06009_),
    .X(_03473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09514_ (.A(_05813_),
    .X(_06010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09515_ (.A1(\design_top.core0.REG1[5][4] ),
    .A2(_06006_),
    .B1(_06010_),
    .B2(_06009_),
    .X(_03472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09516_ (.A(_05817_),
    .X(_06011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09517_ (.A1(\design_top.core0.REG1[5][3] ),
    .A2(_06006_),
    .B1(_06011_),
    .B2(_06009_),
    .X(_03471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09518_ (.A(_05819_),
    .X(_06012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09519_ (.A1(\design_top.core0.REG1[5][2] ),
    .A2(_06006_),
    .B1(_06012_),
    .B2(_06009_),
    .X(_03470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09520_ (.A(_05821_),
    .X(_06013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09521_ (.A1(\design_top.core0.REG1[5][1] ),
    .A2(_05970_),
    .B1(_06013_),
    .B2(_06009_),
    .X(_03469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09522_ (.A(_05823_),
    .X(_06014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09523_ (.A1(\design_top.core0.REG1[5][0] ),
    .A2(_05970_),
    .B1(_06014_),
    .B2(_05973_),
    .X(_03468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _09524_ (.A(_05845_),
    .B(_05913_),
    .C(_01442_),
    .D(_05843_),
    .X(_06015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09525_ (.A(_05931_),
    .B(_06015_),
    .X(_06016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09526_ (.A(_06016_),
    .X(_06017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09527_ (.A(_06017_),
    .X(_06018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09528_ (.A(_06016_),
    .Y(_06019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09529_ (.A(_06019_),
    .X(_06020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09530_ (.A(_06020_),
    .X(_06021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09531_ (.A1(\design_top.core0.REG1[6][31] ),
    .A2(_06018_),
    .B1(_05954_),
    .B2(_06021_),
    .X(_03467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09532_ (.A1(\design_top.core0.REG1[6][30] ),
    .A2(_06018_),
    .B1(_05975_),
    .B2(_06021_),
    .X(_03466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09533_ (.A1(\design_top.core0.REG1[6][29] ),
    .A2(_06018_),
    .B1(_05976_),
    .B2(_06021_),
    .X(_03465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09534_ (.A1(\design_top.core0.REG1[6][28] ),
    .A2(_06018_),
    .B1(_05977_),
    .B2(_06021_),
    .X(_03464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09535_ (.A(_06017_),
    .X(_06022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09536_ (.A1(\design_top.core0.REG1[6][27] ),
    .A2(_06022_),
    .B1(_05979_),
    .B2(_06021_),
    .X(_03463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09537_ (.A(_06020_),
    .X(_06023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09538_ (.A1(\design_top.core0.REG1[6][26] ),
    .A2(_06022_),
    .B1(_05980_),
    .B2(_06023_),
    .X(_03462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09539_ (.A1(\design_top.core0.REG1[6][25] ),
    .A2(_06022_),
    .B1(_05982_),
    .B2(_06023_),
    .X(_03461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09540_ (.A1(\design_top.core0.REG1[6][24] ),
    .A2(_06022_),
    .B1(_05983_),
    .B2(_06023_),
    .X(_03460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09541_ (.A1(\design_top.core0.REG1[6][23] ),
    .A2(_06022_),
    .B1(_05984_),
    .B2(_06023_),
    .X(_03459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09542_ (.A(_06017_),
    .X(_06024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09543_ (.A1(\design_top.core0.REG1[6][22] ),
    .A2(_06024_),
    .B1(_05986_),
    .B2(_06023_),
    .X(_03458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09544_ (.A(_06020_),
    .X(_06025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09545_ (.A1(\design_top.core0.REG1[6][21] ),
    .A2(_06024_),
    .B1(_05987_),
    .B2(_06025_),
    .X(_03457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09546_ (.A1(\design_top.core0.REG1[6][20] ),
    .A2(_06024_),
    .B1(_05989_),
    .B2(_06025_),
    .X(_03456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09547_ (.A1(\design_top.core0.REG1[6][19] ),
    .A2(_06024_),
    .B1(_05990_),
    .B2(_06025_),
    .X(_03455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09548_ (.A1(\design_top.core0.REG1[6][18] ),
    .A2(_06024_),
    .B1(_05991_),
    .B2(_06025_),
    .X(_03454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09549_ (.A(_06016_),
    .X(_06026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09550_ (.A1(\design_top.core0.REG1[6][17] ),
    .A2(_06026_),
    .B1(_05993_),
    .B2(_06025_),
    .X(_03453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09551_ (.A(_06019_),
    .X(_06027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09552_ (.A1(\design_top.core0.REG1[6][16] ),
    .A2(_06026_),
    .B1(_05994_),
    .B2(_06027_),
    .X(_03452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09553_ (.A1(\design_top.core0.REG1[6][15] ),
    .A2(_06026_),
    .B1(_05996_),
    .B2(_06027_),
    .X(_03451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09554_ (.A1(\design_top.core0.REG1[6][14] ),
    .A2(_06026_),
    .B1(_05997_),
    .B2(_06027_),
    .X(_03450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09555_ (.A1(\design_top.core0.REG1[6][13] ),
    .A2(_06020_),
    .B1(_05945_),
    .B2(_06018_),
    .X(_03449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09556_ (.A1(\design_top.core0.REG1[6][12] ),
    .A2(_06026_),
    .B1(_05998_),
    .B2(_06027_),
    .X(_03448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09557_ (.A(_06016_),
    .X(_06028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09558_ (.A1(\design_top.core0.REG1[6][11] ),
    .A2(_06028_),
    .B1(_06000_),
    .B2(_06027_),
    .X(_03447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09559_ (.A(_06019_),
    .X(_06029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09560_ (.A1(\design_top.core0.REG1[6][10] ),
    .A2(_06028_),
    .B1(_06001_),
    .B2(_06029_),
    .X(_03446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09561_ (.A1(\design_top.core0.REG1[6][9] ),
    .A2(_06028_),
    .B1(_06003_),
    .B2(_06029_),
    .X(_03445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09562_ (.A1(\design_top.core0.REG1[6][8] ),
    .A2(_06028_),
    .B1(_06004_),
    .B2(_06029_),
    .X(_03444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09563_ (.A1(\design_top.core0.REG1[6][7] ),
    .A2(_06028_),
    .B1(_06005_),
    .B2(_06029_),
    .X(_03443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09564_ (.A(_06016_),
    .X(_06030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09565_ (.A1(\design_top.core0.REG1[6][6] ),
    .A2(_06030_),
    .B1(_06007_),
    .B2(_06029_),
    .X(_03442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09566_ (.A(_06019_),
    .X(_06031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09567_ (.A1(\design_top.core0.REG1[6][5] ),
    .A2(_06030_),
    .B1(_06008_),
    .B2(_06031_),
    .X(_03441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09568_ (.A1(\design_top.core0.REG1[6][4] ),
    .A2(_06030_),
    .B1(_06010_),
    .B2(_06031_),
    .X(_03440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09569_ (.A1(\design_top.core0.REG1[6][3] ),
    .A2(_06030_),
    .B1(_06011_),
    .B2(_06031_),
    .X(_03439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09570_ (.A1(\design_top.core0.REG1[6][2] ),
    .A2(_06030_),
    .B1(_06012_),
    .B2(_06031_),
    .X(_03438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09571_ (.A1(\design_top.core0.REG1[6][1] ),
    .A2(_06017_),
    .B1(_06013_),
    .B2(_06031_),
    .X(_03437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09572_ (.A1(\design_top.core0.REG1[6][0] ),
    .A2(_06017_),
    .B1(_06014_),
    .B2(_06020_),
    .X(_03436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _09573_ (.A(_05845_),
    .B(_05596_),
    .C(_01442_),
    .D(_05842_),
    .X(_06032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09574_ (.A(_05931_),
    .B(_06032_),
    .X(_06033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09575_ (.A(_06033_),
    .X(_06034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09576_ (.A(_06034_),
    .X(_06035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09577_ (.A(_06033_),
    .Y(_06036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09578_ (.A(_06036_),
    .X(_06037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09579_ (.A(_06037_),
    .X(_06038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09580_ (.A1(\design_top.core0.REG1[7][31] ),
    .A2(_06035_),
    .B1(_05954_),
    .B2(_06038_),
    .X(_03435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09581_ (.A1(\design_top.core0.REG1[7][30] ),
    .A2(_06035_),
    .B1(_05975_),
    .B2(_06038_),
    .X(_03434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09582_ (.A1(\design_top.core0.REG1[7][29] ),
    .A2(_06035_),
    .B1(_05976_),
    .B2(_06038_),
    .X(_03433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09583_ (.A1(\design_top.core0.REG1[7][28] ),
    .A2(_06035_),
    .B1(_05977_),
    .B2(_06038_),
    .X(_03432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09584_ (.A(_06034_),
    .X(_06039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09585_ (.A1(\design_top.core0.REG1[7][27] ),
    .A2(_06039_),
    .B1(_05979_),
    .B2(_06038_),
    .X(_03431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09586_ (.A(_06037_),
    .X(_06040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09587_ (.A1(\design_top.core0.REG1[7][26] ),
    .A2(_06039_),
    .B1(_05980_),
    .B2(_06040_),
    .X(_03430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09588_ (.A1(\design_top.core0.REG1[7][25] ),
    .A2(_06039_),
    .B1(_05982_),
    .B2(_06040_),
    .X(_03429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09589_ (.A1(\design_top.core0.REG1[7][24] ),
    .A2(_06039_),
    .B1(_05983_),
    .B2(_06040_),
    .X(_03428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09590_ (.A1(\design_top.core0.REG1[7][23] ),
    .A2(_06039_),
    .B1(_05984_),
    .B2(_06040_),
    .X(_03427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09591_ (.A(_06034_),
    .X(_06041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09592_ (.A1(\design_top.core0.REG1[7][22] ),
    .A2(_06041_),
    .B1(_05986_),
    .B2(_06040_),
    .X(_03426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09593_ (.A(_06037_),
    .X(_06042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09594_ (.A1(\design_top.core0.REG1[7][21] ),
    .A2(_06041_),
    .B1(_05987_),
    .B2(_06042_),
    .X(_03425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09595_ (.A1(\design_top.core0.REG1[7][20] ),
    .A2(_06041_),
    .B1(_05989_),
    .B2(_06042_),
    .X(_03424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09596_ (.A1(\design_top.core0.REG1[7][19] ),
    .A2(_06041_),
    .B1(_05990_),
    .B2(_06042_),
    .X(_03423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09597_ (.A1(\design_top.core0.REG1[7][18] ),
    .A2(_06041_),
    .B1(_05991_),
    .B2(_06042_),
    .X(_03422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09598_ (.A(_06033_),
    .X(_06043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09599_ (.A1(\design_top.core0.REG1[7][17] ),
    .A2(_06043_),
    .B1(_05993_),
    .B2(_06042_),
    .X(_03421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09600_ (.A(_06036_),
    .X(_06044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09601_ (.A1(\design_top.core0.REG1[7][16] ),
    .A2(_06043_),
    .B1(_05994_),
    .B2(_06044_),
    .X(_03420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09602_ (.A1(\design_top.core0.REG1[7][15] ),
    .A2(_06043_),
    .B1(_05996_),
    .B2(_06044_),
    .X(_03419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09603_ (.A1(\design_top.core0.REG1[7][14] ),
    .A2(_06043_),
    .B1(_05997_),
    .B2(_06044_),
    .X(_03418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09604_ (.A1(\design_top.core0.REG1[7][13] ),
    .A2(_06037_),
    .B1(_05945_),
    .B2(_06035_),
    .X(_03417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09605_ (.A1(\design_top.core0.REG1[7][12] ),
    .A2(_06043_),
    .B1(_05998_),
    .B2(_06044_),
    .X(_03416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09606_ (.A(_06033_),
    .X(_06045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09607_ (.A1(\design_top.core0.REG1[7][11] ),
    .A2(_06045_),
    .B1(_06000_),
    .B2(_06044_),
    .X(_03415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09608_ (.A(_06036_),
    .X(_06046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09609_ (.A1(\design_top.core0.REG1[7][10] ),
    .A2(_06045_),
    .B1(_06001_),
    .B2(_06046_),
    .X(_03414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09610_ (.A1(\design_top.core0.REG1[7][9] ),
    .A2(_06045_),
    .B1(_06003_),
    .B2(_06046_),
    .X(_03413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09611_ (.A1(\design_top.core0.REG1[7][8] ),
    .A2(_06045_),
    .B1(_06004_),
    .B2(_06046_),
    .X(_03412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09612_ (.A1(\design_top.core0.REG1[7][7] ),
    .A2(_06045_),
    .B1(_06005_),
    .B2(_06046_),
    .X(_03411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09613_ (.A(_06033_),
    .X(_06047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09614_ (.A1(\design_top.core0.REG1[7][6] ),
    .A2(_06047_),
    .B1(_06007_),
    .B2(_06046_),
    .X(_03410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09615_ (.A(_06036_),
    .X(_06048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09616_ (.A1(\design_top.core0.REG1[7][5] ),
    .A2(_06047_),
    .B1(_06008_),
    .B2(_06048_),
    .X(_03409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09617_ (.A1(\design_top.core0.REG1[7][4] ),
    .A2(_06047_),
    .B1(_06010_),
    .B2(_06048_),
    .X(_03408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09618_ (.A1(\design_top.core0.REG1[7][3] ),
    .A2(_06047_),
    .B1(_06011_),
    .B2(_06048_),
    .X(_03407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09619_ (.A1(\design_top.core0.REG1[7][2] ),
    .A2(_06047_),
    .B1(_06012_),
    .B2(_06048_),
    .X(_03406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09620_ (.A1(\design_top.core0.REG1[7][1] ),
    .A2(_06034_),
    .B1(_06013_),
    .B2(_06048_),
    .X(_03405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09621_ (.A1(\design_top.core0.REG1[7][0] ),
    .A2(_06034_),
    .B1(_06014_),
    .B2(_06037_),
    .X(_03404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09622_ (.A(_05689_),
    .X(_06049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _09623_ (.A(_05168_),
    .B(_06049_),
    .Y(_00558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09624_ (.A(_05171_),
    .B(_00558_),
    .X(_06050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09625_ (.A(_06050_),
    .X(_06051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09626_ (.A(_06050_),
    .Y(_06052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09627_ (.A(_06052_),
    .X(_06053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09628_ (.A1(_00260_),
    .A2(_06051_),
    .B1(\design_top.MEM[4][7] ),
    .B2(_06053_),
    .X(_03403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09629_ (.A1(_00259_),
    .A2(_06051_),
    .B1(\design_top.MEM[4][6] ),
    .B2(_06053_),
    .X(_03402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09630_ (.A1(_00258_),
    .A2(_06051_),
    .B1(\design_top.MEM[4][5] ),
    .B2(_06053_),
    .X(_03401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09631_ (.A1(_00257_),
    .A2(_06051_),
    .B1(\design_top.MEM[4][4] ),
    .B2(_06053_),
    .X(_03400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09632_ (.A1(_00256_),
    .A2(_06051_),
    .B1(\design_top.MEM[4][3] ),
    .B2(_06053_),
    .X(_03399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09633_ (.A1(_00255_),
    .A2(_06050_),
    .B1(\design_top.MEM[4][2] ),
    .B2(_06052_),
    .X(_03398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09634_ (.A1(_00254_),
    .A2(_06050_),
    .B1(\design_top.MEM[4][1] ),
    .B2(_06052_),
    .X(_03397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09635_ (.A1(_00253_),
    .A2(_06050_),
    .B1(\design_top.MEM[4][0] ),
    .B2(_06052_),
    .X(_03396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09636_ (.A(_05745_),
    .X(_06054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _09637_ (.A(_05841_),
    .B(_05912_),
    .C(_01440_),
    .D(_05913_),
    .X(_06055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09638_ (.A(_06054_),
    .B(_06055_),
    .X(_06056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09639_ (.A(_06056_),
    .X(_06057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09640_ (.A(_06057_),
    .X(_06058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09641_ (.A(_06056_),
    .Y(_06059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09642_ (.A(_06059_),
    .X(_06060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09643_ (.A(_06060_),
    .X(_06061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09644_ (.A1(\design_top.core0.REG1[8][31] ),
    .A2(_06058_),
    .B1(_05954_),
    .B2(_06061_),
    .X(_03395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09645_ (.A1(\design_top.core0.REG1[8][30] ),
    .A2(_06058_),
    .B1(_05975_),
    .B2(_06061_),
    .X(_03394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09646_ (.A1(\design_top.core0.REG1[8][29] ),
    .A2(_06058_),
    .B1(_05976_),
    .B2(_06061_),
    .X(_03393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09647_ (.A1(\design_top.core0.REG1[8][28] ),
    .A2(_06058_),
    .B1(_05977_),
    .B2(_06061_),
    .X(_03392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09648_ (.A(_06057_),
    .X(_06062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09649_ (.A1(\design_top.core0.REG1[8][27] ),
    .A2(_06062_),
    .B1(_05979_),
    .B2(_06061_),
    .X(_03391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09650_ (.A(_06060_),
    .X(_06063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09651_ (.A1(\design_top.core0.REG1[8][26] ),
    .A2(_06062_),
    .B1(_05980_),
    .B2(_06063_),
    .X(_03390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09652_ (.A1(\design_top.core0.REG1[8][25] ),
    .A2(_06062_),
    .B1(_05982_),
    .B2(_06063_),
    .X(_03389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09653_ (.A1(\design_top.core0.REG1[8][24] ),
    .A2(_06062_),
    .B1(_05983_),
    .B2(_06063_),
    .X(_03388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09654_ (.A1(\design_top.core0.REG1[8][23] ),
    .A2(_06062_),
    .B1(_05984_),
    .B2(_06063_),
    .X(_03387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09655_ (.A(_06057_),
    .X(_06064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09656_ (.A1(\design_top.core0.REG1[8][22] ),
    .A2(_06064_),
    .B1(_05986_),
    .B2(_06063_),
    .X(_03386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09657_ (.A(_06060_),
    .X(_06065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09658_ (.A1(\design_top.core0.REG1[8][21] ),
    .A2(_06064_),
    .B1(_05987_),
    .B2(_06065_),
    .X(_03385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09659_ (.A1(\design_top.core0.REG1[8][20] ),
    .A2(_06064_),
    .B1(_05989_),
    .B2(_06065_),
    .X(_03384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09660_ (.A1(\design_top.core0.REG1[8][19] ),
    .A2(_06064_),
    .B1(_05990_),
    .B2(_06065_),
    .X(_03383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09661_ (.A1(\design_top.core0.REG1[8][18] ),
    .A2(_06064_),
    .B1(_05991_),
    .B2(_06065_),
    .X(_03382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09662_ (.A(_06056_),
    .X(_06066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09663_ (.A1(\design_top.core0.REG1[8][17] ),
    .A2(_06066_),
    .B1(_05993_),
    .B2(_06065_),
    .X(_03381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09664_ (.A(_06059_),
    .X(_06067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09665_ (.A1(\design_top.core0.REG1[8][16] ),
    .A2(_06066_),
    .B1(_05994_),
    .B2(_06067_),
    .X(_03380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09666_ (.A1(\design_top.core0.REG1[8][15] ),
    .A2(_06066_),
    .B1(_05996_),
    .B2(_06067_),
    .X(_03379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09667_ (.A1(\design_top.core0.REG1[8][14] ),
    .A2(_06066_),
    .B1(_05997_),
    .B2(_06067_),
    .X(_03378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09668_ (.A(_00045_),
    .X(_06068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09669_ (.A1(\design_top.core0.REG1[8][13] ),
    .A2(_06060_),
    .B1(_06068_),
    .B2(_06058_),
    .X(_03377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09670_ (.A1(\design_top.core0.REG1[8][12] ),
    .A2(_06066_),
    .B1(_05998_),
    .B2(_06067_),
    .X(_03376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09671_ (.A(_06056_),
    .X(_06069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09672_ (.A1(\design_top.core0.REG1[8][11] ),
    .A2(_06069_),
    .B1(_06000_),
    .B2(_06067_),
    .X(_03375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09673_ (.A(_06059_),
    .X(_06070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09674_ (.A1(\design_top.core0.REG1[8][10] ),
    .A2(_06069_),
    .B1(_06001_),
    .B2(_06070_),
    .X(_03374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09675_ (.A1(\design_top.core0.REG1[8][9] ),
    .A2(_06069_),
    .B1(_06003_),
    .B2(_06070_),
    .X(_03373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09676_ (.A1(\design_top.core0.REG1[8][8] ),
    .A2(_06069_),
    .B1(_06004_),
    .B2(_06070_),
    .X(_03372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09677_ (.A1(\design_top.core0.REG1[8][7] ),
    .A2(_06069_),
    .B1(_06005_),
    .B2(_06070_),
    .X(_03371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09678_ (.A(_06056_),
    .X(_06071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09679_ (.A1(\design_top.core0.REG1[8][6] ),
    .A2(_06071_),
    .B1(_06007_),
    .B2(_06070_),
    .X(_03370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09680_ (.A(_06059_),
    .X(_06072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09681_ (.A1(\design_top.core0.REG1[8][5] ),
    .A2(_06071_),
    .B1(_06008_),
    .B2(_06072_),
    .X(_03369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09682_ (.A1(\design_top.core0.REG1[8][4] ),
    .A2(_06071_),
    .B1(_06010_),
    .B2(_06072_),
    .X(_03368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09683_ (.A1(\design_top.core0.REG1[8][3] ),
    .A2(_06071_),
    .B1(_06011_),
    .B2(_06072_),
    .X(_03367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09684_ (.A1(\design_top.core0.REG1[8][2] ),
    .A2(_06071_),
    .B1(_06012_),
    .B2(_06072_),
    .X(_03366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09685_ (.A1(\design_top.core0.REG1[8][1] ),
    .A2(_06057_),
    .B1(_06013_),
    .B2(_06072_),
    .X(_03365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09686_ (.A1(\design_top.core0.REG1[8][0] ),
    .A2(_06057_),
    .B1(_06014_),
    .B2(_06060_),
    .X(_03364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09687_ (.A(\design_top.core0.REG1[0][31] ),
    .Y(_00361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09688_ (.A(_05603_),
    .X(_06073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09689_ (.A(_06073_),
    .B(_05746_),
    .X(_06074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09690_ (.A(_06074_),
    .Y(_06075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _09691_ (.A(_00361_),
    .B(_06075_),
    .Y(_03363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09692_ (.A(_06074_),
    .X(_06076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09693_ (.A(_06076_),
    .X(_06077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09694_ (.A(\design_top.core0.REG1[0][30] ),
    .B(_06077_),
    .X(_03362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09695_ (.A(\design_top.core0.REG1[0][29] ),
    .B(_06077_),
    .X(_03361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09696_ (.A(\design_top.core0.REG1[0][28] ),
    .B(_06077_),
    .X(_03360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09697_ (.A(\design_top.core0.REG1[0][27] ),
    .B(_06077_),
    .X(_03359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09698_ (.A(_06076_),
    .X(_06078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09699_ (.A(\design_top.core0.REG1[0][26] ),
    .B(_06078_),
    .X(_03358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09700_ (.A(\design_top.core0.REG1[0][25] ),
    .B(_06078_),
    .X(_03357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09701_ (.A(\design_top.core0.REG1[0][24] ),
    .B(_06078_),
    .X(_03356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09702_ (.A(\design_top.core0.REG1[0][23] ),
    .B(_06078_),
    .X(_03355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09703_ (.A(\design_top.core0.REG1[0][22] ),
    .B(_06078_),
    .X(_03354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09704_ (.A(_06076_),
    .X(_06079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09705_ (.A(\design_top.core0.REG1[0][21] ),
    .B(_06079_),
    .X(_03353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09706_ (.A(\design_top.core0.REG1[0][20] ),
    .B(_06079_),
    .X(_03352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09707_ (.A(\design_top.core0.REG1[0][19] ),
    .B(_06079_),
    .X(_03351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09708_ (.A(\design_top.core0.REG1[0][18] ),
    .B(_06079_),
    .X(_03350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09709_ (.A(\design_top.core0.REG1[0][17] ),
    .B(_06079_),
    .X(_03349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09710_ (.A(_06076_),
    .X(_06080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09711_ (.A(\design_top.core0.REG1[0][16] ),
    .B(_06080_),
    .X(_03348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09712_ (.A(\design_top.core0.REG1[0][15] ),
    .B(_06080_),
    .X(_03347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09713_ (.A(\design_top.core0.REG1[0][14] ),
    .B(_06080_),
    .X(_03346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09714_ (.A1(\design_top.core0.REG1[0][13] ),
    .A2(_06075_),
    .B1(_06068_),
    .B2(_06077_),
    .X(_03345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09715_ (.A(\design_top.core0.REG1[0][12] ),
    .B(_06080_),
    .X(_03344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09716_ (.A(\design_top.core0.REG1[0][11] ),
    .B(_06080_),
    .X(_03343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09717_ (.A(_06074_),
    .X(_06081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09718_ (.A(\design_top.core0.REG1[0][10] ),
    .B(_06081_),
    .X(_03342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09719_ (.A(\design_top.core0.REG1[0][9] ),
    .B(_06081_),
    .X(_03341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09720_ (.A(\design_top.core0.REG1[0][8] ),
    .B(_06081_),
    .X(_03340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09721_ (.A(\design_top.core0.REG1[0][7] ),
    .B(_06081_),
    .X(_03339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09722_ (.A(\design_top.core0.REG1[0][6] ),
    .B(_06081_),
    .X(_03338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09723_ (.A(_06074_),
    .X(_06082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09724_ (.A(\design_top.core0.REG1[0][5] ),
    .B(_06082_),
    .X(_03337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09725_ (.A(\design_top.core0.REG1[0][4] ),
    .B(_06082_),
    .X(_03336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09726_ (.A(\design_top.core0.REG1[0][3] ),
    .B(_06082_),
    .X(_03335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09727_ (.A(\design_top.core0.REG1[0][2] ),
    .B(_06082_),
    .X(_03334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09728_ (.A(\design_top.core0.REG1[0][1] ),
    .B(_06082_),
    .X(_03333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _09729_ (.A(\design_top.core0.REG1[0][0] ),
    .B(_06076_),
    .X(_03332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _09730_ (.A(_05841_),
    .B(_05912_),
    .C(_05844_),
    .D(_01439_),
    .X(_06083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09731_ (.A(_06054_),
    .B(_06083_),
    .X(_06084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09732_ (.A(_06084_),
    .X(_06085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09733_ (.A(_06085_),
    .X(_06086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09734_ (.A(_05749_),
    .X(_06087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09735_ (.A(_06084_),
    .Y(_06088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09736_ (.A(_06088_),
    .X(_06089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09737_ (.A(_06089_),
    .X(_06090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09738_ (.A1(\design_top.core0.REG1[10][31] ),
    .A2(_06086_),
    .B1(_06087_),
    .B2(_06090_),
    .X(_03331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09739_ (.A1(\design_top.core0.REG1[10][30] ),
    .A2(_06086_),
    .B1(_05975_),
    .B2(_06090_),
    .X(_03330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09740_ (.A1(\design_top.core0.REG1[10][29] ),
    .A2(_06086_),
    .B1(_05976_),
    .B2(_06090_),
    .X(_03329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09741_ (.A1(\design_top.core0.REG1[10][28] ),
    .A2(_06086_),
    .B1(_05977_),
    .B2(_06090_),
    .X(_03328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09742_ (.A(_06085_),
    .X(_06091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09743_ (.A1(\design_top.core0.REG1[10][27] ),
    .A2(_06091_),
    .B1(_05979_),
    .B2(_06090_),
    .X(_03327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09744_ (.A(_06089_),
    .X(_06092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09745_ (.A1(\design_top.core0.REG1[10][26] ),
    .A2(_06091_),
    .B1(_05980_),
    .B2(_06092_),
    .X(_03326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09746_ (.A1(\design_top.core0.REG1[10][25] ),
    .A2(_06091_),
    .B1(_05982_),
    .B2(_06092_),
    .X(_03325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09747_ (.A1(\design_top.core0.REG1[10][24] ),
    .A2(_06091_),
    .B1(_05983_),
    .B2(_06092_),
    .X(_03324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09748_ (.A1(\design_top.core0.REG1[10][23] ),
    .A2(_06091_),
    .B1(_05984_),
    .B2(_06092_),
    .X(_03323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09749_ (.A(_06085_),
    .X(_06093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09750_ (.A1(\design_top.core0.REG1[10][22] ),
    .A2(_06093_),
    .B1(_05986_),
    .B2(_06092_),
    .X(_03322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09751_ (.A(_06089_),
    .X(_06094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09752_ (.A1(\design_top.core0.REG1[10][21] ),
    .A2(_06093_),
    .B1(_05987_),
    .B2(_06094_),
    .X(_03321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09753_ (.A1(\design_top.core0.REG1[10][20] ),
    .A2(_06093_),
    .B1(_05989_),
    .B2(_06094_),
    .X(_03320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09754_ (.A1(\design_top.core0.REG1[10][19] ),
    .A2(_06093_),
    .B1(_05990_),
    .B2(_06094_),
    .X(_03319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09755_ (.A1(\design_top.core0.REG1[10][18] ),
    .A2(_06093_),
    .B1(_05991_),
    .B2(_06094_),
    .X(_03318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09756_ (.A(_06084_),
    .X(_06095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09757_ (.A1(\design_top.core0.REG1[10][17] ),
    .A2(_06095_),
    .B1(_05993_),
    .B2(_06094_),
    .X(_03317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09758_ (.A(_06088_),
    .X(_06096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09759_ (.A1(\design_top.core0.REG1[10][16] ),
    .A2(_06095_),
    .B1(_05994_),
    .B2(_06096_),
    .X(_03316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09760_ (.A1(\design_top.core0.REG1[10][15] ),
    .A2(_06095_),
    .B1(_05996_),
    .B2(_06096_),
    .X(_03315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09761_ (.A1(\design_top.core0.REG1[10][14] ),
    .A2(_06095_),
    .B1(_05997_),
    .B2(_06096_),
    .X(_03314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09762_ (.A1(\design_top.core0.REG1[10][13] ),
    .A2(_06089_),
    .B1(_06068_),
    .B2(_06086_),
    .X(_03313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09763_ (.A1(\design_top.core0.REG1[10][12] ),
    .A2(_06095_),
    .B1(_05998_),
    .B2(_06096_),
    .X(_03312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09764_ (.A(_06084_),
    .X(_06097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09765_ (.A1(\design_top.core0.REG1[10][11] ),
    .A2(_06097_),
    .B1(_06000_),
    .B2(_06096_),
    .X(_03311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09766_ (.A(_06088_),
    .X(_06098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09767_ (.A1(\design_top.core0.REG1[10][10] ),
    .A2(_06097_),
    .B1(_06001_),
    .B2(_06098_),
    .X(_03310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09768_ (.A1(\design_top.core0.REG1[10][9] ),
    .A2(_06097_),
    .B1(_06003_),
    .B2(_06098_),
    .X(_03309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09769_ (.A1(\design_top.core0.REG1[10][8] ),
    .A2(_06097_),
    .B1(_06004_),
    .B2(_06098_),
    .X(_03308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09770_ (.A1(\design_top.core0.REG1[10][7] ),
    .A2(_06097_),
    .B1(_06005_),
    .B2(_06098_),
    .X(_03307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09771_ (.A(_06084_),
    .X(_06099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09772_ (.A1(\design_top.core0.REG1[10][6] ),
    .A2(_06099_),
    .B1(_06007_),
    .B2(_06098_),
    .X(_03306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09773_ (.A(_06088_),
    .X(_06100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09774_ (.A1(\design_top.core0.REG1[10][5] ),
    .A2(_06099_),
    .B1(_06008_),
    .B2(_06100_),
    .X(_03305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09775_ (.A1(\design_top.core0.REG1[10][4] ),
    .A2(_06099_),
    .B1(_06010_),
    .B2(_06100_),
    .X(_03304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09776_ (.A1(\design_top.core0.REG1[10][3] ),
    .A2(_06099_),
    .B1(_06011_),
    .B2(_06100_),
    .X(_03303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09777_ (.A1(\design_top.core0.REG1[10][2] ),
    .A2(_06099_),
    .B1(_06012_),
    .B2(_06100_),
    .X(_03302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09778_ (.A1(\design_top.core0.REG1[10][1] ),
    .A2(_06085_),
    .B1(_06013_),
    .B2(_06100_),
    .X(_03301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09779_ (.A1(\design_top.core0.REG1[10][0] ),
    .A2(_06085_),
    .B1(_06014_),
    .B2(_06089_),
    .X(_03300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _09780_ (.A(_05841_),
    .B(_05912_),
    .C(_05844_),
    .D(_05595_),
    .X(_06101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09781_ (.A(_06054_),
    .B(_06101_),
    .X(_06102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09782_ (.A(_06102_),
    .X(_06103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09783_ (.A(_06103_),
    .X(_06104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09784_ (.A(_06102_),
    .Y(_06105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09785_ (.A(_06105_),
    .X(_06106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09786_ (.A(_06106_),
    .X(_06107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09787_ (.A1(\design_top.core0.REG1[11][31] ),
    .A2(_06104_),
    .B1(_06087_),
    .B2(_06107_),
    .X(_03299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09788_ (.A1(\design_top.core0.REG1[11][30] ),
    .A2(_06104_),
    .B1(_05754_),
    .B2(_06107_),
    .X(_03298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09789_ (.A1(\design_top.core0.REG1[11][29] ),
    .A2(_06104_),
    .B1(_05758_),
    .B2(_06107_),
    .X(_03297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09790_ (.A1(\design_top.core0.REG1[11][28] ),
    .A2(_06104_),
    .B1(_05760_),
    .B2(_06107_),
    .X(_03296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09791_ (.A(_06103_),
    .X(_06108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09792_ (.A1(\design_top.core0.REG1[11][27] ),
    .A2(_06108_),
    .B1(_05762_),
    .B2(_06107_),
    .X(_03295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09793_ (.A(_06106_),
    .X(_06109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09794_ (.A1(\design_top.core0.REG1[11][26] ),
    .A2(_06108_),
    .B1(_05764_),
    .B2(_06109_),
    .X(_03294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09795_ (.A1(\design_top.core0.REG1[11][25] ),
    .A2(_06108_),
    .B1(_05766_),
    .B2(_06109_),
    .X(_03293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09796_ (.A1(\design_top.core0.REG1[11][24] ),
    .A2(_06108_),
    .B1(_05770_),
    .B2(_06109_),
    .X(_03292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09797_ (.A1(\design_top.core0.REG1[11][23] ),
    .A2(_06108_),
    .B1(_05772_),
    .B2(_06109_),
    .X(_03291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09798_ (.A(_06103_),
    .X(_06110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09799_ (.A1(\design_top.core0.REG1[11][22] ),
    .A2(_06110_),
    .B1(_05774_),
    .B2(_06109_),
    .X(_03290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09800_ (.A(_06106_),
    .X(_06111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09801_ (.A1(\design_top.core0.REG1[11][21] ),
    .A2(_06110_),
    .B1(_05776_),
    .B2(_06111_),
    .X(_03289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09802_ (.A1(\design_top.core0.REG1[11][20] ),
    .A2(_06110_),
    .B1(_05778_),
    .B2(_06111_),
    .X(_03288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09803_ (.A1(\design_top.core0.REG1[11][19] ),
    .A2(_06110_),
    .B1(_05782_),
    .B2(_06111_),
    .X(_03287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09804_ (.A1(\design_top.core0.REG1[11][18] ),
    .A2(_06110_),
    .B1(_05784_),
    .B2(_06111_),
    .X(_03286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09805_ (.A(_06102_),
    .X(_06112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09806_ (.A1(\design_top.core0.REG1[11][17] ),
    .A2(_06112_),
    .B1(_05786_),
    .B2(_06111_),
    .X(_03285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09807_ (.A(_06105_),
    .X(_06113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09808_ (.A1(\design_top.core0.REG1[11][16] ),
    .A2(_06112_),
    .B1(_05788_),
    .B2(_06113_),
    .X(_03284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09809_ (.A1(\design_top.core0.REG1[11][15] ),
    .A2(_06112_),
    .B1(_05790_),
    .B2(_06113_),
    .X(_03283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09810_ (.A1(\design_top.core0.REG1[11][14] ),
    .A2(_06112_),
    .B1(_05794_),
    .B2(_06113_),
    .X(_03282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09811_ (.A1(\design_top.core0.REG1[11][13] ),
    .A2(_06106_),
    .B1(_06068_),
    .B2(_06104_),
    .X(_03281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09812_ (.A1(\design_top.core0.REG1[11][12] ),
    .A2(_06112_),
    .B1(_05796_),
    .B2(_06113_),
    .X(_03280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09813_ (.A(_06102_),
    .X(_06114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09814_ (.A1(\design_top.core0.REG1[11][11] ),
    .A2(_06114_),
    .B1(_05798_),
    .B2(_06113_),
    .X(_03279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09815_ (.A(_06105_),
    .X(_06115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09816_ (.A1(\design_top.core0.REG1[11][10] ),
    .A2(_06114_),
    .B1(_05800_),
    .B2(_06115_),
    .X(_03278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09817_ (.A1(\design_top.core0.REG1[11][9] ),
    .A2(_06114_),
    .B1(_05802_),
    .B2(_06115_),
    .X(_03277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09818_ (.A1(\design_top.core0.REG1[11][8] ),
    .A2(_06114_),
    .B1(_05806_),
    .B2(_06115_),
    .X(_03276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09819_ (.A1(\design_top.core0.REG1[11][7] ),
    .A2(_06114_),
    .B1(_05808_),
    .B2(_06115_),
    .X(_03275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09820_ (.A(_06102_),
    .X(_06116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09821_ (.A1(\design_top.core0.REG1[11][6] ),
    .A2(_06116_),
    .B1(_05810_),
    .B2(_06115_),
    .X(_03274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09822_ (.A(_06105_),
    .X(_06117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09823_ (.A1(\design_top.core0.REG1[11][5] ),
    .A2(_06116_),
    .B1(_05812_),
    .B2(_06117_),
    .X(_03273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09824_ (.A1(\design_top.core0.REG1[11][4] ),
    .A2(_06116_),
    .B1(_05814_),
    .B2(_06117_),
    .X(_03272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09825_ (.A1(\design_top.core0.REG1[11][3] ),
    .A2(_06116_),
    .B1(_05818_),
    .B2(_06117_),
    .X(_03271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09826_ (.A1(\design_top.core0.REG1[11][2] ),
    .A2(_06116_),
    .B1(_05820_),
    .B2(_06117_),
    .X(_03270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09827_ (.A1(\design_top.core0.REG1[11][1] ),
    .A2(_06103_),
    .B1(_05822_),
    .B2(_06117_),
    .X(_03269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09828_ (.A1(\design_top.core0.REG1[11][0] ),
    .A2(_06103_),
    .B1(_05824_),
    .B2(_06106_),
    .X(_03268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _09829_ (.A(_05594_),
    .B(_05913_),
    .C(_05597_),
    .D(_05842_),
    .X(_06118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09830_ (.A(_06054_),
    .B(_06118_),
    .X(_06119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09831_ (.A(_06119_),
    .X(_06120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09832_ (.A(_06120_),
    .X(_06121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09833_ (.A(_06119_),
    .Y(_06122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09834_ (.A(_06122_),
    .X(_06123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09835_ (.A(_06123_),
    .X(_06124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09836_ (.A1(\design_top.core0.REG1[12][31] ),
    .A2(_06121_),
    .B1(_06087_),
    .B2(_06124_),
    .X(_03267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09837_ (.A1(\design_top.core0.REG1[12][30] ),
    .A2(_06121_),
    .B1(_05754_),
    .B2(_06124_),
    .X(_03266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09838_ (.A1(\design_top.core0.REG1[12][29] ),
    .A2(_06121_),
    .B1(_05758_),
    .B2(_06124_),
    .X(_03265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09839_ (.A1(\design_top.core0.REG1[12][28] ),
    .A2(_06121_),
    .B1(_05760_),
    .B2(_06124_),
    .X(_03264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09840_ (.A(_06120_),
    .X(_06125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09841_ (.A1(\design_top.core0.REG1[12][27] ),
    .A2(_06125_),
    .B1(_05762_),
    .B2(_06124_),
    .X(_03263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09842_ (.A(_06123_),
    .X(_06126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09843_ (.A1(\design_top.core0.REG1[12][26] ),
    .A2(_06125_),
    .B1(_05764_),
    .B2(_06126_),
    .X(_03262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09844_ (.A1(\design_top.core0.REG1[12][25] ),
    .A2(_06125_),
    .B1(_05766_),
    .B2(_06126_),
    .X(_03261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09845_ (.A1(\design_top.core0.REG1[12][24] ),
    .A2(_06125_),
    .B1(_05770_),
    .B2(_06126_),
    .X(_03260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09846_ (.A1(\design_top.core0.REG1[12][23] ),
    .A2(_06125_),
    .B1(_05772_),
    .B2(_06126_),
    .X(_03259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09847_ (.A(_06120_),
    .X(_06127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09848_ (.A1(\design_top.core0.REG1[12][22] ),
    .A2(_06127_),
    .B1(_05774_),
    .B2(_06126_),
    .X(_03258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09849_ (.A(_06123_),
    .X(_06128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09850_ (.A1(\design_top.core0.REG1[12][21] ),
    .A2(_06127_),
    .B1(_05776_),
    .B2(_06128_),
    .X(_03257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09851_ (.A1(\design_top.core0.REG1[12][20] ),
    .A2(_06127_),
    .B1(_05778_),
    .B2(_06128_),
    .X(_03256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09852_ (.A1(\design_top.core0.REG1[12][19] ),
    .A2(_06127_),
    .B1(_05782_),
    .B2(_06128_),
    .X(_03255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09853_ (.A1(\design_top.core0.REG1[12][18] ),
    .A2(_06127_),
    .B1(_05784_),
    .B2(_06128_),
    .X(_03254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09854_ (.A(_06119_),
    .X(_06129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09855_ (.A1(\design_top.core0.REG1[12][17] ),
    .A2(_06129_),
    .B1(_05786_),
    .B2(_06128_),
    .X(_03253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09856_ (.A(_06122_),
    .X(_06130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09857_ (.A1(\design_top.core0.REG1[12][16] ),
    .A2(_06129_),
    .B1(_05788_),
    .B2(_06130_),
    .X(_03252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09858_ (.A1(\design_top.core0.REG1[12][15] ),
    .A2(_06129_),
    .B1(_05790_),
    .B2(_06130_),
    .X(_03251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09859_ (.A1(\design_top.core0.REG1[12][14] ),
    .A2(_06129_),
    .B1(_05794_),
    .B2(_06130_),
    .X(_03250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09860_ (.A1(\design_top.core0.REG1[12][13] ),
    .A2(_06123_),
    .B1(_06068_),
    .B2(_06121_),
    .X(_03249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09861_ (.A1(\design_top.core0.REG1[12][12] ),
    .A2(_06129_),
    .B1(_05796_),
    .B2(_06130_),
    .X(_03248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09862_ (.A(_06119_),
    .X(_06131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09863_ (.A1(\design_top.core0.REG1[12][11] ),
    .A2(_06131_),
    .B1(_05798_),
    .B2(_06130_),
    .X(_03247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09864_ (.A(_06122_),
    .X(_06132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09865_ (.A1(\design_top.core0.REG1[12][10] ),
    .A2(_06131_),
    .B1(_05800_),
    .B2(_06132_),
    .X(_03246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09866_ (.A1(\design_top.core0.REG1[12][9] ),
    .A2(_06131_),
    .B1(_05802_),
    .B2(_06132_),
    .X(_03245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09867_ (.A1(\design_top.core0.REG1[12][8] ),
    .A2(_06131_),
    .B1(_05806_),
    .B2(_06132_),
    .X(_03244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09868_ (.A1(\design_top.core0.REG1[12][7] ),
    .A2(_06131_),
    .B1(_05808_),
    .B2(_06132_),
    .X(_03243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09869_ (.A(_06119_),
    .X(_06133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09870_ (.A1(\design_top.core0.REG1[12][6] ),
    .A2(_06133_),
    .B1(_05810_),
    .B2(_06132_),
    .X(_03242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09871_ (.A(_06122_),
    .X(_06134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09872_ (.A1(\design_top.core0.REG1[12][5] ),
    .A2(_06133_),
    .B1(_05812_),
    .B2(_06134_),
    .X(_03241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09873_ (.A1(\design_top.core0.REG1[12][4] ),
    .A2(_06133_),
    .B1(_05814_),
    .B2(_06134_),
    .X(_03240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09874_ (.A1(\design_top.core0.REG1[12][3] ),
    .A2(_06133_),
    .B1(_05818_),
    .B2(_06134_),
    .X(_03239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09875_ (.A1(\design_top.core0.REG1[12][2] ),
    .A2(_06133_),
    .B1(_05820_),
    .B2(_06134_),
    .X(_03238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09876_ (.A1(\design_top.core0.REG1[12][1] ),
    .A2(_06120_),
    .B1(_05822_),
    .B2(_06134_),
    .X(_03237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09877_ (.A1(\design_top.core0.REG1[12][0] ),
    .A2(_06120_),
    .B1(_05824_),
    .B2(_06123_),
    .X(_03236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _09878_ (.A(_01440_),
    .B(_05596_),
    .C(_05597_),
    .D(_05842_),
    .X(_06135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09879_ (.A(_06054_),
    .B(_06135_),
    .X(_06136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09880_ (.A(_06136_),
    .X(_06137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09881_ (.A(_06137_),
    .X(_06138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09882_ (.A(_06136_),
    .Y(_06139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09883_ (.A(_06139_),
    .X(_06140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09884_ (.A(_06140_),
    .X(_06141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09885_ (.A1(\design_top.core0.REG1[13][31] ),
    .A2(_06138_),
    .B1(_06087_),
    .B2(_06141_),
    .X(_03235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09886_ (.A1(\design_top.core0.REG1[13][30] ),
    .A2(_06138_),
    .B1(_05754_),
    .B2(_06141_),
    .X(_03234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09887_ (.A1(\design_top.core0.REG1[13][29] ),
    .A2(_06138_),
    .B1(_05758_),
    .B2(_06141_),
    .X(_03233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09888_ (.A1(\design_top.core0.REG1[13][28] ),
    .A2(_06138_),
    .B1(_05760_),
    .B2(_06141_),
    .X(_03232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09889_ (.A(_06137_),
    .X(_06142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09890_ (.A1(\design_top.core0.REG1[13][27] ),
    .A2(_06142_),
    .B1(_05762_),
    .B2(_06141_),
    .X(_03231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09891_ (.A(_06140_),
    .X(_06143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09892_ (.A1(\design_top.core0.REG1[13][26] ),
    .A2(_06142_),
    .B1(_05764_),
    .B2(_06143_),
    .X(_03230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09893_ (.A1(\design_top.core0.REG1[13][25] ),
    .A2(_06142_),
    .B1(_05766_),
    .B2(_06143_),
    .X(_03229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09894_ (.A1(\design_top.core0.REG1[13][24] ),
    .A2(_06142_),
    .B1(_05770_),
    .B2(_06143_),
    .X(_03228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09895_ (.A1(\design_top.core0.REG1[13][23] ),
    .A2(_06142_),
    .B1(_05772_),
    .B2(_06143_),
    .X(_03227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09896_ (.A(_06137_),
    .X(_06144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09897_ (.A1(\design_top.core0.REG1[13][22] ),
    .A2(_06144_),
    .B1(_05774_),
    .B2(_06143_),
    .X(_03226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09898_ (.A(_06140_),
    .X(_06145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09899_ (.A1(\design_top.core0.REG1[13][21] ),
    .A2(_06144_),
    .B1(_05776_),
    .B2(_06145_),
    .X(_03225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09900_ (.A1(\design_top.core0.REG1[13][20] ),
    .A2(_06144_),
    .B1(_05778_),
    .B2(_06145_),
    .X(_03224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09901_ (.A1(\design_top.core0.REG1[13][19] ),
    .A2(_06144_),
    .B1(_05782_),
    .B2(_06145_),
    .X(_03223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09902_ (.A1(\design_top.core0.REG1[13][18] ),
    .A2(_06144_),
    .B1(_05784_),
    .B2(_06145_),
    .X(_03222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09903_ (.A(_06136_),
    .X(_06146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09904_ (.A1(\design_top.core0.REG1[13][17] ),
    .A2(_06146_),
    .B1(_05786_),
    .B2(_06145_),
    .X(_03221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09905_ (.A(_06139_),
    .X(_06147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09906_ (.A1(\design_top.core0.REG1[13][16] ),
    .A2(_06146_),
    .B1(_05788_),
    .B2(_06147_),
    .X(_03220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09907_ (.A1(\design_top.core0.REG1[13][15] ),
    .A2(_06146_),
    .B1(_05790_),
    .B2(_06147_),
    .X(_03219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09908_ (.A1(\design_top.core0.REG1[13][14] ),
    .A2(_06146_),
    .B1(_05794_),
    .B2(_06147_),
    .X(_03218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09909_ (.A1(\design_top.core0.REG1[13][13] ),
    .A2(_06140_),
    .B1(_05655_),
    .B2(_06138_),
    .X(_03217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09910_ (.A1(\design_top.core0.REG1[13][12] ),
    .A2(_06146_),
    .B1(_05796_),
    .B2(_06147_),
    .X(_03216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09911_ (.A(_06136_),
    .X(_06148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09912_ (.A1(\design_top.core0.REG1[13][11] ),
    .A2(_06148_),
    .B1(_05798_),
    .B2(_06147_),
    .X(_03215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09913_ (.A(_06139_),
    .X(_06149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09914_ (.A1(\design_top.core0.REG1[13][10] ),
    .A2(_06148_),
    .B1(_05800_),
    .B2(_06149_),
    .X(_03214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09915_ (.A1(\design_top.core0.REG1[13][9] ),
    .A2(_06148_),
    .B1(_05802_),
    .B2(_06149_),
    .X(_03213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09916_ (.A1(\design_top.core0.REG1[13][8] ),
    .A2(_06148_),
    .B1(_05806_),
    .B2(_06149_),
    .X(_03212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09917_ (.A1(\design_top.core0.REG1[13][7] ),
    .A2(_06148_),
    .B1(_05808_),
    .B2(_06149_),
    .X(_03211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09918_ (.A(_06136_),
    .X(_06150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09919_ (.A1(\design_top.core0.REG1[13][6] ),
    .A2(_06150_),
    .B1(_05810_),
    .B2(_06149_),
    .X(_03210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09920_ (.A(_06139_),
    .X(_06151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09921_ (.A1(\design_top.core0.REG1[13][5] ),
    .A2(_06150_),
    .B1(_05812_),
    .B2(_06151_),
    .X(_03209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09922_ (.A1(\design_top.core0.REG1[13][4] ),
    .A2(_06150_),
    .B1(_05814_),
    .B2(_06151_),
    .X(_03208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09923_ (.A1(\design_top.core0.REG1[13][3] ),
    .A2(_06150_),
    .B1(_05818_),
    .B2(_06151_),
    .X(_03207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09924_ (.A1(\design_top.core0.REG1[13][2] ),
    .A2(_06150_),
    .B1(_05820_),
    .B2(_06151_),
    .X(_03206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09925_ (.A1(\design_top.core0.REG1[13][1] ),
    .A2(_06137_),
    .B1(_05822_),
    .B2(_06151_),
    .X(_03205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09926_ (.A1(\design_top.core0.REG1[13][0] ),
    .A2(_06137_),
    .B1(_05824_),
    .B2(_06140_),
    .X(_03204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _09927_ (.A(_05841_),
    .B(_05843_),
    .C(_05844_),
    .D(_01439_),
    .X(_06152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09928_ (.A(_05745_),
    .B(_06152_),
    .X(_06153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09929_ (.A(_06153_),
    .X(_06154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09930_ (.A(_06154_),
    .X(_06155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09931_ (.A(_06153_),
    .Y(_06156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09932_ (.A(_06156_),
    .X(_06157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09933_ (.A(_06157_),
    .X(_06158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09934_ (.A1(\design_top.core0.REG1[14][31] ),
    .A2(_06155_),
    .B1(_06087_),
    .B2(_06158_),
    .X(_03203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09935_ (.A1(\design_top.core0.REG1[14][30] ),
    .A2(_06155_),
    .B1(_05754_),
    .B2(_06158_),
    .X(_03202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09936_ (.A1(\design_top.core0.REG1[14][29] ),
    .A2(_06155_),
    .B1(_05758_),
    .B2(_06158_),
    .X(_03201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09937_ (.A1(\design_top.core0.REG1[14][28] ),
    .A2(_06155_),
    .B1(_05760_),
    .B2(_06158_),
    .X(_03200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09938_ (.A(_06154_),
    .X(_06159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09939_ (.A1(\design_top.core0.REG1[14][27] ),
    .A2(_06159_),
    .B1(_05762_),
    .B2(_06158_),
    .X(_03199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09940_ (.A(_06157_),
    .X(_06160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09941_ (.A1(\design_top.core0.REG1[14][26] ),
    .A2(_06159_),
    .B1(_05764_),
    .B2(_06160_),
    .X(_03198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09942_ (.A1(\design_top.core0.REG1[14][25] ),
    .A2(_06159_),
    .B1(_05766_),
    .B2(_06160_),
    .X(_03197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09943_ (.A1(\design_top.core0.REG1[14][24] ),
    .A2(_06159_),
    .B1(_05770_),
    .B2(_06160_),
    .X(_03196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09944_ (.A1(\design_top.core0.REG1[14][23] ),
    .A2(_06159_),
    .B1(_05772_),
    .B2(_06160_),
    .X(_03195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09945_ (.A(_06154_),
    .X(_06161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09946_ (.A1(\design_top.core0.REG1[14][22] ),
    .A2(_06161_),
    .B1(_05774_),
    .B2(_06160_),
    .X(_03194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09947_ (.A(_06157_),
    .X(_06162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09948_ (.A1(\design_top.core0.REG1[14][21] ),
    .A2(_06161_),
    .B1(_05776_),
    .B2(_06162_),
    .X(_03193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09949_ (.A1(\design_top.core0.REG1[14][20] ),
    .A2(_06161_),
    .B1(_05778_),
    .B2(_06162_),
    .X(_03192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09950_ (.A1(\design_top.core0.REG1[14][19] ),
    .A2(_06161_),
    .B1(_05782_),
    .B2(_06162_),
    .X(_03191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09951_ (.A1(\design_top.core0.REG1[14][18] ),
    .A2(_06161_),
    .B1(_05784_),
    .B2(_06162_),
    .X(_03190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09952_ (.A(_06153_),
    .X(_06163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09953_ (.A1(\design_top.core0.REG1[14][17] ),
    .A2(_06163_),
    .B1(_05786_),
    .B2(_06162_),
    .X(_03189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09954_ (.A(_06156_),
    .X(_06164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09955_ (.A1(\design_top.core0.REG1[14][16] ),
    .A2(_06163_),
    .B1(_05788_),
    .B2(_06164_),
    .X(_03188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09956_ (.A1(\design_top.core0.REG1[14][15] ),
    .A2(_06163_),
    .B1(_05790_),
    .B2(_06164_),
    .X(_03187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09957_ (.A1(\design_top.core0.REG1[14][14] ),
    .A2(_06163_),
    .B1(_05794_),
    .B2(_06164_),
    .X(_03186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _09958_ (.A1(\design_top.core0.REG1[14][13] ),
    .A2(_06157_),
    .B1(_05655_),
    .B2(_06155_),
    .X(_03185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09959_ (.A1(\design_top.core0.REG1[14][12] ),
    .A2(_06163_),
    .B1(_05796_),
    .B2(_06164_),
    .X(_03184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09960_ (.A(_06153_),
    .X(_06165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09961_ (.A1(\design_top.core0.REG1[14][11] ),
    .A2(_06165_),
    .B1(_05798_),
    .B2(_06164_),
    .X(_03183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09962_ (.A(_06156_),
    .X(_06166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09963_ (.A1(\design_top.core0.REG1[14][10] ),
    .A2(_06165_),
    .B1(_05800_),
    .B2(_06166_),
    .X(_03182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09964_ (.A1(\design_top.core0.REG1[14][9] ),
    .A2(_06165_),
    .B1(_05802_),
    .B2(_06166_),
    .X(_03181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09965_ (.A1(\design_top.core0.REG1[14][8] ),
    .A2(_06165_),
    .B1(_05806_),
    .B2(_06166_),
    .X(_03180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09966_ (.A1(\design_top.core0.REG1[14][7] ),
    .A2(_06165_),
    .B1(_05808_),
    .B2(_06166_),
    .X(_03179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09967_ (.A(_06153_),
    .X(_06167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09968_ (.A1(\design_top.core0.REG1[14][6] ),
    .A2(_06167_),
    .B1(_05810_),
    .B2(_06166_),
    .X(_03178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09969_ (.A(_06156_),
    .X(_06168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09970_ (.A1(\design_top.core0.REG1[14][5] ),
    .A2(_06167_),
    .B1(_05812_),
    .B2(_06168_),
    .X(_03177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09971_ (.A1(\design_top.core0.REG1[14][4] ),
    .A2(_06167_),
    .B1(_05814_),
    .B2(_06168_),
    .X(_03176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09972_ (.A1(\design_top.core0.REG1[14][3] ),
    .A2(_06167_),
    .B1(_05818_),
    .B2(_06168_),
    .X(_03175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09973_ (.A1(\design_top.core0.REG1[14][2] ),
    .A2(_06167_),
    .B1(_05820_),
    .B2(_06168_),
    .X(_03174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09974_ (.A1(\design_top.core0.REG1[14][1] ),
    .A2(_06154_),
    .B1(_05822_),
    .B2(_06168_),
    .X(_03173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09975_ (.A1(\design_top.core0.REG1[14][0] ),
    .A2(_06154_),
    .B1(_05824_),
    .B2(_06157_),
    .X(_03172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _09976_ (.A(_05206_),
    .B(_06049_),
    .Y(_00557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09977_ (.A(_05209_),
    .B(_00557_),
    .X(_06169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09978_ (.A(_06169_),
    .X(_06170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09979_ (.A(_06169_),
    .Y(_06171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09980_ (.A(_06171_),
    .X(_06172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09981_ (.A1(_00268_),
    .A2(_06170_),
    .B1(\design_top.MEM[5][7] ),
    .B2(_06172_),
    .X(_03171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09982_ (.A1(_00267_),
    .A2(_06170_),
    .B1(\design_top.MEM[5][6] ),
    .B2(_06172_),
    .X(_03170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09983_ (.A1(_00266_),
    .A2(_06170_),
    .B1(\design_top.MEM[5][5] ),
    .B2(_06172_),
    .X(_03169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09984_ (.A1(_00265_),
    .A2(_06170_),
    .B1(\design_top.MEM[5][4] ),
    .B2(_06172_),
    .X(_03168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09985_ (.A1(_00264_),
    .A2(_06170_),
    .B1(\design_top.MEM[5][3] ),
    .B2(_06172_),
    .X(_03167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09986_ (.A1(_00263_),
    .A2(_06169_),
    .B1(\design_top.MEM[5][2] ),
    .B2(_06171_),
    .X(_03166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09987_ (.A1(_00262_),
    .A2(_06169_),
    .B1(\design_top.MEM[5][1] ),
    .B2(_06171_),
    .X(_03165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09988_ (.A1(_00261_),
    .A2(_06169_),
    .B1(\design_top.MEM[5][0] ),
    .B2(_06171_),
    .X(_03164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _09989_ (.A(_05220_),
    .B(_06049_),
    .Y(_00556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09990_ (.A(_05223_),
    .B(_00556_),
    .X(_06173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09991_ (.A(_06173_),
    .X(_06174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09992_ (.A(_06173_),
    .Y(_06175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09993_ (.A(_06175_),
    .X(_06176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09994_ (.A1(_00276_),
    .A2(_06174_),
    .B1(\design_top.MEM[6][7] ),
    .B2(_06176_),
    .X(_03163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09995_ (.A1(_00275_),
    .A2(_06174_),
    .B1(\design_top.MEM[6][6] ),
    .B2(_06176_),
    .X(_03162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09996_ (.A1(_00274_),
    .A2(_06174_),
    .B1(\design_top.MEM[6][5] ),
    .B2(_06176_),
    .X(_03161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09997_ (.A1(_00273_),
    .A2(_06174_),
    .B1(\design_top.MEM[6][4] ),
    .B2(_06176_),
    .X(_03160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09998_ (.A1(_00272_),
    .A2(_06174_),
    .B1(\design_top.MEM[6][3] ),
    .B2(_06176_),
    .X(_03159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _09999_ (.A1(_00271_),
    .A2(_06173_),
    .B1(\design_top.MEM[6][2] ),
    .B2(_06175_),
    .X(_03158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10000_ (.A1(_00270_),
    .A2(_06173_),
    .B1(\design_top.MEM[6][1] ),
    .B2(_06175_),
    .X(_03157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10001_ (.A1(_00269_),
    .A2(_06173_),
    .B1(\design_top.MEM[6][0] ),
    .B2(_06175_),
    .X(_03156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10002_ (.A(_05749_),
    .X(_06177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10003_ (.A(_05846_),
    .X(_06178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10004_ (.A(_06178_),
    .X(_06179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10005_ (.A(_06179_),
    .X(_06180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10006_ (.A(_06178_),
    .Y(_06181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10007_ (.A(_06181_),
    .X(_06182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10008_ (.A(_06182_),
    .X(_06183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10009_ (.A1(_06177_),
    .A2(_06180_),
    .B1(\design_top.core0.REG2[15][31] ),
    .B2(_06183_),
    .X(_03155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10010_ (.A(_05753_),
    .X(_06184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10011_ (.A1(_06184_),
    .A2(_06180_),
    .B1(\design_top.core0.REG2[15][30] ),
    .B2(_06183_),
    .X(_03154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10012_ (.A(_05757_),
    .X(_06185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10013_ (.A1(_06185_),
    .A2(_06180_),
    .B1(\design_top.core0.REG2[15][29] ),
    .B2(_06183_),
    .X(_03153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10014_ (.A(_05759_),
    .X(_06186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10015_ (.A1(_06186_),
    .A2(_06180_),
    .B1(\design_top.core0.REG2[15][28] ),
    .B2(_06183_),
    .X(_03152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10016_ (.A(_05761_),
    .X(_06187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10017_ (.A1(_06187_),
    .A2(_06180_),
    .B1(\design_top.core0.REG2[15][27] ),
    .B2(_06183_),
    .X(_03151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10018_ (.A(_05763_),
    .X(_06188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10019_ (.A(_06179_),
    .X(_06189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10020_ (.A(_06182_),
    .X(_06190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10021_ (.A1(_06188_),
    .A2(_06189_),
    .B1(\design_top.core0.REG2[15][26] ),
    .B2(_06190_),
    .X(_03150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10022_ (.A(_05765_),
    .X(_06191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10023_ (.A1(_06191_),
    .A2(_06189_),
    .B1(\design_top.core0.REG2[15][25] ),
    .B2(_06190_),
    .X(_03149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10024_ (.A(_05769_),
    .X(_06192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10025_ (.A1(_06192_),
    .A2(_06189_),
    .B1(\design_top.core0.REG2[15][24] ),
    .B2(_06190_),
    .X(_03148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10026_ (.A(_05771_),
    .X(_06193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10027_ (.A1(_06193_),
    .A2(_06189_),
    .B1(\design_top.core0.REG2[15][23] ),
    .B2(_06190_),
    .X(_03147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10028_ (.A(_05773_),
    .X(_06194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10029_ (.A1(_06194_),
    .A2(_06189_),
    .B1(\design_top.core0.REG2[15][22] ),
    .B2(_06190_),
    .X(_03146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10030_ (.A(_05775_),
    .X(_06195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10031_ (.A(_06179_),
    .X(_06196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10032_ (.A(_06182_),
    .X(_06197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10033_ (.A1(_06195_),
    .A2(_06196_),
    .B1(\design_top.core0.REG2[15][21] ),
    .B2(_06197_),
    .X(_03145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10034_ (.A(_05777_),
    .X(_06198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10035_ (.A1(_06198_),
    .A2(_06196_),
    .B1(\design_top.core0.REG2[15][20] ),
    .B2(_06197_),
    .X(_03144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10036_ (.A(_05781_),
    .X(_06199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10037_ (.A1(_06199_),
    .A2(_06196_),
    .B1(\design_top.core0.REG2[15][19] ),
    .B2(_06197_),
    .X(_03143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10038_ (.A(_05783_),
    .X(_06200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10039_ (.A1(_06200_),
    .A2(_06196_),
    .B1(\design_top.core0.REG2[15][18] ),
    .B2(_06197_),
    .X(_03142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10040_ (.A(_05785_),
    .X(_06201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10041_ (.A1(_06201_),
    .A2(_06196_),
    .B1(\design_top.core0.REG2[15][17] ),
    .B2(_06197_),
    .X(_03141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10042_ (.A(_05787_),
    .X(_06202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10043_ (.A(_06178_),
    .X(_06203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10044_ (.A(_06181_),
    .X(_06204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10045_ (.A1(_06202_),
    .A2(_06203_),
    .B1(\design_top.core0.REG2[15][16] ),
    .B2(_06204_),
    .X(_03140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10046_ (.A(_05789_),
    .X(_06205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10047_ (.A1(_06205_),
    .A2(_06203_),
    .B1(\design_top.core0.REG2[15][15] ),
    .B2(_06204_),
    .X(_03139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10048_ (.A(_05793_),
    .X(_06206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10049_ (.A1(_06206_),
    .A2(_06203_),
    .B1(\design_top.core0.REG2[15][14] ),
    .B2(_06204_),
    .X(_03138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10050_ (.A1(\design_top.core0.REG2[15][13] ),
    .A2(_06179_),
    .B1(_05656_),
    .B2(_06182_),
    .X(_03137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10051_ (.A(_05795_),
    .X(_06207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10052_ (.A1(_06207_),
    .A2(_06203_),
    .B1(\design_top.core0.REG2[15][12] ),
    .B2(_06204_),
    .X(_03136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10053_ (.A(_05797_),
    .X(_06208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10054_ (.A1(_06208_),
    .A2(_06203_),
    .B1(\design_top.core0.REG2[15][11] ),
    .B2(_06204_),
    .X(_03135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10055_ (.A(_05799_),
    .X(_06209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10056_ (.A(_06178_),
    .X(_06210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10057_ (.A(_06181_),
    .X(_06211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10058_ (.A1(_06209_),
    .A2(_06210_),
    .B1(\design_top.core0.REG2[15][10] ),
    .B2(_06211_),
    .X(_03134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10059_ (.A(_05801_),
    .X(_06212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10060_ (.A1(_06212_),
    .A2(_06210_),
    .B1(\design_top.core0.REG2[15][9] ),
    .B2(_06211_),
    .X(_03133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10061_ (.A(_05805_),
    .X(_06213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10062_ (.A1(_06213_),
    .A2(_06210_),
    .B1(\design_top.core0.REG2[15][8] ),
    .B2(_06211_),
    .X(_03132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10063_ (.A(_05807_),
    .X(_06214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10064_ (.A1(_06214_),
    .A2(_06210_),
    .B1(\design_top.core0.REG2[15][7] ),
    .B2(_06211_),
    .X(_03131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10065_ (.A(_05809_),
    .X(_06215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10066_ (.A1(_06215_),
    .A2(_06210_),
    .B1(\design_top.core0.REG2[15][6] ),
    .B2(_06211_),
    .X(_03130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10067_ (.A(_05811_),
    .X(_06216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10068_ (.A(_06178_),
    .X(_06217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10069_ (.A(_06181_),
    .X(_06218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10070_ (.A1(_06216_),
    .A2(_06217_),
    .B1(\design_top.core0.REG2[15][5] ),
    .B2(_06218_),
    .X(_03129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10071_ (.A(_05813_),
    .X(_06219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10072_ (.A1(_06219_),
    .A2(_06217_),
    .B1(\design_top.core0.REG2[15][4] ),
    .B2(_06218_),
    .X(_03128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10073_ (.A(_05817_),
    .X(_06220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10074_ (.A1(_06220_),
    .A2(_06217_),
    .B1(\design_top.core0.REG2[15][3] ),
    .B2(_06218_),
    .X(_03127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10075_ (.A(_05819_),
    .X(_06221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10076_ (.A1(_06221_),
    .A2(_06217_),
    .B1(\design_top.core0.REG2[15][2] ),
    .B2(_06218_),
    .X(_03126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10077_ (.A(_05821_),
    .X(_06222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10078_ (.A1(_06222_),
    .A2(_06217_),
    .B1(\design_top.core0.REG2[15][1] ),
    .B2(_06218_),
    .X(_03125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10079_ (.A(_05823_),
    .X(_06223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10080_ (.A1(_06223_),
    .A2(_06179_),
    .B1(\design_top.core0.REG2[15][0] ),
    .B2(_06182_),
    .X(_03124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10081_ (.A(_05895_),
    .X(_06224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10082_ (.A(_06224_),
    .X(_06225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10083_ (.A(_06225_),
    .X(_06226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10084_ (.A(_06224_),
    .Y(_06227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10085_ (.A(_06227_),
    .X(_06228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10086_ (.A(_06228_),
    .X(_06229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10087_ (.A1(_06177_),
    .A2(_06226_),
    .B1(\design_top.core0.REG2[1][31] ),
    .B2(_06229_),
    .X(_03123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10088_ (.A1(_06184_),
    .A2(_06226_),
    .B1(\design_top.core0.REG2[1][30] ),
    .B2(_06229_),
    .X(_03122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10089_ (.A1(_06185_),
    .A2(_06226_),
    .B1(\design_top.core0.REG2[1][29] ),
    .B2(_06229_),
    .X(_03121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10090_ (.A1(_06186_),
    .A2(_06226_),
    .B1(\design_top.core0.REG2[1][28] ),
    .B2(_06229_),
    .X(_03120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10091_ (.A1(_06187_),
    .A2(_06226_),
    .B1(\design_top.core0.REG2[1][27] ),
    .B2(_06229_),
    .X(_03119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10092_ (.A(_06225_),
    .X(_06230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10093_ (.A(_06228_),
    .X(_06231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10094_ (.A1(_06188_),
    .A2(_06230_),
    .B1(\design_top.core0.REG2[1][26] ),
    .B2(_06231_),
    .X(_03118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10095_ (.A1(_06191_),
    .A2(_06230_),
    .B1(\design_top.core0.REG2[1][25] ),
    .B2(_06231_),
    .X(_03117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10096_ (.A1(_06192_),
    .A2(_06230_),
    .B1(\design_top.core0.REG2[1][24] ),
    .B2(_06231_),
    .X(_03116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10097_ (.A1(_06193_),
    .A2(_06230_),
    .B1(\design_top.core0.REG2[1][23] ),
    .B2(_06231_),
    .X(_03115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10098_ (.A1(_06194_),
    .A2(_06230_),
    .B1(\design_top.core0.REG2[1][22] ),
    .B2(_06231_),
    .X(_03114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10099_ (.A(_06225_),
    .X(_06232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10100_ (.A(_06228_),
    .X(_06233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10101_ (.A1(_06195_),
    .A2(_06232_),
    .B1(\design_top.core0.REG2[1][21] ),
    .B2(_06233_),
    .X(_03113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10102_ (.A1(_06198_),
    .A2(_06232_),
    .B1(\design_top.core0.REG2[1][20] ),
    .B2(_06233_),
    .X(_03112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10103_ (.A1(_06199_),
    .A2(_06232_),
    .B1(\design_top.core0.REG2[1][19] ),
    .B2(_06233_),
    .X(_03111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10104_ (.A1(_06200_),
    .A2(_06232_),
    .B1(\design_top.core0.REG2[1][18] ),
    .B2(_06233_),
    .X(_03110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10105_ (.A1(_06201_),
    .A2(_06232_),
    .B1(\design_top.core0.REG2[1][17] ),
    .B2(_06233_),
    .X(_03109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10106_ (.A(_06224_),
    .X(_06234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10107_ (.A(_06227_),
    .X(_06235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10108_ (.A1(_06202_),
    .A2(_06234_),
    .B1(\design_top.core0.REG2[1][16] ),
    .B2(_06235_),
    .X(_03108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10109_ (.A1(_06205_),
    .A2(_06234_),
    .B1(\design_top.core0.REG2[1][15] ),
    .B2(_06235_),
    .X(_03107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10110_ (.A1(_06206_),
    .A2(_06234_),
    .B1(\design_top.core0.REG2[1][14] ),
    .B2(_06235_),
    .X(_03106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10111_ (.A1(\design_top.core0.REG2[1][13] ),
    .A2(_06225_),
    .B1(_05656_),
    .B2(_06228_),
    .X(_03105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10112_ (.A1(_06207_),
    .A2(_06234_),
    .B1(\design_top.core0.REG2[1][12] ),
    .B2(_06235_),
    .X(_03104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10113_ (.A1(_06208_),
    .A2(_06234_),
    .B1(\design_top.core0.REG2[1][11] ),
    .B2(_06235_),
    .X(_03103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10114_ (.A(_06224_),
    .X(_06236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10115_ (.A(_06227_),
    .X(_06237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10116_ (.A1(_06209_),
    .A2(_06236_),
    .B1(\design_top.core0.REG2[1][10] ),
    .B2(_06237_),
    .X(_03102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10117_ (.A1(_06212_),
    .A2(_06236_),
    .B1(\design_top.core0.REG2[1][9] ),
    .B2(_06237_),
    .X(_03101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10118_ (.A1(_06213_),
    .A2(_06236_),
    .B1(\design_top.core0.REG2[1][8] ),
    .B2(_06237_),
    .X(_03100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10119_ (.A1(_06214_),
    .A2(_06236_),
    .B1(\design_top.core0.REG2[1][7] ),
    .B2(_06237_),
    .X(_03099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10120_ (.A1(_06215_),
    .A2(_06236_),
    .B1(\design_top.core0.REG2[1][6] ),
    .B2(_06237_),
    .X(_03098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10121_ (.A(_06224_),
    .X(_06238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10122_ (.A(_06227_),
    .X(_06239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10123_ (.A1(_06216_),
    .A2(_06238_),
    .B1(\design_top.core0.REG2[1][5] ),
    .B2(_06239_),
    .X(_03097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10124_ (.A1(_06219_),
    .A2(_06238_),
    .B1(\design_top.core0.REG2[1][4] ),
    .B2(_06239_),
    .X(_03096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10125_ (.A1(_06220_),
    .A2(_06238_),
    .B1(\design_top.core0.REG2[1][3] ),
    .B2(_06239_),
    .X(_03095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10126_ (.A1(_06221_),
    .A2(_06238_),
    .B1(\design_top.core0.REG2[1][2] ),
    .B2(_06239_),
    .X(_03094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10127_ (.A1(_06222_),
    .A2(_06238_),
    .B1(\design_top.core0.REG2[1][1] ),
    .B2(_06239_),
    .X(_03093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10128_ (.A1(_06223_),
    .A2(_06225_),
    .B1(\design_top.core0.REG2[1][0] ),
    .B2(_06228_),
    .X(_03092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10129_ (.A(_05914_),
    .X(_06240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10130_ (.A(_06240_),
    .X(_06241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10131_ (.A(_06241_),
    .X(_06242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10132_ (.A(_06240_),
    .Y(_06243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10133_ (.A(_06243_),
    .X(_06244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10134_ (.A(_06244_),
    .X(_06245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10135_ (.A1(_06177_),
    .A2(_06242_),
    .B1(\design_top.core0.REG2[2][31] ),
    .B2(_06245_),
    .X(_03091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10136_ (.A1(_06184_),
    .A2(_06242_),
    .B1(\design_top.core0.REG2[2][30] ),
    .B2(_06245_),
    .X(_03090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10137_ (.A1(_06185_),
    .A2(_06242_),
    .B1(\design_top.core0.REG2[2][29] ),
    .B2(_06245_),
    .X(_03089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10138_ (.A1(_06186_),
    .A2(_06242_),
    .B1(\design_top.core0.REG2[2][28] ),
    .B2(_06245_),
    .X(_03088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10139_ (.A1(_06187_),
    .A2(_06242_),
    .B1(\design_top.core0.REG2[2][27] ),
    .B2(_06245_),
    .X(_03087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10140_ (.A(_06241_),
    .X(_06246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10141_ (.A(_06244_),
    .X(_06247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10142_ (.A1(_06188_),
    .A2(_06246_),
    .B1(\design_top.core0.REG2[2][26] ),
    .B2(_06247_),
    .X(_03086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10143_ (.A1(_06191_),
    .A2(_06246_),
    .B1(\design_top.core0.REG2[2][25] ),
    .B2(_06247_),
    .X(_03085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10144_ (.A1(_06192_),
    .A2(_06246_),
    .B1(\design_top.core0.REG2[2][24] ),
    .B2(_06247_),
    .X(_03084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10145_ (.A1(_06193_),
    .A2(_06246_),
    .B1(\design_top.core0.REG2[2][23] ),
    .B2(_06247_),
    .X(_03083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10146_ (.A1(_06194_),
    .A2(_06246_),
    .B1(\design_top.core0.REG2[2][22] ),
    .B2(_06247_),
    .X(_03082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10147_ (.A(_06241_),
    .X(_06248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10148_ (.A(_06244_),
    .X(_06249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10149_ (.A1(_06195_),
    .A2(_06248_),
    .B1(\design_top.core0.REG2[2][21] ),
    .B2(_06249_),
    .X(_03081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10150_ (.A1(_06198_),
    .A2(_06248_),
    .B1(\design_top.core0.REG2[2][20] ),
    .B2(_06249_),
    .X(_03080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10151_ (.A1(_06199_),
    .A2(_06248_),
    .B1(\design_top.core0.REG2[2][19] ),
    .B2(_06249_),
    .X(_03079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10152_ (.A1(_06200_),
    .A2(_06248_),
    .B1(\design_top.core0.REG2[2][18] ),
    .B2(_06249_),
    .X(_03078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10153_ (.A1(_06201_),
    .A2(_06248_),
    .B1(\design_top.core0.REG2[2][17] ),
    .B2(_06249_),
    .X(_03077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10154_ (.A(_06240_),
    .X(_06250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10155_ (.A(_06243_),
    .X(_06251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10156_ (.A1(_06202_),
    .A2(_06250_),
    .B1(\design_top.core0.REG2[2][16] ),
    .B2(_06251_),
    .X(_03076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10157_ (.A1(_06205_),
    .A2(_06250_),
    .B1(\design_top.core0.REG2[2][15] ),
    .B2(_06251_),
    .X(_03075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10158_ (.A1(_06206_),
    .A2(_06250_),
    .B1(\design_top.core0.REG2[2][14] ),
    .B2(_06251_),
    .X(_03074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10159_ (.A1(\design_top.core0.REG2[2][13] ),
    .A2(_06241_),
    .B1(_05656_),
    .B2(_06244_),
    .X(_03073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10160_ (.A1(_06207_),
    .A2(_06250_),
    .B1(\design_top.core0.REG2[2][12] ),
    .B2(_06251_),
    .X(_03072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10161_ (.A1(_06208_),
    .A2(_06250_),
    .B1(\design_top.core0.REG2[2][11] ),
    .B2(_06251_),
    .X(_03071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10162_ (.A(_06240_),
    .X(_06252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10163_ (.A(_06243_),
    .X(_06253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10164_ (.A1(_06209_),
    .A2(_06252_),
    .B1(\design_top.core0.REG2[2][10] ),
    .B2(_06253_),
    .X(_03070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10165_ (.A1(_06212_),
    .A2(_06252_),
    .B1(\design_top.core0.REG2[2][9] ),
    .B2(_06253_),
    .X(_03069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10166_ (.A1(_06213_),
    .A2(_06252_),
    .B1(\design_top.core0.REG2[2][8] ),
    .B2(_06253_),
    .X(_03068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10167_ (.A1(_06214_),
    .A2(_06252_),
    .B1(\design_top.core0.REG2[2][7] ),
    .B2(_06253_),
    .X(_03067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10168_ (.A1(_06215_),
    .A2(_06252_),
    .B1(\design_top.core0.REG2[2][6] ),
    .B2(_06253_),
    .X(_03066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10169_ (.A(_06240_),
    .X(_06254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10170_ (.A(_06243_),
    .X(_06255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10171_ (.A1(_06216_),
    .A2(_06254_),
    .B1(\design_top.core0.REG2[2][5] ),
    .B2(_06255_),
    .X(_03065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10172_ (.A1(_06219_),
    .A2(_06254_),
    .B1(\design_top.core0.REG2[2][4] ),
    .B2(_06255_),
    .X(_03064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10173_ (.A1(_06220_),
    .A2(_06254_),
    .B1(\design_top.core0.REG2[2][3] ),
    .B2(_06255_),
    .X(_03063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10174_ (.A1(_06221_),
    .A2(_06254_),
    .B1(\design_top.core0.REG2[2][2] ),
    .B2(_06255_),
    .X(_03062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10175_ (.A1(_06222_),
    .A2(_06254_),
    .B1(\design_top.core0.REG2[2][1] ),
    .B2(_06255_),
    .X(_03061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10176_ (.A1(_06223_),
    .A2(_06241_),
    .B1(\design_top.core0.REG2[2][0] ),
    .B2(_06244_),
    .X(_03060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10177_ (.A(_05932_),
    .X(_06256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10178_ (.A(_06256_),
    .X(_06257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10179_ (.A(_06257_),
    .X(_06258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10180_ (.A(_06256_),
    .Y(_06259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10181_ (.A(_06259_),
    .X(_06260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10182_ (.A(_06260_),
    .X(_06261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10183_ (.A1(_06177_),
    .A2(_06258_),
    .B1(\design_top.core0.REG2[3][31] ),
    .B2(_06261_),
    .X(_03059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10184_ (.A1(_06184_),
    .A2(_06258_),
    .B1(\design_top.core0.REG2[3][30] ),
    .B2(_06261_),
    .X(_03058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10185_ (.A1(_06185_),
    .A2(_06258_),
    .B1(\design_top.core0.REG2[3][29] ),
    .B2(_06261_),
    .X(_03057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10186_ (.A1(_06186_),
    .A2(_06258_),
    .B1(\design_top.core0.REG2[3][28] ),
    .B2(_06261_),
    .X(_03056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10187_ (.A1(_06187_),
    .A2(_06258_),
    .B1(\design_top.core0.REG2[3][27] ),
    .B2(_06261_),
    .X(_03055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10188_ (.A(_06257_),
    .X(_06262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10189_ (.A(_06260_),
    .X(_06263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10190_ (.A1(_06188_),
    .A2(_06262_),
    .B1(\design_top.core0.REG2[3][26] ),
    .B2(_06263_),
    .X(_03054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10191_ (.A1(_06191_),
    .A2(_06262_),
    .B1(\design_top.core0.REG2[3][25] ),
    .B2(_06263_),
    .X(_03053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10192_ (.A1(_06192_),
    .A2(_06262_),
    .B1(\design_top.core0.REG2[3][24] ),
    .B2(_06263_),
    .X(_03052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10193_ (.A1(_06193_),
    .A2(_06262_),
    .B1(\design_top.core0.REG2[3][23] ),
    .B2(_06263_),
    .X(_03051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10194_ (.A1(_06194_),
    .A2(_06262_),
    .B1(\design_top.core0.REG2[3][22] ),
    .B2(_06263_),
    .X(_03050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10195_ (.A(_06257_),
    .X(_06264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10196_ (.A(_06260_),
    .X(_06265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10197_ (.A1(_06195_),
    .A2(_06264_),
    .B1(\design_top.core0.REG2[3][21] ),
    .B2(_06265_),
    .X(_03049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10198_ (.A1(_06198_),
    .A2(_06264_),
    .B1(\design_top.core0.REG2[3][20] ),
    .B2(_06265_),
    .X(_03048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10199_ (.A1(_06199_),
    .A2(_06264_),
    .B1(\design_top.core0.REG2[3][19] ),
    .B2(_06265_),
    .X(_03047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10200_ (.A1(_06200_),
    .A2(_06264_),
    .B1(\design_top.core0.REG2[3][18] ),
    .B2(_06265_),
    .X(_03046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10201_ (.A1(_06201_),
    .A2(_06264_),
    .B1(\design_top.core0.REG2[3][17] ),
    .B2(_06265_),
    .X(_03045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10202_ (.A(_06256_),
    .X(_06266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10203_ (.A(_06259_),
    .X(_06267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10204_ (.A1(_06202_),
    .A2(_06266_),
    .B1(\design_top.core0.REG2[3][16] ),
    .B2(_06267_),
    .X(_03044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10205_ (.A1(_06205_),
    .A2(_06266_),
    .B1(\design_top.core0.REG2[3][15] ),
    .B2(_06267_),
    .X(_03043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10206_ (.A1(_06206_),
    .A2(_06266_),
    .B1(\design_top.core0.REG2[3][14] ),
    .B2(_06267_),
    .X(_03042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10207_ (.A(_05655_),
    .X(_06268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10208_ (.A1(\design_top.core0.REG2[3][13] ),
    .A2(_06257_),
    .B1(_06268_),
    .B2(_06260_),
    .X(_03041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10209_ (.A1(_06207_),
    .A2(_06266_),
    .B1(\design_top.core0.REG2[3][12] ),
    .B2(_06267_),
    .X(_03040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10210_ (.A1(_06208_),
    .A2(_06266_),
    .B1(\design_top.core0.REG2[3][11] ),
    .B2(_06267_),
    .X(_03039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10211_ (.A(_06256_),
    .X(_06269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10212_ (.A(_06259_),
    .X(_06270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10213_ (.A1(_06209_),
    .A2(_06269_),
    .B1(\design_top.core0.REG2[3][10] ),
    .B2(_06270_),
    .X(_03038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10214_ (.A1(_06212_),
    .A2(_06269_),
    .B1(\design_top.core0.REG2[3][9] ),
    .B2(_06270_),
    .X(_03037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10215_ (.A1(_06213_),
    .A2(_06269_),
    .B1(\design_top.core0.REG2[3][8] ),
    .B2(_06270_),
    .X(_03036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10216_ (.A1(_06214_),
    .A2(_06269_),
    .B1(\design_top.core0.REG2[3][7] ),
    .B2(_06270_),
    .X(_03035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10217_ (.A1(_06215_),
    .A2(_06269_),
    .B1(\design_top.core0.REG2[3][6] ),
    .B2(_06270_),
    .X(_03034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10218_ (.A(_06256_),
    .X(_06271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10219_ (.A(_06259_),
    .X(_06272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10220_ (.A1(_06216_),
    .A2(_06271_),
    .B1(\design_top.core0.REG2[3][5] ),
    .B2(_06272_),
    .X(_03033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10221_ (.A1(_06219_),
    .A2(_06271_),
    .B1(\design_top.core0.REG2[3][4] ),
    .B2(_06272_),
    .X(_03032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10222_ (.A1(_06220_),
    .A2(_06271_),
    .B1(\design_top.core0.REG2[3][3] ),
    .B2(_06272_),
    .X(_03031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10223_ (.A1(_06221_),
    .A2(_06271_),
    .B1(\design_top.core0.REG2[3][2] ),
    .B2(_06272_),
    .X(_03030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10224_ (.A1(_06222_),
    .A2(_06271_),
    .B1(\design_top.core0.REG2[3][1] ),
    .B2(_06272_),
    .X(_03029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10225_ (.A1(_06223_),
    .A2(_06257_),
    .B1(\design_top.core0.REG2[3][0] ),
    .B2(_06260_),
    .X(_03028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10226_ (.A(_05950_),
    .X(_06273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10227_ (.A(_06273_),
    .X(_06274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10228_ (.A(_06274_),
    .X(_06275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10229_ (.A(_06273_),
    .Y(_06276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10230_ (.A(_06276_),
    .X(_06277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10231_ (.A(_06277_),
    .X(_06278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10232_ (.A1(_06177_),
    .A2(_06275_),
    .B1(\design_top.core0.REG2[4][31] ),
    .B2(_06278_),
    .X(_03027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10233_ (.A1(_06184_),
    .A2(_06275_),
    .B1(\design_top.core0.REG2[4][30] ),
    .B2(_06278_),
    .X(_03026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10234_ (.A1(_06185_),
    .A2(_06275_),
    .B1(\design_top.core0.REG2[4][29] ),
    .B2(_06278_),
    .X(_03025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10235_ (.A1(_06186_),
    .A2(_06275_),
    .B1(\design_top.core0.REG2[4][28] ),
    .B2(_06278_),
    .X(_03024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10236_ (.A1(_06187_),
    .A2(_06275_),
    .B1(\design_top.core0.REG2[4][27] ),
    .B2(_06278_),
    .X(_03023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10237_ (.A(_06274_),
    .X(_06279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10238_ (.A(_06277_),
    .X(_06280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10239_ (.A1(_06188_),
    .A2(_06279_),
    .B1(\design_top.core0.REG2[4][26] ),
    .B2(_06280_),
    .X(_03022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10240_ (.A1(_06191_),
    .A2(_06279_),
    .B1(\design_top.core0.REG2[4][25] ),
    .B2(_06280_),
    .X(_03021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10241_ (.A1(_06192_),
    .A2(_06279_),
    .B1(\design_top.core0.REG2[4][24] ),
    .B2(_06280_),
    .X(_03020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10242_ (.A1(_06193_),
    .A2(_06279_),
    .B1(\design_top.core0.REG2[4][23] ),
    .B2(_06280_),
    .X(_03019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10243_ (.A1(_06194_),
    .A2(_06279_),
    .B1(\design_top.core0.REG2[4][22] ),
    .B2(_06280_),
    .X(_03018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10244_ (.A(_06274_),
    .X(_06281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10245_ (.A(_06277_),
    .X(_06282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10246_ (.A1(_06195_),
    .A2(_06281_),
    .B1(\design_top.core0.REG2[4][21] ),
    .B2(_06282_),
    .X(_03017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10247_ (.A1(_06198_),
    .A2(_06281_),
    .B1(\design_top.core0.REG2[4][20] ),
    .B2(_06282_),
    .X(_03016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10248_ (.A1(_06199_),
    .A2(_06281_),
    .B1(\design_top.core0.REG2[4][19] ),
    .B2(_06282_),
    .X(_03015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10249_ (.A1(_06200_),
    .A2(_06281_),
    .B1(\design_top.core0.REG2[4][18] ),
    .B2(_06282_),
    .X(_03014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10250_ (.A1(_06201_),
    .A2(_06281_),
    .B1(\design_top.core0.REG2[4][17] ),
    .B2(_06282_),
    .X(_03013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10251_ (.A(_06273_),
    .X(_06283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10252_ (.A(_06276_),
    .X(_06284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10253_ (.A1(_06202_),
    .A2(_06283_),
    .B1(\design_top.core0.REG2[4][16] ),
    .B2(_06284_),
    .X(_03012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10254_ (.A1(_06205_),
    .A2(_06283_),
    .B1(\design_top.core0.REG2[4][15] ),
    .B2(_06284_),
    .X(_03011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10255_ (.A1(_06206_),
    .A2(_06283_),
    .B1(\design_top.core0.REG2[4][14] ),
    .B2(_06284_),
    .X(_03010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10256_ (.A1(\design_top.core0.REG2[4][13] ),
    .A2(_06274_),
    .B1(_06268_),
    .B2(_06277_),
    .X(_03009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10257_ (.A1(_06207_),
    .A2(_06283_),
    .B1(\design_top.core0.REG2[4][12] ),
    .B2(_06284_),
    .X(_03008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10258_ (.A1(_06208_),
    .A2(_06283_),
    .B1(\design_top.core0.REG2[4][11] ),
    .B2(_06284_),
    .X(_03007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10259_ (.A(_06273_),
    .X(_06285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10260_ (.A(_06276_),
    .X(_06286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10261_ (.A1(_06209_),
    .A2(_06285_),
    .B1(\design_top.core0.REG2[4][10] ),
    .B2(_06286_),
    .X(_03006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10262_ (.A1(_06212_),
    .A2(_06285_),
    .B1(\design_top.core0.REG2[4][9] ),
    .B2(_06286_),
    .X(_03005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10263_ (.A1(_06213_),
    .A2(_06285_),
    .B1(\design_top.core0.REG2[4][8] ),
    .B2(_06286_),
    .X(_03004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10264_ (.A1(_06214_),
    .A2(_06285_),
    .B1(\design_top.core0.REG2[4][7] ),
    .B2(_06286_),
    .X(_03003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10265_ (.A1(_06215_),
    .A2(_06285_),
    .B1(\design_top.core0.REG2[4][6] ),
    .B2(_06286_),
    .X(_03002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10266_ (.A(_06273_),
    .X(_06287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10267_ (.A(_06276_),
    .X(_06288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10268_ (.A1(_06216_),
    .A2(_06287_),
    .B1(\design_top.core0.REG2[4][5] ),
    .B2(_06288_),
    .X(_03001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10269_ (.A1(_06219_),
    .A2(_06287_),
    .B1(\design_top.core0.REG2[4][4] ),
    .B2(_06288_),
    .X(_03000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10270_ (.A1(_06220_),
    .A2(_06287_),
    .B1(\design_top.core0.REG2[4][3] ),
    .B2(_06288_),
    .X(_02999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10271_ (.A1(_06221_),
    .A2(_06287_),
    .B1(\design_top.core0.REG2[4][2] ),
    .B2(_06288_),
    .X(_02998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10272_ (.A1(_06222_),
    .A2(_06287_),
    .B1(\design_top.core0.REG2[4][1] ),
    .B2(_06288_),
    .X(_02997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10273_ (.A1(_06223_),
    .A2(_06274_),
    .B1(\design_top.core0.REG2[4][0] ),
    .B2(_06277_),
    .X(_02996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10274_ (.A(_05234_),
    .B(_06049_),
    .Y(_00555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10275_ (.A(_05237_),
    .B(_00555_),
    .X(_06289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10276_ (.A(_06289_),
    .X(_06290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10277_ (.A(_06289_),
    .Y(_06291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10278_ (.A(_06291_),
    .X(_06292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10279_ (.A1(_00284_),
    .A2(_06290_),
    .B1(\design_top.MEM[7][7] ),
    .B2(_06292_),
    .X(_02995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10280_ (.A1(_00283_),
    .A2(_06290_),
    .B1(\design_top.MEM[7][6] ),
    .B2(_06292_),
    .X(_02994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10281_ (.A1(_00282_),
    .A2(_06290_),
    .B1(\design_top.MEM[7][5] ),
    .B2(_06292_),
    .X(_02993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10282_ (.A1(_00281_),
    .A2(_06290_),
    .B1(\design_top.MEM[7][4] ),
    .B2(_06292_),
    .X(_02992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10283_ (.A1(_00280_),
    .A2(_06290_),
    .B1(\design_top.MEM[7][3] ),
    .B2(_06292_),
    .X(_02991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10284_ (.A1(_00279_),
    .A2(_06289_),
    .B1(\design_top.MEM[7][2] ),
    .B2(_06291_),
    .X(_02990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10285_ (.A1(_00278_),
    .A2(_06289_),
    .B1(\design_top.MEM[7][1] ),
    .B2(_06291_),
    .X(_02989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10286_ (.A1(_00277_),
    .A2(_06289_),
    .B1(\design_top.MEM[7][0] ),
    .B2(_06291_),
    .X(_02988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10287_ (.A(_05749_),
    .X(_06293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10288_ (.A(_05968_),
    .X(_06294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10289_ (.A(_06294_),
    .X(_06295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10290_ (.A(_06295_),
    .X(_06296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10291_ (.A(_06294_),
    .Y(_06297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10292_ (.A(_06297_),
    .X(_06298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10293_ (.A(_06298_),
    .X(_06299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10294_ (.A1(_06293_),
    .A2(_06296_),
    .B1(\design_top.core0.REG2[5][31] ),
    .B2(_06299_),
    .X(_02987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10295_ (.A(_05753_),
    .X(_06300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10296_ (.A1(_06300_),
    .A2(_06296_),
    .B1(\design_top.core0.REG2[5][30] ),
    .B2(_06299_),
    .X(_02986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10297_ (.A(_05757_),
    .X(_06301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10298_ (.A1(_06301_),
    .A2(_06296_),
    .B1(\design_top.core0.REG2[5][29] ),
    .B2(_06299_),
    .X(_02985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10299_ (.A(_05759_),
    .X(_06302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10300_ (.A1(_06302_),
    .A2(_06296_),
    .B1(\design_top.core0.REG2[5][28] ),
    .B2(_06299_),
    .X(_02984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10301_ (.A(_05761_),
    .X(_06303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10302_ (.A1(_06303_),
    .A2(_06296_),
    .B1(\design_top.core0.REG2[5][27] ),
    .B2(_06299_),
    .X(_02983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10303_ (.A(_05763_),
    .X(_06304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10304_ (.A(_06295_),
    .X(_06305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10305_ (.A(_06298_),
    .X(_06306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10306_ (.A1(_06304_),
    .A2(_06305_),
    .B1(\design_top.core0.REG2[5][26] ),
    .B2(_06306_),
    .X(_02982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10307_ (.A(_05765_),
    .X(_06307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10308_ (.A1(_06307_),
    .A2(_06305_),
    .B1(\design_top.core0.REG2[5][25] ),
    .B2(_06306_),
    .X(_02981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10309_ (.A(_05769_),
    .X(_06308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10310_ (.A1(_06308_),
    .A2(_06305_),
    .B1(\design_top.core0.REG2[5][24] ),
    .B2(_06306_),
    .X(_02980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10311_ (.A(_05771_),
    .X(_06309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10312_ (.A1(_06309_),
    .A2(_06305_),
    .B1(\design_top.core0.REG2[5][23] ),
    .B2(_06306_),
    .X(_02979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10313_ (.A(_05773_),
    .X(_06310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10314_ (.A1(_06310_),
    .A2(_06305_),
    .B1(\design_top.core0.REG2[5][22] ),
    .B2(_06306_),
    .X(_02978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10315_ (.A(_05775_),
    .X(_06311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10316_ (.A(_06295_),
    .X(_06312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10317_ (.A(_06298_),
    .X(_06313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10318_ (.A1(_06311_),
    .A2(_06312_),
    .B1(\design_top.core0.REG2[5][21] ),
    .B2(_06313_),
    .X(_02977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10319_ (.A(_05777_),
    .X(_06314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10320_ (.A1(_06314_),
    .A2(_06312_),
    .B1(\design_top.core0.REG2[5][20] ),
    .B2(_06313_),
    .X(_02976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10321_ (.A(_05781_),
    .X(_06315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10322_ (.A1(_06315_),
    .A2(_06312_),
    .B1(\design_top.core0.REG2[5][19] ),
    .B2(_06313_),
    .X(_02975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10323_ (.A(_05783_),
    .X(_06316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10324_ (.A1(_06316_),
    .A2(_06312_),
    .B1(\design_top.core0.REG2[5][18] ),
    .B2(_06313_),
    .X(_02974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10325_ (.A(_05785_),
    .X(_06317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10326_ (.A1(_06317_),
    .A2(_06312_),
    .B1(\design_top.core0.REG2[5][17] ),
    .B2(_06313_),
    .X(_02973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10327_ (.A(_05787_),
    .X(_06318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10328_ (.A(_06294_),
    .X(_06319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10329_ (.A(_06297_),
    .X(_06320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10330_ (.A1(_06318_),
    .A2(_06319_),
    .B1(\design_top.core0.REG2[5][16] ),
    .B2(_06320_),
    .X(_02972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10331_ (.A(_05789_),
    .X(_06321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10332_ (.A1(_06321_),
    .A2(_06319_),
    .B1(\design_top.core0.REG2[5][15] ),
    .B2(_06320_),
    .X(_02971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10333_ (.A(_05793_),
    .X(_06322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10334_ (.A1(_06322_),
    .A2(_06319_),
    .B1(\design_top.core0.REG2[5][14] ),
    .B2(_06320_),
    .X(_02970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10335_ (.A1(\design_top.core0.REG2[5][13] ),
    .A2(_06295_),
    .B1(_06268_),
    .B2(_06298_),
    .X(_02969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10336_ (.A(_05795_),
    .X(_06323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10337_ (.A1(_06323_),
    .A2(_06319_),
    .B1(\design_top.core0.REG2[5][12] ),
    .B2(_06320_),
    .X(_02968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10338_ (.A(_05797_),
    .X(_06324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10339_ (.A1(_06324_),
    .A2(_06319_),
    .B1(\design_top.core0.REG2[5][11] ),
    .B2(_06320_),
    .X(_02967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10340_ (.A(_05799_),
    .X(_06325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10341_ (.A(_06294_),
    .X(_06326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10342_ (.A(_06297_),
    .X(_06327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10343_ (.A1(_06325_),
    .A2(_06326_),
    .B1(\design_top.core0.REG2[5][10] ),
    .B2(_06327_),
    .X(_02966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10344_ (.A(_05801_),
    .X(_06328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10345_ (.A1(_06328_),
    .A2(_06326_),
    .B1(\design_top.core0.REG2[5][9] ),
    .B2(_06327_),
    .X(_02965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10346_ (.A(_05805_),
    .X(_06329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10347_ (.A1(_06329_),
    .A2(_06326_),
    .B1(\design_top.core0.REG2[5][8] ),
    .B2(_06327_),
    .X(_02964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10348_ (.A(_05807_),
    .X(_06330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10349_ (.A1(_06330_),
    .A2(_06326_),
    .B1(\design_top.core0.REG2[5][7] ),
    .B2(_06327_),
    .X(_02963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10350_ (.A(_05809_),
    .X(_06331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10351_ (.A1(_06331_),
    .A2(_06326_),
    .B1(\design_top.core0.REG2[5][6] ),
    .B2(_06327_),
    .X(_02962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10352_ (.A(_05811_),
    .X(_06332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10353_ (.A(_06294_),
    .X(_06333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10354_ (.A(_06297_),
    .X(_06334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10355_ (.A1(_06332_),
    .A2(_06333_),
    .B1(\design_top.core0.REG2[5][5] ),
    .B2(_06334_),
    .X(_02961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10356_ (.A(_05813_),
    .X(_06335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10357_ (.A1(_06335_),
    .A2(_06333_),
    .B1(\design_top.core0.REG2[5][4] ),
    .B2(_06334_),
    .X(_02960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10358_ (.A(_05817_),
    .X(_06336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10359_ (.A1(_06336_),
    .A2(_06333_),
    .B1(\design_top.core0.REG2[5][3] ),
    .B2(_06334_),
    .X(_02959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10360_ (.A(_05819_),
    .X(_06337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10361_ (.A1(_06337_),
    .A2(_06333_),
    .B1(\design_top.core0.REG2[5][2] ),
    .B2(_06334_),
    .X(_02958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10362_ (.A(_05821_),
    .X(_06338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10363_ (.A1(_06338_),
    .A2(_06333_),
    .B1(\design_top.core0.REG2[5][1] ),
    .B2(_06334_),
    .X(_02957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10364_ (.A(_05823_),
    .X(_06339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10365_ (.A1(_06339_),
    .A2(_06295_),
    .B1(\design_top.core0.REG2[5][0] ),
    .B2(_06298_),
    .X(_02956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10366_ (.A(_06015_),
    .X(_06340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10367_ (.A(_06340_),
    .X(_06341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10368_ (.A(_06341_),
    .X(_06342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10369_ (.A(_06340_),
    .Y(_06343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10370_ (.A(_06343_),
    .X(_06344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10371_ (.A(_06344_),
    .X(_06345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10372_ (.A1(_06293_),
    .A2(_06342_),
    .B1(\design_top.core0.REG2[6][31] ),
    .B2(_06345_),
    .X(_02955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10373_ (.A1(_06300_),
    .A2(_06342_),
    .B1(\design_top.core0.REG2[6][30] ),
    .B2(_06345_),
    .X(_02954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10374_ (.A1(_06301_),
    .A2(_06342_),
    .B1(\design_top.core0.REG2[6][29] ),
    .B2(_06345_),
    .X(_02953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10375_ (.A1(_06302_),
    .A2(_06342_),
    .B1(\design_top.core0.REG2[6][28] ),
    .B2(_06345_),
    .X(_02952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10376_ (.A1(_06303_),
    .A2(_06342_),
    .B1(\design_top.core0.REG2[6][27] ),
    .B2(_06345_),
    .X(_02951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10377_ (.A(_06341_),
    .X(_06346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10378_ (.A(_06344_),
    .X(_06347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10379_ (.A1(_06304_),
    .A2(_06346_),
    .B1(\design_top.core0.REG2[6][26] ),
    .B2(_06347_),
    .X(_02950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10380_ (.A1(_06307_),
    .A2(_06346_),
    .B1(\design_top.core0.REG2[6][25] ),
    .B2(_06347_),
    .X(_02949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10381_ (.A1(_06308_),
    .A2(_06346_),
    .B1(\design_top.core0.REG2[6][24] ),
    .B2(_06347_),
    .X(_02948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10382_ (.A1(_06309_),
    .A2(_06346_),
    .B1(\design_top.core0.REG2[6][23] ),
    .B2(_06347_),
    .X(_02947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10383_ (.A1(_06310_),
    .A2(_06346_),
    .B1(\design_top.core0.REG2[6][22] ),
    .B2(_06347_),
    .X(_02946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10384_ (.A(_06341_),
    .X(_06348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10385_ (.A(_06344_),
    .X(_06349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10386_ (.A1(_06311_),
    .A2(_06348_),
    .B1(\design_top.core0.REG2[6][21] ),
    .B2(_06349_),
    .X(_02945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10387_ (.A1(_06314_),
    .A2(_06348_),
    .B1(\design_top.core0.REG2[6][20] ),
    .B2(_06349_),
    .X(_02944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10388_ (.A1(_06315_),
    .A2(_06348_),
    .B1(\design_top.core0.REG2[6][19] ),
    .B2(_06349_),
    .X(_02943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10389_ (.A1(_06316_),
    .A2(_06348_),
    .B1(\design_top.core0.REG2[6][18] ),
    .B2(_06349_),
    .X(_02942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10390_ (.A1(_06317_),
    .A2(_06348_),
    .B1(\design_top.core0.REG2[6][17] ),
    .B2(_06349_),
    .X(_02941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10391_ (.A(_06340_),
    .X(_06350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10392_ (.A(_06343_),
    .X(_06351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10393_ (.A1(_06318_),
    .A2(_06350_),
    .B1(\design_top.core0.REG2[6][16] ),
    .B2(_06351_),
    .X(_02940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10394_ (.A1(_06321_),
    .A2(_06350_),
    .B1(\design_top.core0.REG2[6][15] ),
    .B2(_06351_),
    .X(_02939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10395_ (.A1(_06322_),
    .A2(_06350_),
    .B1(\design_top.core0.REG2[6][14] ),
    .B2(_06351_),
    .X(_02938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10396_ (.A1(\design_top.core0.REG2[6][13] ),
    .A2(_06341_),
    .B1(_06268_),
    .B2(_06344_),
    .X(_02937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10397_ (.A1(_06323_),
    .A2(_06350_),
    .B1(\design_top.core0.REG2[6][12] ),
    .B2(_06351_),
    .X(_02936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10398_ (.A1(_06324_),
    .A2(_06350_),
    .B1(\design_top.core0.REG2[6][11] ),
    .B2(_06351_),
    .X(_02935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10399_ (.A(_06340_),
    .X(_06352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10400_ (.A(_06343_),
    .X(_06353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10401_ (.A1(_06325_),
    .A2(_06352_),
    .B1(\design_top.core0.REG2[6][10] ),
    .B2(_06353_),
    .X(_02934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10402_ (.A1(_06328_),
    .A2(_06352_),
    .B1(\design_top.core0.REG2[6][9] ),
    .B2(_06353_),
    .X(_02933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10403_ (.A1(_06329_),
    .A2(_06352_),
    .B1(\design_top.core0.REG2[6][8] ),
    .B2(_06353_),
    .X(_02932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10404_ (.A1(_06330_),
    .A2(_06352_),
    .B1(\design_top.core0.REG2[6][7] ),
    .B2(_06353_),
    .X(_02931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10405_ (.A1(_06331_),
    .A2(_06352_),
    .B1(\design_top.core0.REG2[6][6] ),
    .B2(_06353_),
    .X(_02930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10406_ (.A(_06340_),
    .X(_06354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10407_ (.A(_06343_),
    .X(_06355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10408_ (.A1(_06332_),
    .A2(_06354_),
    .B1(\design_top.core0.REG2[6][5] ),
    .B2(_06355_),
    .X(_02929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10409_ (.A1(_06335_),
    .A2(_06354_),
    .B1(\design_top.core0.REG2[6][4] ),
    .B2(_06355_),
    .X(_02928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10410_ (.A1(_06336_),
    .A2(_06354_),
    .B1(\design_top.core0.REG2[6][3] ),
    .B2(_06355_),
    .X(_02927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10411_ (.A1(_06337_),
    .A2(_06354_),
    .B1(\design_top.core0.REG2[6][2] ),
    .B2(_06355_),
    .X(_02926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10412_ (.A1(_06338_),
    .A2(_06354_),
    .B1(\design_top.core0.REG2[6][1] ),
    .B2(_06355_),
    .X(_02925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10413_ (.A1(_06339_),
    .A2(_06341_),
    .B1(\design_top.core0.REG2[6][0] ),
    .B2(_06344_),
    .X(_02924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10414_ (.A(_06032_),
    .X(_06356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10415_ (.A(_06356_),
    .X(_06357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10416_ (.A(_06357_),
    .X(_06358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10417_ (.A(_06356_),
    .Y(_06359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10418_ (.A(_06359_),
    .X(_06360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10419_ (.A(_06360_),
    .X(_06361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10420_ (.A1(_06293_),
    .A2(_06358_),
    .B1(\design_top.core0.REG2[7][31] ),
    .B2(_06361_),
    .X(_02923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10421_ (.A1(_06300_),
    .A2(_06358_),
    .B1(\design_top.core0.REG2[7][30] ),
    .B2(_06361_),
    .X(_02922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10422_ (.A1(_06301_),
    .A2(_06358_),
    .B1(\design_top.core0.REG2[7][29] ),
    .B2(_06361_),
    .X(_02921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10423_ (.A1(_06302_),
    .A2(_06358_),
    .B1(\design_top.core0.REG2[7][28] ),
    .B2(_06361_),
    .X(_02920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10424_ (.A1(_06303_),
    .A2(_06358_),
    .B1(\design_top.core0.REG2[7][27] ),
    .B2(_06361_),
    .X(_02919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10425_ (.A(_06357_),
    .X(_06362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10426_ (.A(_06360_),
    .X(_06363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10427_ (.A1(_06304_),
    .A2(_06362_),
    .B1(\design_top.core0.REG2[7][26] ),
    .B2(_06363_),
    .X(_02918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10428_ (.A1(_06307_),
    .A2(_06362_),
    .B1(\design_top.core0.REG2[7][25] ),
    .B2(_06363_),
    .X(_02917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10429_ (.A1(_06308_),
    .A2(_06362_),
    .B1(\design_top.core0.REG2[7][24] ),
    .B2(_06363_),
    .X(_02916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10430_ (.A1(_06309_),
    .A2(_06362_),
    .B1(\design_top.core0.REG2[7][23] ),
    .B2(_06363_),
    .X(_02915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10431_ (.A1(_06310_),
    .A2(_06362_),
    .B1(\design_top.core0.REG2[7][22] ),
    .B2(_06363_),
    .X(_02914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10432_ (.A(_06357_),
    .X(_06364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10433_ (.A(_06360_),
    .X(_06365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10434_ (.A1(_06311_),
    .A2(_06364_),
    .B1(\design_top.core0.REG2[7][21] ),
    .B2(_06365_),
    .X(_02913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10435_ (.A1(_06314_),
    .A2(_06364_),
    .B1(\design_top.core0.REG2[7][20] ),
    .B2(_06365_),
    .X(_02912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10436_ (.A1(_06315_),
    .A2(_06364_),
    .B1(\design_top.core0.REG2[7][19] ),
    .B2(_06365_),
    .X(_02911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10437_ (.A1(_06316_),
    .A2(_06364_),
    .B1(\design_top.core0.REG2[7][18] ),
    .B2(_06365_),
    .X(_02910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10438_ (.A1(_06317_),
    .A2(_06364_),
    .B1(\design_top.core0.REG2[7][17] ),
    .B2(_06365_),
    .X(_02909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10439_ (.A(_06356_),
    .X(_06366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10440_ (.A(_06359_),
    .X(_06367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10441_ (.A1(_06318_),
    .A2(_06366_),
    .B1(\design_top.core0.REG2[7][16] ),
    .B2(_06367_),
    .X(_02908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10442_ (.A1(_06321_),
    .A2(_06366_),
    .B1(\design_top.core0.REG2[7][15] ),
    .B2(_06367_),
    .X(_02907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10443_ (.A1(_06322_),
    .A2(_06366_),
    .B1(\design_top.core0.REG2[7][14] ),
    .B2(_06367_),
    .X(_02906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10444_ (.A1(\design_top.core0.REG2[7][13] ),
    .A2(_06357_),
    .B1(_06268_),
    .B2(_06360_),
    .X(_02905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10445_ (.A1(_06323_),
    .A2(_06366_),
    .B1(\design_top.core0.REG2[7][12] ),
    .B2(_06367_),
    .X(_02904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10446_ (.A1(_06324_),
    .A2(_06366_),
    .B1(\design_top.core0.REG2[7][11] ),
    .B2(_06367_),
    .X(_02903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10447_ (.A(_06356_),
    .X(_06368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10448_ (.A(_06359_),
    .X(_06369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10449_ (.A1(_06325_),
    .A2(_06368_),
    .B1(\design_top.core0.REG2[7][10] ),
    .B2(_06369_),
    .X(_02902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10450_ (.A1(_06328_),
    .A2(_06368_),
    .B1(\design_top.core0.REG2[7][9] ),
    .B2(_06369_),
    .X(_02901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10451_ (.A1(_06329_),
    .A2(_06368_),
    .B1(\design_top.core0.REG2[7][8] ),
    .B2(_06369_),
    .X(_02900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10452_ (.A1(_06330_),
    .A2(_06368_),
    .B1(\design_top.core0.REG2[7][7] ),
    .B2(_06369_),
    .X(_02899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10453_ (.A1(_06331_),
    .A2(_06368_),
    .B1(\design_top.core0.REG2[7][6] ),
    .B2(_06369_),
    .X(_02898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10454_ (.A(_06356_),
    .X(_06370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10455_ (.A(_06359_),
    .X(_06371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10456_ (.A1(_06332_),
    .A2(_06370_),
    .B1(\design_top.core0.REG2[7][5] ),
    .B2(_06371_),
    .X(_02897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10457_ (.A1(_06335_),
    .A2(_06370_),
    .B1(\design_top.core0.REG2[7][4] ),
    .B2(_06371_),
    .X(_02896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10458_ (.A1(_06336_),
    .A2(_06370_),
    .B1(\design_top.core0.REG2[7][3] ),
    .B2(_06371_),
    .X(_02895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10459_ (.A1(_06337_),
    .A2(_06370_),
    .B1(\design_top.core0.REG2[7][2] ),
    .B2(_06371_),
    .X(_02894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10460_ (.A1(_06338_),
    .A2(_06370_),
    .B1(\design_top.core0.REG2[7][1] ),
    .B2(_06371_),
    .X(_02893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10461_ (.A1(_06339_),
    .A2(_06357_),
    .B1(\design_top.core0.REG2[7][0] ),
    .B2(_06360_),
    .X(_02892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10462_ (.A(_06055_),
    .X(_06372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10463_ (.A(_06372_),
    .X(_06373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10464_ (.A(_06373_),
    .X(_06374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10465_ (.A(_06372_),
    .Y(_06375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10466_ (.A(_06375_),
    .X(_06376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10467_ (.A(_06376_),
    .X(_06377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10468_ (.A1(_06293_),
    .A2(_06374_),
    .B1(\design_top.core0.REG2[8][31] ),
    .B2(_06377_),
    .X(_02891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10469_ (.A1(_06300_),
    .A2(_06374_),
    .B1(\design_top.core0.REG2[8][30] ),
    .B2(_06377_),
    .X(_02890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10470_ (.A1(_06301_),
    .A2(_06374_),
    .B1(\design_top.core0.REG2[8][29] ),
    .B2(_06377_),
    .X(_02889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10471_ (.A1(_06302_),
    .A2(_06374_),
    .B1(\design_top.core0.REG2[8][28] ),
    .B2(_06377_),
    .X(_02888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10472_ (.A1(_06303_),
    .A2(_06374_),
    .B1(\design_top.core0.REG2[8][27] ),
    .B2(_06377_),
    .X(_02887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10473_ (.A(_06373_),
    .X(_06378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10474_ (.A(_06376_),
    .X(_06379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10475_ (.A1(_06304_),
    .A2(_06378_),
    .B1(\design_top.core0.REG2[8][26] ),
    .B2(_06379_),
    .X(_02886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10476_ (.A1(_06307_),
    .A2(_06378_),
    .B1(\design_top.core0.REG2[8][25] ),
    .B2(_06379_),
    .X(_02885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10477_ (.A1(_06308_),
    .A2(_06378_),
    .B1(\design_top.core0.REG2[8][24] ),
    .B2(_06379_),
    .X(_02884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10478_ (.A1(_06309_),
    .A2(_06378_),
    .B1(\design_top.core0.REG2[8][23] ),
    .B2(_06379_),
    .X(_02883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10479_ (.A1(_06310_),
    .A2(_06378_),
    .B1(\design_top.core0.REG2[8][22] ),
    .B2(_06379_),
    .X(_02882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10480_ (.A(_06373_),
    .X(_06380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10481_ (.A(_06376_),
    .X(_06381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10482_ (.A1(_06311_),
    .A2(_06380_),
    .B1(\design_top.core0.REG2[8][21] ),
    .B2(_06381_),
    .X(_02881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10483_ (.A1(_06314_),
    .A2(_06380_),
    .B1(\design_top.core0.REG2[8][20] ),
    .B2(_06381_),
    .X(_02880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10484_ (.A1(_06315_),
    .A2(_06380_),
    .B1(\design_top.core0.REG2[8][19] ),
    .B2(_06381_),
    .X(_02879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10485_ (.A1(_06316_),
    .A2(_06380_),
    .B1(\design_top.core0.REG2[8][18] ),
    .B2(_06381_),
    .X(_02878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10486_ (.A1(_06317_),
    .A2(_06380_),
    .B1(\design_top.core0.REG2[8][17] ),
    .B2(_06381_),
    .X(_02877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10487_ (.A(_06372_),
    .X(_06382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10488_ (.A(_06375_),
    .X(_06383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10489_ (.A1(_06318_),
    .A2(_06382_),
    .B1(\design_top.core0.REG2[8][16] ),
    .B2(_06383_),
    .X(_02876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10490_ (.A1(_06321_),
    .A2(_06382_),
    .B1(\design_top.core0.REG2[8][15] ),
    .B2(_06383_),
    .X(_02875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10491_ (.A1(_06322_),
    .A2(_06382_),
    .B1(\design_top.core0.REG2[8][14] ),
    .B2(_06383_),
    .X(_02874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10492_ (.A(_05655_),
    .X(_06384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10493_ (.A1(\design_top.core0.REG2[8][13] ),
    .A2(_06373_),
    .B1(_06384_),
    .B2(_06376_),
    .X(_02873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10494_ (.A1(_06323_),
    .A2(_06382_),
    .B1(\design_top.core0.REG2[8][12] ),
    .B2(_06383_),
    .X(_02872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10495_ (.A1(_06324_),
    .A2(_06382_),
    .B1(\design_top.core0.REG2[8][11] ),
    .B2(_06383_),
    .X(_02871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10496_ (.A(_06372_),
    .X(_06385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10497_ (.A(_06375_),
    .X(_06386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10498_ (.A1(_06325_),
    .A2(_06385_),
    .B1(\design_top.core0.REG2[8][10] ),
    .B2(_06386_),
    .X(_02870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10499_ (.A1(_06328_),
    .A2(_06385_),
    .B1(\design_top.core0.REG2[8][9] ),
    .B2(_06386_),
    .X(_02869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10500_ (.A1(_06329_),
    .A2(_06385_),
    .B1(\design_top.core0.REG2[8][8] ),
    .B2(_06386_),
    .X(_02868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10501_ (.A1(_06330_),
    .A2(_06385_),
    .B1(\design_top.core0.REG2[8][7] ),
    .B2(_06386_),
    .X(_02867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10502_ (.A1(_06331_),
    .A2(_06385_),
    .B1(\design_top.core0.REG2[8][6] ),
    .B2(_06386_),
    .X(_02866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10503_ (.A(_06372_),
    .X(_06387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10504_ (.A(_06375_),
    .X(_06388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10505_ (.A1(_06332_),
    .A2(_06387_),
    .B1(\design_top.core0.REG2[8][5] ),
    .B2(_06388_),
    .X(_02865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10506_ (.A1(_06335_),
    .A2(_06387_),
    .B1(\design_top.core0.REG2[8][4] ),
    .B2(_06388_),
    .X(_02864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10507_ (.A1(_06336_),
    .A2(_06387_),
    .B1(\design_top.core0.REG2[8][3] ),
    .B2(_06388_),
    .X(_02863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10508_ (.A1(_06337_),
    .A2(_06387_),
    .B1(\design_top.core0.REG2[8][2] ),
    .B2(_06388_),
    .X(_02862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10509_ (.A1(_06338_),
    .A2(_06387_),
    .B1(\design_top.core0.REG2[8][1] ),
    .B2(_06388_),
    .X(_02861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10510_ (.A1(_06339_),
    .A2(_06373_),
    .B1(\design_top.core0.REG2[8][0] ),
    .B2(_06376_),
    .X(_02860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10511_ (.A(_06073_),
    .X(_06389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10512_ (.A(_06389_),
    .X(_06390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10513_ (.A(\design_top.core0.REG2[0][31] ),
    .B(_06390_),
    .X(_02859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10514_ (.A(\design_top.core0.REG2[0][30] ),
    .B(_06390_),
    .X(_02858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10515_ (.A(\design_top.core0.REG2[0][29] ),
    .B(_06390_),
    .X(_02857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10516_ (.A(\design_top.core0.REG2[0][28] ),
    .B(_06390_),
    .X(_02856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10517_ (.A(\design_top.core0.REG2[0][27] ),
    .B(_06390_),
    .X(_02855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10518_ (.A(_06389_),
    .X(_06391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10519_ (.A(\design_top.core0.REG2[0][26] ),
    .B(_06391_),
    .X(_02854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10520_ (.A(\design_top.core0.REG2[0][25] ),
    .B(_06391_),
    .X(_02853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10521_ (.A(\design_top.core0.REG2[0][24] ),
    .B(_06391_),
    .X(_02852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10522_ (.A(\design_top.core0.REG2[0][23] ),
    .B(_06391_),
    .X(_02851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10523_ (.A(\design_top.core0.REG2[0][22] ),
    .B(_06391_),
    .X(_02850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10524_ (.A(_06389_),
    .X(_06392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10525_ (.A(\design_top.core0.REG2[0][21] ),
    .B(_06392_),
    .X(_02849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10526_ (.A(\design_top.core0.REG2[0][20] ),
    .B(_06392_),
    .X(_02848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10527_ (.A(\design_top.core0.REG2[0][19] ),
    .B(_06392_),
    .X(_02847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10528_ (.A(\design_top.core0.REG2[0][18] ),
    .B(_06392_),
    .X(_02846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10529_ (.A(\design_top.core0.REG2[0][17] ),
    .B(_06392_),
    .X(_02845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10530_ (.A(_06073_),
    .X(_06393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10531_ (.A(\design_top.core0.REG2[0][16] ),
    .B(_06393_),
    .X(_02844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10532_ (.A(\design_top.core0.REG2[0][15] ),
    .B(_06393_),
    .X(_02843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10533_ (.A(\design_top.core0.REG2[0][14] ),
    .B(_06393_),
    .X(_02842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10534_ (.A1(\design_top.core0.REG2[0][13] ),
    .A2(_06389_),
    .B1(_06384_),
    .B2(_05604_),
    .X(_02841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10535_ (.A(\design_top.core0.REG2[0][12] ),
    .B(_06393_),
    .X(_02840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10536_ (.A(\design_top.core0.REG2[0][11] ),
    .B(_06393_),
    .X(_02839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10537_ (.A(_06073_),
    .X(_06394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10538_ (.A(\design_top.core0.REG2[0][10] ),
    .B(_06394_),
    .X(_02838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10539_ (.A(\design_top.core0.REG2[0][9] ),
    .B(_06394_),
    .X(_02837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10540_ (.A(\design_top.core0.REG2[0][8] ),
    .B(_06394_),
    .X(_02836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10541_ (.A(\design_top.core0.REG2[0][7] ),
    .B(_06394_),
    .X(_02835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10542_ (.A(\design_top.core0.REG2[0][6] ),
    .B(_06394_),
    .X(_02834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10543_ (.A(_06073_),
    .X(_06395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10544_ (.A(\design_top.core0.REG2[0][5] ),
    .B(_06395_),
    .X(_02833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10545_ (.A(\design_top.core0.REG2[0][4] ),
    .B(_06395_),
    .X(_02832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10546_ (.A(\design_top.core0.REG2[0][3] ),
    .B(_06395_),
    .X(_02831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10547_ (.A(\design_top.core0.REG2[0][2] ),
    .B(_06395_),
    .X(_02830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10548_ (.A(\design_top.core0.REG2[0][1] ),
    .B(_06395_),
    .X(_02829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10549_ (.A(\design_top.core0.REG2[0][0] ),
    .B(_06389_),
    .X(_02828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10550_ (.A(_06083_),
    .X(_06396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10551_ (.A(_06396_),
    .X(_06397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10552_ (.A(_06397_),
    .X(_06398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10553_ (.A(_06396_),
    .Y(_06399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10554_ (.A(_06399_),
    .X(_06400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10555_ (.A(_06400_),
    .X(_06401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10556_ (.A1(_06293_),
    .A2(_06398_),
    .B1(\design_top.core0.REG2[10][31] ),
    .B2(_06401_),
    .X(_02827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10557_ (.A1(_06300_),
    .A2(_06398_),
    .B1(\design_top.core0.REG2[10][30] ),
    .B2(_06401_),
    .X(_02826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10558_ (.A1(_06301_),
    .A2(_06398_),
    .B1(\design_top.core0.REG2[10][29] ),
    .B2(_06401_),
    .X(_02825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10559_ (.A1(_06302_),
    .A2(_06398_),
    .B1(\design_top.core0.REG2[10][28] ),
    .B2(_06401_),
    .X(_02824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10560_ (.A1(_06303_),
    .A2(_06398_),
    .B1(\design_top.core0.REG2[10][27] ),
    .B2(_06401_),
    .X(_02823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10561_ (.A(_06397_),
    .X(_06402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10562_ (.A(_06400_),
    .X(_06403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10563_ (.A1(_06304_),
    .A2(_06402_),
    .B1(\design_top.core0.REG2[10][26] ),
    .B2(_06403_),
    .X(_02822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10564_ (.A1(_06307_),
    .A2(_06402_),
    .B1(\design_top.core0.REG2[10][25] ),
    .B2(_06403_),
    .X(_02821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10565_ (.A1(_06308_),
    .A2(_06402_),
    .B1(\design_top.core0.REG2[10][24] ),
    .B2(_06403_),
    .X(_02820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10566_ (.A1(_06309_),
    .A2(_06402_),
    .B1(\design_top.core0.REG2[10][23] ),
    .B2(_06403_),
    .X(_02819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10567_ (.A1(_06310_),
    .A2(_06402_),
    .B1(\design_top.core0.REG2[10][22] ),
    .B2(_06403_),
    .X(_02818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10568_ (.A(_06397_),
    .X(_06404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10569_ (.A(_06400_),
    .X(_06405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10570_ (.A1(_06311_),
    .A2(_06404_),
    .B1(\design_top.core0.REG2[10][21] ),
    .B2(_06405_),
    .X(_02817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10571_ (.A1(_06314_),
    .A2(_06404_),
    .B1(\design_top.core0.REG2[10][20] ),
    .B2(_06405_),
    .X(_02816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10572_ (.A1(_06315_),
    .A2(_06404_),
    .B1(\design_top.core0.REG2[10][19] ),
    .B2(_06405_),
    .X(_02815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10573_ (.A1(_06316_),
    .A2(_06404_),
    .B1(\design_top.core0.REG2[10][18] ),
    .B2(_06405_),
    .X(_02814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10574_ (.A1(_06317_),
    .A2(_06404_),
    .B1(\design_top.core0.REG2[10][17] ),
    .B2(_06405_),
    .X(_02813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10575_ (.A(_06396_),
    .X(_06406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10576_ (.A(_06399_),
    .X(_06407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10577_ (.A1(_06318_),
    .A2(_06406_),
    .B1(\design_top.core0.REG2[10][16] ),
    .B2(_06407_),
    .X(_02812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10578_ (.A1(_06321_),
    .A2(_06406_),
    .B1(\design_top.core0.REG2[10][15] ),
    .B2(_06407_),
    .X(_02811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10579_ (.A1(_06322_),
    .A2(_06406_),
    .B1(\design_top.core0.REG2[10][14] ),
    .B2(_06407_),
    .X(_02810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10580_ (.A1(\design_top.core0.REG2[10][13] ),
    .A2(_06397_),
    .B1(_06384_),
    .B2(_06400_),
    .X(_02809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10581_ (.A1(_06323_),
    .A2(_06406_),
    .B1(\design_top.core0.REG2[10][12] ),
    .B2(_06407_),
    .X(_02808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10582_ (.A1(_06324_),
    .A2(_06406_),
    .B1(\design_top.core0.REG2[10][11] ),
    .B2(_06407_),
    .X(_02807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10583_ (.A(_06396_),
    .X(_06408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10584_ (.A(_06399_),
    .X(_06409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10585_ (.A1(_06325_),
    .A2(_06408_),
    .B1(\design_top.core0.REG2[10][10] ),
    .B2(_06409_),
    .X(_02806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10586_ (.A1(_06328_),
    .A2(_06408_),
    .B1(\design_top.core0.REG2[10][9] ),
    .B2(_06409_),
    .X(_02805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10587_ (.A1(_06329_),
    .A2(_06408_),
    .B1(\design_top.core0.REG2[10][8] ),
    .B2(_06409_),
    .X(_02804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10588_ (.A1(_06330_),
    .A2(_06408_),
    .B1(\design_top.core0.REG2[10][7] ),
    .B2(_06409_),
    .X(_02803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10589_ (.A1(_06331_),
    .A2(_06408_),
    .B1(\design_top.core0.REG2[10][6] ),
    .B2(_06409_),
    .X(_02802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10590_ (.A(_06396_),
    .X(_06410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10591_ (.A(_06399_),
    .X(_06411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10592_ (.A1(_06332_),
    .A2(_06410_),
    .B1(\design_top.core0.REG2[10][5] ),
    .B2(_06411_),
    .X(_02801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10593_ (.A1(_06335_),
    .A2(_06410_),
    .B1(\design_top.core0.REG2[10][4] ),
    .B2(_06411_),
    .X(_02800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10594_ (.A1(_06336_),
    .A2(_06410_),
    .B1(\design_top.core0.REG2[10][3] ),
    .B2(_06411_),
    .X(_02799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10595_ (.A1(_06337_),
    .A2(_06410_),
    .B1(\design_top.core0.REG2[10][2] ),
    .B2(_06411_),
    .X(_02798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10596_ (.A1(_06338_),
    .A2(_06410_),
    .B1(\design_top.core0.REG2[10][1] ),
    .B2(_06411_),
    .X(_02797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10597_ (.A1(_06339_),
    .A2(_06397_),
    .B1(\design_top.core0.REG2[10][0] ),
    .B2(_06400_),
    .X(_02796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10598_ (.A(_06101_),
    .X(_06412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10599_ (.A(_06412_),
    .X(_06413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10600_ (.A(_06413_),
    .X(_06414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10601_ (.A(_06412_),
    .Y(_06415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10602_ (.A(_06415_),
    .X(_06416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10603_ (.A(_06416_),
    .X(_06417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10604_ (.A1(_05609_),
    .A2(_06414_),
    .B1(\design_top.core0.REG2[11][31] ),
    .B2(_06417_),
    .X(_02795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10605_ (.A1(_05612_),
    .A2(_06414_),
    .B1(\design_top.core0.REG2[11][30] ),
    .B2(_06417_),
    .X(_02794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10606_ (.A1(_05615_),
    .A2(_06414_),
    .B1(\design_top.core0.REG2[11][29] ),
    .B2(_06417_),
    .X(_02793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10607_ (.A1(_05617_),
    .A2(_06414_),
    .B1(\design_top.core0.REG2[11][28] ),
    .B2(_06417_),
    .X(_02792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10608_ (.A1(_05619_),
    .A2(_06414_),
    .B1(\design_top.core0.REG2[11][27] ),
    .B2(_06417_),
    .X(_02791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10609_ (.A(_06413_),
    .X(_06418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10610_ (.A(_06416_),
    .X(_06419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10611_ (.A1(_05622_),
    .A2(_06418_),
    .B1(\design_top.core0.REG2[11][26] ),
    .B2(_06419_),
    .X(_02790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10612_ (.A1(_05625_),
    .A2(_06418_),
    .B1(\design_top.core0.REG2[11][25] ),
    .B2(_06419_),
    .X(_02789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10613_ (.A1(_05628_),
    .A2(_06418_),
    .B1(\design_top.core0.REG2[11][24] ),
    .B2(_06419_),
    .X(_02788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10614_ (.A1(_05630_),
    .A2(_06418_),
    .B1(\design_top.core0.REG2[11][23] ),
    .B2(_06419_),
    .X(_02787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10615_ (.A1(_05632_),
    .A2(_06418_),
    .B1(\design_top.core0.REG2[11][22] ),
    .B2(_06419_),
    .X(_02786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10616_ (.A(_06413_),
    .X(_06420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10617_ (.A(_06416_),
    .X(_06421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10618_ (.A1(_05635_),
    .A2(_06420_),
    .B1(\design_top.core0.REG2[11][21] ),
    .B2(_06421_),
    .X(_02785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10619_ (.A1(_05638_),
    .A2(_06420_),
    .B1(\design_top.core0.REG2[11][20] ),
    .B2(_06421_),
    .X(_02784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10620_ (.A1(_05641_),
    .A2(_06420_),
    .B1(\design_top.core0.REG2[11][19] ),
    .B2(_06421_),
    .X(_02783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10621_ (.A1(_05643_),
    .A2(_06420_),
    .B1(\design_top.core0.REG2[11][18] ),
    .B2(_06421_),
    .X(_02782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10622_ (.A1(_05645_),
    .A2(_06420_),
    .B1(\design_top.core0.REG2[11][17] ),
    .B2(_06421_),
    .X(_02781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10623_ (.A(_06412_),
    .X(_06422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10624_ (.A(_06415_),
    .X(_06423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10625_ (.A1(_05648_),
    .A2(_06422_),
    .B1(\design_top.core0.REG2[11][16] ),
    .B2(_06423_),
    .X(_02780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10626_ (.A1(_05651_),
    .A2(_06422_),
    .B1(\design_top.core0.REG2[11][15] ),
    .B2(_06423_),
    .X(_02779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10627_ (.A1(_05654_),
    .A2(_06422_),
    .B1(\design_top.core0.REG2[11][14] ),
    .B2(_06423_),
    .X(_02778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10628_ (.A1(\design_top.core0.REG2[11][13] ),
    .A2(_06413_),
    .B1(_06384_),
    .B2(_06416_),
    .X(_02777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10629_ (.A1(_05658_),
    .A2(_06422_),
    .B1(\design_top.core0.REG2[11][12] ),
    .B2(_06423_),
    .X(_02776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10630_ (.A1(_05660_),
    .A2(_06422_),
    .B1(\design_top.core0.REG2[11][11] ),
    .B2(_06423_),
    .X(_02775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10631_ (.A(_06412_),
    .X(_06424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10632_ (.A(_06415_),
    .X(_06425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10633_ (.A1(_05663_),
    .A2(_06424_),
    .B1(\design_top.core0.REG2[11][10] ),
    .B2(_06425_),
    .X(_02774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10634_ (.A1(_05666_),
    .A2(_06424_),
    .B1(\design_top.core0.REG2[11][9] ),
    .B2(_06425_),
    .X(_02773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10635_ (.A1(_05669_),
    .A2(_06424_),
    .B1(\design_top.core0.REG2[11][8] ),
    .B2(_06425_),
    .X(_02772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10636_ (.A1(_05671_),
    .A2(_06424_),
    .B1(\design_top.core0.REG2[11][7] ),
    .B2(_06425_),
    .X(_02771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10637_ (.A1(_05673_),
    .A2(_06424_),
    .B1(\design_top.core0.REG2[11][6] ),
    .B2(_06425_),
    .X(_02770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10638_ (.A(_06412_),
    .X(_06426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10639_ (.A(_06415_),
    .X(_06427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10640_ (.A1(_05676_),
    .A2(_06426_),
    .B1(\design_top.core0.REG2[11][5] ),
    .B2(_06427_),
    .X(_02769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10641_ (.A1(_05679_),
    .A2(_06426_),
    .B1(\design_top.core0.REG2[11][4] ),
    .B2(_06427_),
    .X(_02768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10642_ (.A1(_05682_),
    .A2(_06426_),
    .B1(\design_top.core0.REG2[11][3] ),
    .B2(_06427_),
    .X(_02767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10643_ (.A1(_05684_),
    .A2(_06426_),
    .B1(\design_top.core0.REG2[11][2] ),
    .B2(_06427_),
    .X(_02766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10644_ (.A1(_05686_),
    .A2(_06426_),
    .B1(\design_top.core0.REG2[11][1] ),
    .B2(_06427_),
    .X(_02765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10645_ (.A1(_05688_),
    .A2(_06413_),
    .B1(\design_top.core0.REG2[11][0] ),
    .B2(_06416_),
    .X(_02764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10646_ (.A(_06118_),
    .X(_06428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10647_ (.A(_06428_),
    .X(_06429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10648_ (.A(_06429_),
    .X(_06430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10649_ (.A(_06428_),
    .Y(_06431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10650_ (.A(_06431_),
    .X(_06432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10651_ (.A(_06432_),
    .X(_06433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10652_ (.A1(_05609_),
    .A2(_06430_),
    .B1(\design_top.core0.REG2[12][31] ),
    .B2(_06433_),
    .X(_02763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10653_ (.A1(_05612_),
    .A2(_06430_),
    .B1(\design_top.core0.REG2[12][30] ),
    .B2(_06433_),
    .X(_02762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10654_ (.A1(_05615_),
    .A2(_06430_),
    .B1(\design_top.core0.REG2[12][29] ),
    .B2(_06433_),
    .X(_02761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10655_ (.A1(_05617_),
    .A2(_06430_),
    .B1(\design_top.core0.REG2[12][28] ),
    .B2(_06433_),
    .X(_02760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10656_ (.A1(_05619_),
    .A2(_06430_),
    .B1(\design_top.core0.REG2[12][27] ),
    .B2(_06433_),
    .X(_02759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10657_ (.A(_06429_),
    .X(_06434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10658_ (.A(_06432_),
    .X(_06435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10659_ (.A1(_05622_),
    .A2(_06434_),
    .B1(\design_top.core0.REG2[12][26] ),
    .B2(_06435_),
    .X(_02758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10660_ (.A1(_05625_),
    .A2(_06434_),
    .B1(\design_top.core0.REG2[12][25] ),
    .B2(_06435_),
    .X(_02757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10661_ (.A1(_05628_),
    .A2(_06434_),
    .B1(\design_top.core0.REG2[12][24] ),
    .B2(_06435_),
    .X(_02756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10662_ (.A1(_05630_),
    .A2(_06434_),
    .B1(\design_top.core0.REG2[12][23] ),
    .B2(_06435_),
    .X(_02755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10663_ (.A1(_05632_),
    .A2(_06434_),
    .B1(\design_top.core0.REG2[12][22] ),
    .B2(_06435_),
    .X(_02754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10664_ (.A(_06429_),
    .X(_06436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10665_ (.A(_06432_),
    .X(_06437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10666_ (.A1(_05635_),
    .A2(_06436_),
    .B1(\design_top.core0.REG2[12][21] ),
    .B2(_06437_),
    .X(_02753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10667_ (.A1(_05638_),
    .A2(_06436_),
    .B1(\design_top.core0.REG2[12][20] ),
    .B2(_06437_),
    .X(_02752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10668_ (.A1(_05641_),
    .A2(_06436_),
    .B1(\design_top.core0.REG2[12][19] ),
    .B2(_06437_),
    .X(_02751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10669_ (.A1(_05643_),
    .A2(_06436_),
    .B1(\design_top.core0.REG2[12][18] ),
    .B2(_06437_),
    .X(_02750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10670_ (.A1(_05645_),
    .A2(_06436_),
    .B1(\design_top.core0.REG2[12][17] ),
    .B2(_06437_),
    .X(_02749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10671_ (.A(_06428_),
    .X(_06438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10672_ (.A(_06431_),
    .X(_06439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10673_ (.A1(_05648_),
    .A2(_06438_),
    .B1(\design_top.core0.REG2[12][16] ),
    .B2(_06439_),
    .X(_02748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10674_ (.A1(_05651_),
    .A2(_06438_),
    .B1(\design_top.core0.REG2[12][15] ),
    .B2(_06439_),
    .X(_02747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10675_ (.A1(_05654_),
    .A2(_06438_),
    .B1(\design_top.core0.REG2[12][14] ),
    .B2(_06439_),
    .X(_02746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10676_ (.A1(\design_top.core0.REG2[12][13] ),
    .A2(_06429_),
    .B1(_06384_),
    .B2(_06432_),
    .X(_02745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10677_ (.A1(_05658_),
    .A2(_06438_),
    .B1(\design_top.core0.REG2[12][12] ),
    .B2(_06439_),
    .X(_02744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10678_ (.A1(_05660_),
    .A2(_06438_),
    .B1(\design_top.core0.REG2[12][11] ),
    .B2(_06439_),
    .X(_02743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10679_ (.A(_06428_),
    .X(_06440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10680_ (.A(_06431_),
    .X(_06441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10681_ (.A1(_05663_),
    .A2(_06440_),
    .B1(\design_top.core0.REG2[12][10] ),
    .B2(_06441_),
    .X(_02742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10682_ (.A1(_05666_),
    .A2(_06440_),
    .B1(\design_top.core0.REG2[12][9] ),
    .B2(_06441_),
    .X(_02741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10683_ (.A1(_05669_),
    .A2(_06440_),
    .B1(\design_top.core0.REG2[12][8] ),
    .B2(_06441_),
    .X(_02740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10684_ (.A1(_05671_),
    .A2(_06440_),
    .B1(\design_top.core0.REG2[12][7] ),
    .B2(_06441_),
    .X(_02739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10685_ (.A1(_05673_),
    .A2(_06440_),
    .B1(\design_top.core0.REG2[12][6] ),
    .B2(_06441_),
    .X(_02738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10686_ (.A(_06428_),
    .X(_06442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10687_ (.A(_06431_),
    .X(_06443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10688_ (.A1(_05676_),
    .A2(_06442_),
    .B1(\design_top.core0.REG2[12][5] ),
    .B2(_06443_),
    .X(_02737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10689_ (.A1(_05679_),
    .A2(_06442_),
    .B1(\design_top.core0.REG2[12][4] ),
    .B2(_06443_),
    .X(_02736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10690_ (.A1(_05682_),
    .A2(_06442_),
    .B1(\design_top.core0.REG2[12][3] ),
    .B2(_06443_),
    .X(_02735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10691_ (.A1(_05684_),
    .A2(_06442_),
    .B1(\design_top.core0.REG2[12][2] ),
    .B2(_06443_),
    .X(_02734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10692_ (.A1(_05686_),
    .A2(_06442_),
    .B1(\design_top.core0.REG2[12][1] ),
    .B2(_06443_),
    .X(_02733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10693_ (.A1(_05688_),
    .A2(_06429_),
    .B1(\design_top.core0.REG2[12][0] ),
    .B2(_06432_),
    .X(_02732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10694_ (.A(_06135_),
    .X(_06444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10695_ (.A(_06444_),
    .X(_06445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10696_ (.A(_06445_),
    .X(_06446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10697_ (.A(_06444_),
    .Y(_06447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10698_ (.A(_06447_),
    .X(_06448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10699_ (.A(_06448_),
    .X(_06449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10700_ (.A1(_05609_),
    .A2(_06446_),
    .B1(\design_top.core0.REG2[13][31] ),
    .B2(_06449_),
    .X(_02731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10701_ (.A1(_05612_),
    .A2(_06446_),
    .B1(\design_top.core0.REG2[13][30] ),
    .B2(_06449_),
    .X(_02730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10702_ (.A1(_05615_),
    .A2(_06446_),
    .B1(\design_top.core0.REG2[13][29] ),
    .B2(_06449_),
    .X(_02729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10703_ (.A1(_05617_),
    .A2(_06446_),
    .B1(\design_top.core0.REG2[13][28] ),
    .B2(_06449_),
    .X(_02728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10704_ (.A1(_05619_),
    .A2(_06446_),
    .B1(\design_top.core0.REG2[13][27] ),
    .B2(_06449_),
    .X(_02727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10705_ (.A(_06445_),
    .X(_06450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10706_ (.A(_06448_),
    .X(_06451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10707_ (.A1(_05622_),
    .A2(_06450_),
    .B1(\design_top.core0.REG2[13][26] ),
    .B2(_06451_),
    .X(_02726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10708_ (.A1(_05625_),
    .A2(_06450_),
    .B1(\design_top.core0.REG2[13][25] ),
    .B2(_06451_),
    .X(_02725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10709_ (.A1(_05628_),
    .A2(_06450_),
    .B1(\design_top.core0.REG2[13][24] ),
    .B2(_06451_),
    .X(_02724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10710_ (.A1(_05630_),
    .A2(_06450_),
    .B1(\design_top.core0.REG2[13][23] ),
    .B2(_06451_),
    .X(_02723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10711_ (.A1(_05632_),
    .A2(_06450_),
    .B1(\design_top.core0.REG2[13][22] ),
    .B2(_06451_),
    .X(_02722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10712_ (.A(_06445_),
    .X(_06452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10713_ (.A(_06448_),
    .X(_06453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10714_ (.A1(_05635_),
    .A2(_06452_),
    .B1(\design_top.core0.REG2[13][21] ),
    .B2(_06453_),
    .X(_02721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10715_ (.A1(_05638_),
    .A2(_06452_),
    .B1(\design_top.core0.REG2[13][20] ),
    .B2(_06453_),
    .X(_02720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10716_ (.A1(_05641_),
    .A2(_06452_),
    .B1(\design_top.core0.REG2[13][19] ),
    .B2(_06453_),
    .X(_02719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10717_ (.A1(_05643_),
    .A2(_06452_),
    .B1(\design_top.core0.REG2[13][18] ),
    .B2(_06453_),
    .X(_02718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10718_ (.A1(_05645_),
    .A2(_06452_),
    .B1(\design_top.core0.REG2[13][17] ),
    .B2(_06453_),
    .X(_02717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10719_ (.A(_06444_),
    .X(_06454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10720_ (.A(_06447_),
    .X(_06455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10721_ (.A1(_05648_),
    .A2(_06454_),
    .B1(\design_top.core0.REG2[13][16] ),
    .B2(_06455_),
    .X(_02716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10722_ (.A1(_05651_),
    .A2(_06454_),
    .B1(\design_top.core0.REG2[13][15] ),
    .B2(_06455_),
    .X(_02715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10723_ (.A1(_05654_),
    .A2(_06454_),
    .B1(\design_top.core0.REG2[13][14] ),
    .B2(_06455_),
    .X(_02714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10724_ (.A1(\design_top.core0.REG2[13][13] ),
    .A2(_06445_),
    .B1(_05876_),
    .B2(_06448_),
    .X(_02713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10725_ (.A1(_05658_),
    .A2(_06454_),
    .B1(\design_top.core0.REG2[13][12] ),
    .B2(_06455_),
    .X(_02712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10726_ (.A1(_05660_),
    .A2(_06454_),
    .B1(\design_top.core0.REG2[13][11] ),
    .B2(_06455_),
    .X(_02711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10727_ (.A(_06444_),
    .X(_06456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10728_ (.A(_06447_),
    .X(_06457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10729_ (.A1(_05663_),
    .A2(_06456_),
    .B1(\design_top.core0.REG2[13][10] ),
    .B2(_06457_),
    .X(_02710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10730_ (.A1(_05666_),
    .A2(_06456_),
    .B1(\design_top.core0.REG2[13][9] ),
    .B2(_06457_),
    .X(_02709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10731_ (.A1(_05669_),
    .A2(_06456_),
    .B1(\design_top.core0.REG2[13][8] ),
    .B2(_06457_),
    .X(_02708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10732_ (.A1(_05671_),
    .A2(_06456_),
    .B1(\design_top.core0.REG2[13][7] ),
    .B2(_06457_),
    .X(_02707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10733_ (.A1(_05673_),
    .A2(_06456_),
    .B1(\design_top.core0.REG2[13][6] ),
    .B2(_06457_),
    .X(_02706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10734_ (.A(_06444_),
    .X(_06458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10735_ (.A(_06447_),
    .X(_06459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10736_ (.A1(_05676_),
    .A2(_06458_),
    .B1(\design_top.core0.REG2[13][5] ),
    .B2(_06459_),
    .X(_02705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10737_ (.A1(_05679_),
    .A2(_06458_),
    .B1(\design_top.core0.REG2[13][4] ),
    .B2(_06459_),
    .X(_02704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10738_ (.A1(_05682_),
    .A2(_06458_),
    .B1(\design_top.core0.REG2[13][3] ),
    .B2(_06459_),
    .X(_02703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10739_ (.A1(_05684_),
    .A2(_06458_),
    .B1(\design_top.core0.REG2[13][2] ),
    .B2(_06459_),
    .X(_02702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10740_ (.A1(_05686_),
    .A2(_06458_),
    .B1(\design_top.core0.REG2[13][1] ),
    .B2(_06459_),
    .X(_02701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10741_ (.A1(_05688_),
    .A2(_06445_),
    .B1(\design_top.core0.REG2[13][0] ),
    .B2(_06448_),
    .X(_02700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10742_ (.A(_06152_),
    .X(_06460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10743_ (.A(_06460_),
    .X(_06461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10744_ (.A(_06461_),
    .X(_06462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10745_ (.A(_06460_),
    .Y(_06463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10746_ (.A(_06463_),
    .X(_06464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10747_ (.A(_06464_),
    .X(_06465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10748_ (.A1(_05609_),
    .A2(_06462_),
    .B1(\design_top.core0.REG2[14][31] ),
    .B2(_06465_),
    .X(_02699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10749_ (.A1(_05612_),
    .A2(_06462_),
    .B1(\design_top.core0.REG2[14][30] ),
    .B2(_06465_),
    .X(_02698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10750_ (.A1(_05615_),
    .A2(_06462_),
    .B1(\design_top.core0.REG2[14][29] ),
    .B2(_06465_),
    .X(_02697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10751_ (.A1(_05617_),
    .A2(_06462_),
    .B1(\design_top.core0.REG2[14][28] ),
    .B2(_06465_),
    .X(_02696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10752_ (.A1(_05619_),
    .A2(_06462_),
    .B1(\design_top.core0.REG2[14][27] ),
    .B2(_06465_),
    .X(_02695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10753_ (.A(_06461_),
    .X(_06466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10754_ (.A(_06464_),
    .X(_06467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10755_ (.A1(_05622_),
    .A2(_06466_),
    .B1(\design_top.core0.REG2[14][26] ),
    .B2(_06467_),
    .X(_02694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10756_ (.A1(_05625_),
    .A2(_06466_),
    .B1(\design_top.core0.REG2[14][25] ),
    .B2(_06467_),
    .X(_02693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10757_ (.A1(_05628_),
    .A2(_06466_),
    .B1(\design_top.core0.REG2[14][24] ),
    .B2(_06467_),
    .X(_02692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10758_ (.A1(_05630_),
    .A2(_06466_),
    .B1(\design_top.core0.REG2[14][23] ),
    .B2(_06467_),
    .X(_02691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10759_ (.A1(_05632_),
    .A2(_06466_),
    .B1(\design_top.core0.REG2[14][22] ),
    .B2(_06467_),
    .X(_02690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10760_ (.A(_06461_),
    .X(_06468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10761_ (.A(_06464_),
    .X(_06469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10762_ (.A1(_05635_),
    .A2(_06468_),
    .B1(\design_top.core0.REG2[14][21] ),
    .B2(_06469_),
    .X(_02689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10763_ (.A1(_05638_),
    .A2(_06468_),
    .B1(\design_top.core0.REG2[14][20] ),
    .B2(_06469_),
    .X(_02688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10764_ (.A1(_05641_),
    .A2(_06468_),
    .B1(\design_top.core0.REG2[14][19] ),
    .B2(_06469_),
    .X(_02687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10765_ (.A1(_05643_),
    .A2(_06468_),
    .B1(\design_top.core0.REG2[14][18] ),
    .B2(_06469_),
    .X(_02686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10766_ (.A1(_05645_),
    .A2(_06468_),
    .B1(\design_top.core0.REG2[14][17] ),
    .B2(_06469_),
    .X(_02685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10767_ (.A(_06460_),
    .X(_06470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10768_ (.A(_06463_),
    .X(_06471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10769_ (.A1(_05648_),
    .A2(_06470_),
    .B1(\design_top.core0.REG2[14][16] ),
    .B2(_06471_),
    .X(_02684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10770_ (.A1(_05651_),
    .A2(_06470_),
    .B1(\design_top.core0.REG2[14][15] ),
    .B2(_06471_),
    .X(_02683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10771_ (.A1(_05654_),
    .A2(_06470_),
    .B1(\design_top.core0.REG2[14][14] ),
    .B2(_06471_),
    .X(_02682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10772_ (.A1(\design_top.core0.REG2[14][13] ),
    .A2(_06461_),
    .B1(_05876_),
    .B2(_06464_),
    .X(_02681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10773_ (.A1(_05658_),
    .A2(_06470_),
    .B1(\design_top.core0.REG2[14][12] ),
    .B2(_06471_),
    .X(_02680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10774_ (.A1(_05660_),
    .A2(_06470_),
    .B1(\design_top.core0.REG2[14][11] ),
    .B2(_06471_),
    .X(_02679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10775_ (.A(_06460_),
    .X(_06472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10776_ (.A(_06463_),
    .X(_06473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10777_ (.A1(_05663_),
    .A2(_06472_),
    .B1(\design_top.core0.REG2[14][10] ),
    .B2(_06473_),
    .X(_02678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10778_ (.A1(_05666_),
    .A2(_06472_),
    .B1(\design_top.core0.REG2[14][9] ),
    .B2(_06473_),
    .X(_02677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10779_ (.A1(_05669_),
    .A2(_06472_),
    .B1(\design_top.core0.REG2[14][8] ),
    .B2(_06473_),
    .X(_02676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10780_ (.A1(_05671_),
    .A2(_06472_),
    .B1(\design_top.core0.REG2[14][7] ),
    .B2(_06473_),
    .X(_02675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10781_ (.A1(_05673_),
    .A2(_06472_),
    .B1(\design_top.core0.REG2[14][6] ),
    .B2(_06473_),
    .X(_02674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10782_ (.A(_06460_),
    .X(_06474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10783_ (.A(_06463_),
    .X(_06475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10784_ (.A1(_05676_),
    .A2(_06474_),
    .B1(\design_top.core0.REG2[14][5] ),
    .B2(_06475_),
    .X(_02673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10785_ (.A1(_05679_),
    .A2(_06474_),
    .B1(\design_top.core0.REG2[14][4] ),
    .B2(_06475_),
    .X(_02672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10786_ (.A1(_05682_),
    .A2(_06474_),
    .B1(\design_top.core0.REG2[14][3] ),
    .B2(_06475_),
    .X(_02671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10787_ (.A1(_05684_),
    .A2(_06474_),
    .B1(\design_top.core0.REG2[14][2] ),
    .B2(_06475_),
    .X(_02670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10788_ (.A1(_05686_),
    .A2(_06474_),
    .B1(\design_top.core0.REG2[14][1] ),
    .B2(_06475_),
    .X(_02669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10789_ (.A1(_05688_),
    .A2(_06461_),
    .B1(\design_top.core0.REG2[14][0] ),
    .B2(_06464_),
    .X(_02668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10790_ (.A(_05248_),
    .B(_06049_),
    .Y(_00554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10791_ (.A(_05251_),
    .B(_00554_),
    .X(_06476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10792_ (.A(_06476_),
    .X(_06477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10793_ (.A(_06476_),
    .Y(_06478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10794_ (.A(_06478_),
    .X(_06479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10795_ (.A1(_00292_),
    .A2(_06477_),
    .B1(\design_top.MEM[8][7] ),
    .B2(_06479_),
    .X(_02667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10796_ (.A1(_00291_),
    .A2(_06477_),
    .B1(\design_top.MEM[8][6] ),
    .B2(_06479_),
    .X(_02666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10797_ (.A1(_00290_),
    .A2(_06477_),
    .B1(\design_top.MEM[8][5] ),
    .B2(_06479_),
    .X(_02665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10798_ (.A1(_00289_),
    .A2(_06477_),
    .B1(\design_top.MEM[8][4] ),
    .B2(_06479_),
    .X(_02664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10799_ (.A1(_00288_),
    .A2(_06477_),
    .B1(\design_top.MEM[8][3] ),
    .B2(_06479_),
    .X(_02663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10800_ (.A1(_00287_),
    .A2(_06476_),
    .B1(\design_top.MEM[8][2] ),
    .B2(_06478_),
    .X(_02662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10801_ (.A1(_00286_),
    .A2(_06476_),
    .B1(\design_top.MEM[8][1] ),
    .B2(_06478_),
    .X(_02661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10802_ (.A1(_00285_),
    .A2(_06476_),
    .B1(\design_top.MEM[8][0] ),
    .B2(_06478_),
    .X(_02660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10803_ (.A(_04876_),
    .B(_05689_),
    .Y(_00550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10804_ (.A(_04886_),
    .B(_00550_),
    .X(_06480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10805_ (.A(_06480_),
    .X(_06481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10806_ (.A(_06480_),
    .Y(_06482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10807_ (.A(_06482_),
    .X(_06483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10808_ (.A1(_00300_),
    .A2(_06481_),
    .B1(\design_top.MEM[9][7] ),
    .B2(_06483_),
    .X(_02659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10809_ (.A1(_00299_),
    .A2(_06481_),
    .B1(\design_top.MEM[9][6] ),
    .B2(_06483_),
    .X(_02658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10810_ (.A1(_00298_),
    .A2(_06481_),
    .B1(\design_top.MEM[9][5] ),
    .B2(_06483_),
    .X(_02657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10811_ (.A1(_00297_),
    .A2(_06481_),
    .B1(\design_top.MEM[9][4] ),
    .B2(_06483_),
    .X(_02656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10812_ (.A1(_00296_),
    .A2(_06481_),
    .B1(\design_top.MEM[9][3] ),
    .B2(_06483_),
    .X(_02655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10813_ (.A1(_00295_),
    .A2(_06480_),
    .B1(\design_top.MEM[9][2] ),
    .B2(_06482_),
    .X(_02654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10814_ (.A1(_00294_),
    .A2(_06480_),
    .B1(\design_top.MEM[9][1] ),
    .B2(_06482_),
    .X(_02653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10815_ (.A1(_00293_),
    .A2(_06480_),
    .B1(\design_top.MEM[9][0] ),
    .B2(_06482_),
    .X(_02652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10816_ (.A(_05274_),
    .Y(_06484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10817_ (.A(_05014_),
    .B(_06484_),
    .X(_06485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10818_ (.A(_04906_),
    .B(_05018_),
    .X(_06486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10819_ (.A(_06485_),
    .B(_06486_),
    .X(_06487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10820_ (.A(_06487_),
    .X(_06488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10821_ (.A(_06487_),
    .Y(_06489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10822_ (.A(_06489_),
    .X(_06490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10823_ (.A1(\design_top.GPIOFF[15] ),
    .A2(_06488_),
    .B1(\design_top.DATAO[31] ),
    .B2(_06490_),
    .X(_02651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10824_ (.A1(\design_top.GPIOFF[14] ),
    .A2(_06488_),
    .B1(\design_top.DATAO[30] ),
    .B2(_06490_),
    .X(_02650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10825_ (.A1(\design_top.GPIOFF[13] ),
    .A2(_06488_),
    .B1(\design_top.DATAO[29] ),
    .B2(_06490_),
    .X(_02649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10826_ (.A1(\design_top.GPIOFF[12] ),
    .A2(_06488_),
    .B1(\design_top.DATAO[28] ),
    .B2(_06490_),
    .X(_02648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10827_ (.A1(\design_top.GPIOFF[11] ),
    .A2(_06488_),
    .B1(\design_top.DATAO[27] ),
    .B2(_06490_),
    .X(_02647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10828_ (.A(_06487_),
    .X(_06491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10829_ (.A(_06489_),
    .X(_06492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10830_ (.A1(\design_top.GPIOFF[10] ),
    .A2(_06491_),
    .B1(\design_top.DATAO[26] ),
    .B2(_06492_),
    .X(_02646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10831_ (.A1(\design_top.GPIOFF[9] ),
    .A2(_06491_),
    .B1(\design_top.DATAO[25] ),
    .B2(_06492_),
    .X(_02645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10832_ (.A1(\design_top.GPIOFF[8] ),
    .A2(_06491_),
    .B1(\design_top.DATAO[24] ),
    .B2(_06492_),
    .X(_02644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10833_ (.A1(\design_top.GPIOFF[7] ),
    .A2(_06491_),
    .B1(\design_top.DATAO[23] ),
    .B2(_06492_),
    .X(_02643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10834_ (.A1(\design_top.GPIOFF[6] ),
    .A2(_06491_),
    .B1(\design_top.DATAO[22] ),
    .B2(_06492_),
    .X(_02642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10835_ (.A(_06487_),
    .X(_06493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10836_ (.A(_06489_),
    .X(_06494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10837_ (.A1(\design_top.GPIOFF[5] ),
    .A2(_06493_),
    .B1(\design_top.DATAO[21] ),
    .B2(_06494_),
    .X(_02641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10838_ (.A1(\design_top.GPIOFF[4] ),
    .A2(_06493_),
    .B1(\design_top.DATAO[20] ),
    .B2(_06494_),
    .X(_02640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10839_ (.A1(\design_top.GPIOFF[3] ),
    .A2(_06493_),
    .B1(\design_top.DATAO[19] ),
    .B2(_06494_),
    .X(_02639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10840_ (.A1(\design_top.GPIOFF[2] ),
    .A2(_06493_),
    .B1(\design_top.DATAO[18] ),
    .B2(_06494_),
    .X(_02638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10841_ (.A1(\design_top.GPIOFF[1] ),
    .A2(_06493_),
    .B1(\design_top.DATAO[17] ),
    .B2(_06494_),
    .X(_02637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10842_ (.A1(io_out[15]),
    .A2(_06487_),
    .B1(\design_top.DATAO[16] ),
    .B2(_06489_),
    .X(_02636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10843_ (.A(_00548_),
    .B(_06486_),
    .X(_06495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10844_ (.A(_06495_),
    .X(_06496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10845_ (.A(_06495_),
    .Y(_06497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10846_ (.A(_06497_),
    .X(_06498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10847_ (.A1(\design_top.LEDFF[15] ),
    .A2(_06496_),
    .B1(\design_top.DATAO[15] ),
    .B2(_06498_),
    .X(_02635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10848_ (.A1(\design_top.LEDFF[14] ),
    .A2(_06496_),
    .B1(\design_top.DATAO[14] ),
    .B2(_06498_),
    .X(_02634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10849_ (.A1(\design_top.LEDFF[13] ),
    .A2(_06496_),
    .B1(\design_top.DATAO[13] ),
    .B2(_06498_),
    .X(_02633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10850_ (.A1(\design_top.LEDFF[12] ),
    .A2(_06496_),
    .B1(\design_top.DATAO[12] ),
    .B2(_06498_),
    .X(_02632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10851_ (.A1(\design_top.LEDFF[11] ),
    .A2(_06496_),
    .B1(\design_top.DATAO[11] ),
    .B2(_06498_),
    .X(_02631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10852_ (.A(_06495_),
    .X(_06499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10853_ (.A(_06497_),
    .X(_06500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10854_ (.A1(\design_top.LEDFF[10] ),
    .A2(_06499_),
    .B1(\design_top.DATAO[10] ),
    .B2(_06500_),
    .X(_02630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10855_ (.A1(\design_top.LEDFF[9] ),
    .A2(_06499_),
    .B1(\design_top.DATAO[9] ),
    .B2(_06500_),
    .X(_02629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10856_ (.A1(\design_top.LEDFF[8] ),
    .A2(_06499_),
    .B1(\design_top.DATAO[8] ),
    .B2(_06500_),
    .X(_02628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10857_ (.A1(\design_top.LEDFF[7] ),
    .A2(_06499_),
    .B1(\design_top.DATAO[7] ),
    .B2(_06500_),
    .X(_02627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10858_ (.A1(\design_top.LEDFF[6] ),
    .A2(_06499_),
    .B1(\design_top.DATAO[6] ),
    .B2(_06500_),
    .X(_02626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10859_ (.A(_06495_),
    .X(_06501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10860_ (.A(_06497_),
    .X(_06502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10861_ (.A1(\design_top.LEDFF[5] ),
    .A2(_06501_),
    .B1(\design_top.DATAO[5] ),
    .B2(_06502_),
    .X(_02625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10862_ (.A1(\design_top.LEDFF[4] ),
    .A2(_06501_),
    .B1(\design_top.DATAO[4] ),
    .B2(_06502_),
    .X(_02624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10863_ (.A1(io_out[11]),
    .A2(_06501_),
    .B1(\design_top.DATAO[3] ),
    .B2(_06502_),
    .X(_02623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10864_ (.A1(io_out[10]),
    .A2(_06501_),
    .B1(\design_top.DATAO[2] ),
    .B2(_06502_),
    .X(_02622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10865_ (.A1(io_out[9]),
    .A2(_06501_),
    .B1(\design_top.DATAO[1] ),
    .B2(_06502_),
    .X(_02621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10866_ (.A1(io_out[8]),
    .A2(_06495_),
    .B1(\design_top.DATAO[0] ),
    .B2(_06497_),
    .X(_02620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10867_ (.A1(\design_top.ROMFF2[31] ),
    .A2(_05470_),
    .B1(\design_top.ROMFF[31] ),
    .B2(\design_top.HLT ),
    .X(_02619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10868_ (.A1(\design_top.ROMFF2[30] ),
    .A2(_05470_),
    .B1(\design_top.ROMFF[30] ),
    .B2(\design_top.HLT ),
    .X(_02618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10869_ (.A1(\design_top.ROMFF2[29] ),
    .A2(_05470_),
    .B1(\design_top.ROMFF[29] ),
    .B2(\design_top.HLT ),
    .X(_02617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10870_ (.A(_05419_),
    .X(_06503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10871_ (.A1(\design_top.ROMFF2[28] ),
    .A2(_05470_),
    .B1(\design_top.ROMFF[28] ),
    .B2(_06503_),
    .X(_02616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10872_ (.A(_05424_),
    .X(_06504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10873_ (.A1(\design_top.ROMFF2[27] ),
    .A2(_06504_),
    .B1(\design_top.ROMFF[27] ),
    .B2(_06503_),
    .X(_02615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10874_ (.A1(\design_top.ROMFF2[26] ),
    .A2(_06504_),
    .B1(\design_top.ROMFF[26] ),
    .B2(_06503_),
    .X(_02614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10875_ (.A1(\design_top.ROMFF2[25] ),
    .A2(_06504_),
    .B1(\design_top.ROMFF[25] ),
    .B2(_06503_),
    .X(_02613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10876_ (.A1(\design_top.ROMFF2[24] ),
    .A2(_06504_),
    .B1(\design_top.ROMFF[24] ),
    .B2(_06503_),
    .X(_02612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10877_ (.A(_05318_),
    .X(_06505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10878_ (.A(_06505_),
    .X(_06506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10879_ (.A1(\design_top.ROMFF2[23] ),
    .A2(_06504_),
    .B1(\design_top.ROMFF[23] ),
    .B2(_06506_),
    .X(_02611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10880_ (.A(_05383_),
    .X(_06507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10881_ (.A(_06507_),
    .X(_06508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10882_ (.A1(\design_top.ROMFF2[22] ),
    .A2(_06508_),
    .B1(\design_top.ROMFF[22] ),
    .B2(_06506_),
    .X(_02610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10883_ (.A1(\design_top.ROMFF2[21] ),
    .A2(_06508_),
    .B1(\design_top.ROMFF[21] ),
    .B2(_06506_),
    .X(_02609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10884_ (.A1(\design_top.ROMFF2[20] ),
    .A2(_06508_),
    .B1(\design_top.ROMFF[20] ),
    .B2(_06506_),
    .X(_02608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10885_ (.A1(\design_top.ROMFF2[19] ),
    .A2(_06508_),
    .B1(\design_top.ROMFF[19] ),
    .B2(_06506_),
    .X(_02607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10886_ (.A(_06505_),
    .X(_06509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10887_ (.A1(\design_top.ROMFF2[18] ),
    .A2(_06508_),
    .B1(\design_top.ROMFF[18] ),
    .B2(_06509_),
    .X(_02606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10888_ (.A(_06507_),
    .X(_06510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10889_ (.A1(\design_top.ROMFF2[17] ),
    .A2(_06510_),
    .B1(\design_top.ROMFF[17] ),
    .B2(_06509_),
    .X(_02605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10890_ (.A1(\design_top.ROMFF2[16] ),
    .A2(_06510_),
    .B1(\design_top.ROMFF[16] ),
    .B2(_06509_),
    .X(_02604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10891_ (.A1(\design_top.ROMFF2[15] ),
    .A2(_06510_),
    .B1(\design_top.ROMFF[15] ),
    .B2(_06509_),
    .X(_02603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10892_ (.A1(\design_top.ROMFF2[14] ),
    .A2(_06510_),
    .B1(\design_top.ROMFF[14] ),
    .B2(_06509_),
    .X(_02602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10893_ (.A(_06505_),
    .X(_06511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10894_ (.A1(\design_top.ROMFF2[13] ),
    .A2(_06510_),
    .B1(\design_top.ROMFF[13] ),
    .B2(_06511_),
    .X(_02601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10895_ (.A(_06507_),
    .X(_06512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10896_ (.A1(\design_top.ROMFF2[12] ),
    .A2(_06512_),
    .B1(\design_top.ROMFF[12] ),
    .B2(_06511_),
    .X(_02600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10897_ (.A1(\design_top.ROMFF2[11] ),
    .A2(_06512_),
    .B1(\design_top.ROMFF[11] ),
    .B2(_06511_),
    .X(_02599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10898_ (.A1(\design_top.ROMFF2[10] ),
    .A2(_06512_),
    .B1(\design_top.ROMFF[10] ),
    .B2(_06511_),
    .X(_02598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10899_ (.A1(\design_top.ROMFF2[9] ),
    .A2(_06512_),
    .B1(\design_top.ROMFF[9] ),
    .B2(_06511_),
    .X(_02597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10900_ (.A(_06505_),
    .X(_06513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10901_ (.A1(\design_top.ROMFF2[8] ),
    .A2(_06512_),
    .B1(\design_top.ROMFF[8] ),
    .B2(_06513_),
    .X(_02596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10902_ (.A(_06507_),
    .X(_06514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10903_ (.A1(\design_top.ROMFF2[7] ),
    .A2(_06514_),
    .B1(\design_top.ROMFF[7] ),
    .B2(_06513_),
    .X(_02595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10904_ (.A1(\design_top.ROMFF2[6] ),
    .A2(_06514_),
    .B1(\design_top.ROMFF[6] ),
    .B2(_06513_),
    .X(_02594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10905_ (.A1(\design_top.ROMFF2[5] ),
    .A2(_06514_),
    .B1(\design_top.ROMFF[5] ),
    .B2(_06513_),
    .X(_02593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10906_ (.A1(\design_top.ROMFF2[4] ),
    .A2(_06514_),
    .B1(\design_top.ROMFF[4] ),
    .B2(_06513_),
    .X(_02592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10907_ (.A(_06505_),
    .X(_06515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10908_ (.A1(\design_top.ROMFF2[3] ),
    .A2(_06514_),
    .B1(\design_top.ROMFF[3] ),
    .B2(_06515_),
    .X(_02591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10909_ (.A(_06507_),
    .X(_06516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10910_ (.A1(\design_top.ROMFF2[2] ),
    .A2(_06516_),
    .B1(\design_top.ROMFF[2] ),
    .B2(_06515_),
    .X(_02590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10911_ (.A1(\design_top.ROMFF2[1] ),
    .A2(_06516_),
    .B1(\design_top.ROMFF[1] ),
    .B2(_06515_),
    .X(_02589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10912_ (.A1(\design_top.ROMFF2[0] ),
    .A2(_06516_),
    .B1(\design_top.ROMFF[0] ),
    .B2(_06515_),
    .X(_02588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10913_ (.A1(\design_top.uart0.UART_XREQ ),
    .A2(_05538_),
    .B1(\design_top.uart0.UART_XACK ),
    .B2(_05546_),
    .X(_02587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10914_ (.A(\design_top.uart0.UART_RACK ),
    .Y(_06517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _10915_ (.A0(_06517_),
    .A1(\design_top.uart0.UART_RREQ ),
    .S(_05554_),
    .X(_02586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10916_ (.A(\design_top.uart0.UART_RXDFF[2] ),
    .X(_06518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _10917_ (.A(_05562_),
    .B(_05561_),
    .C(_05552_),
    .D(_05548_),
    .X(_06519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _10918_ (.A0(_06518_),
    .A1(\design_top.uart0.UART_RFIFO[7] ),
    .S(_06519_),
    .X(_02585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _10919_ (.A(_05562_),
    .B(_05564_),
    .C(_05552_),
    .D(_05485_),
    .X(_06520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _10920_ (.A0(_06518_),
    .A1(\design_top.uart0.UART_RFIFO[6] ),
    .S(_06520_),
    .X(_02584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10921_ (.A(_05551_),
    .X(_06521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _10922_ (.A(_05553_),
    .B(_05561_),
    .C(_06521_),
    .D(_05485_),
    .X(_06522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _10923_ (.A0(_06518_),
    .A1(\design_top.uart0.UART_RFIFO[5] ),
    .S(_06522_),
    .X(_02583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _10924_ (.A(_05552_),
    .B(_05548_),
    .C(_05553_),
    .D(_05564_),
    .X(_06523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _10925_ (.A0(_06518_),
    .A1(\design_top.uart0.UART_RFIFO[4] ),
    .S(_06523_),
    .X(_02582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _10926_ (.A(_05562_),
    .B(_05561_),
    .C(_06521_),
    .D(_05558_),
    .X(_06524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _10927_ (.A0(\design_top.uart0.UART_RXDFF[2] ),
    .A1(\design_top.uart0.UART_RFIFO[3] ),
    .S(_06524_),
    .X(_02581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _10928_ (.A(_05562_),
    .B(_05564_),
    .C(_06521_),
    .D(_05558_),
    .X(_06525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _10929_ (.A0(\design_top.uart0.UART_RXDFF[2] ),
    .A1(\design_top.uart0.UART_RFIFO[2] ),
    .S(_06525_),
    .X(_02580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _10930_ (.A(_05553_),
    .B(_05549_),
    .C(_06521_),
    .D(_05558_),
    .X(_06526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _10931_ (.A0(\design_top.uart0.UART_RXDFF[2] ),
    .A1(\design_top.uart0.UART_RFIFO[1] ),
    .S(_06526_),
    .X(_02579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _10932_ (.A(_05553_),
    .B(_05564_),
    .C(_06521_),
    .D(_05558_),
    .X(_06527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _10933_ (.A0(\design_top.uart0.UART_RXDFF[2] ),
    .A1(\design_top.uart0.UART_RFIFO[0] ),
    .S(_06527_),
    .X(_02578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10934_ (.A1(\design_top.core0.NXPC[31] ),
    .A2(_06516_),
    .B1(\design_top.core0.PC[31] ),
    .B2(_06515_),
    .X(_02577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10935_ (.A(_05318_),
    .X(_06528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10936_ (.A(_06528_),
    .X(_06529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10937_ (.A1(\design_top.core0.NXPC[30] ),
    .A2(_06516_),
    .B1(\design_top.core0.PC[30] ),
    .B2(_06529_),
    .X(_02576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10938_ (.A(_05383_),
    .X(_06530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10939_ (.A(_06530_),
    .X(_06531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10940_ (.A1(\design_top.core0.NXPC[29] ),
    .A2(_06531_),
    .B1(\design_top.core0.PC[29] ),
    .B2(_06529_),
    .X(_02575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10941_ (.A1(\design_top.core0.NXPC[28] ),
    .A2(_06531_),
    .B1(\design_top.core0.PC[28] ),
    .B2(_06529_),
    .X(_02574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10942_ (.A1(\design_top.core0.NXPC[27] ),
    .A2(_06531_),
    .B1(\design_top.core0.PC[27] ),
    .B2(_06529_),
    .X(_02573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10943_ (.A1(\design_top.core0.NXPC[26] ),
    .A2(_06531_),
    .B1(\design_top.core0.PC[26] ),
    .B2(_06529_),
    .X(_02572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10944_ (.A(_06528_),
    .X(_06532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10945_ (.A1(\design_top.core0.NXPC[25] ),
    .A2(_06531_),
    .B1(\design_top.core0.PC[25] ),
    .B2(_06532_),
    .X(_02571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10946_ (.A(_06530_),
    .X(_06533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10947_ (.A1(\design_top.core0.NXPC[24] ),
    .A2(_06533_),
    .B1(\design_top.core0.PC[24] ),
    .B2(_06532_),
    .X(_02570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10948_ (.A1(\design_top.core0.NXPC[23] ),
    .A2(_06533_),
    .B1(\design_top.core0.PC[23] ),
    .B2(_06532_),
    .X(_02569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10949_ (.A1(\design_top.core0.NXPC[22] ),
    .A2(_06533_),
    .B1(\design_top.core0.PC[22] ),
    .B2(_06532_),
    .X(_02568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10950_ (.A1(\design_top.core0.NXPC[21] ),
    .A2(_06533_),
    .B1(\design_top.core0.PC[21] ),
    .B2(_06532_),
    .X(_02567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10951_ (.A(_06528_),
    .X(_06534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10952_ (.A1(\design_top.core0.NXPC[20] ),
    .A2(_06533_),
    .B1(\design_top.core0.PC[20] ),
    .B2(_06534_),
    .X(_02566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10953_ (.A(_06530_),
    .X(_06535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10954_ (.A1(\design_top.core0.NXPC[19] ),
    .A2(_06535_),
    .B1(\design_top.core0.PC[19] ),
    .B2(_06534_),
    .X(_02565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10955_ (.A1(\design_top.core0.NXPC[18] ),
    .A2(_06535_),
    .B1(\design_top.core0.PC[18] ),
    .B2(_06534_),
    .X(_02564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10956_ (.A1(\design_top.core0.NXPC[17] ),
    .A2(_06535_),
    .B1(\design_top.core0.PC[17] ),
    .B2(_06534_),
    .X(_02563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10957_ (.A1(\design_top.core0.NXPC[16] ),
    .A2(_06535_),
    .B1(\design_top.core0.PC[16] ),
    .B2(_06534_),
    .X(_02562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10958_ (.A(_06528_),
    .X(_06536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10959_ (.A1(\design_top.core0.NXPC[15] ),
    .A2(_06535_),
    .B1(\design_top.core0.PC[15] ),
    .B2(_06536_),
    .X(_02561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10960_ (.A(_06530_),
    .X(_06537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10961_ (.A1(\design_top.core0.NXPC[14] ),
    .A2(_06537_),
    .B1(\design_top.core0.PC[14] ),
    .B2(_06536_),
    .X(_02560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10962_ (.A1(\design_top.core0.NXPC[13] ),
    .A2(_06537_),
    .B1(\design_top.core0.PC[13] ),
    .B2(_06536_),
    .X(_02559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10963_ (.A1(\design_top.core0.NXPC[12] ),
    .A2(_06537_),
    .B1(\design_top.core0.PC[12] ),
    .B2(_06536_),
    .X(_02558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10964_ (.A1(\design_top.core0.NXPC[11] ),
    .A2(_06537_),
    .B1(\design_top.core0.PC[11] ),
    .B2(_06536_),
    .X(_02557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10965_ (.A(_06528_),
    .X(_06538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10966_ (.A1(\design_top.core0.NXPC[10] ),
    .A2(_06537_),
    .B1(\design_top.core0.PC[10] ),
    .B2(_06538_),
    .X(_02556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10967_ (.A(_06530_),
    .X(_06539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10968_ (.A1(\design_top.core0.NXPC[9] ),
    .A2(_06539_),
    .B1(\design_top.core0.PC[9] ),
    .B2(_06538_),
    .X(_02555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10969_ (.A1(\design_top.core0.NXPC[8] ),
    .A2(_06539_),
    .B1(\design_top.core0.PC[8] ),
    .B2(_06538_),
    .X(_02554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10970_ (.A1(\design_top.core0.NXPC[7] ),
    .A2(_06539_),
    .B1(\design_top.core0.PC[7] ),
    .B2(_06538_),
    .X(_02553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10971_ (.A1(\design_top.core0.NXPC[6] ),
    .A2(_06539_),
    .B1(\design_top.core0.PC[6] ),
    .B2(_06538_),
    .X(_02552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10972_ (.A(_05318_),
    .X(_06540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10973_ (.A(_06540_),
    .X(_06541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10974_ (.A1(\design_top.core0.NXPC[5] ),
    .A2(_06539_),
    .B1(\design_top.core0.PC[5] ),
    .B2(_06541_),
    .X(_02551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10975_ (.A(_05383_),
    .X(_06542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10976_ (.A(_06542_),
    .X(_06543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10977_ (.A1(\design_top.core0.NXPC[4] ),
    .A2(_06543_),
    .B1(\design_top.core0.PC[4] ),
    .B2(_06541_),
    .X(_02550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10978_ (.A1(\design_top.core0.NXPC[3] ),
    .A2(_06543_),
    .B1(\design_top.core0.PC[3] ),
    .B2(_06541_),
    .X(_02549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10979_ (.A1(\design_top.core0.NXPC[2] ),
    .A2(_06543_),
    .B1(\design_top.core0.PC[2] ),
    .B2(_06541_),
    .X(_02548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10980_ (.A1(\design_top.core0.NXPC[1] ),
    .A2(_06543_),
    .B1(\design_top.core0.PC[1] ),
    .B2(_06541_),
    .X(_02547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10981_ (.A(_06540_),
    .X(_06544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10982_ (.A1(\design_top.core0.NXPC[0] ),
    .A2(_06543_),
    .B1(\design_top.core0.PC[0] ),
    .B2(_06544_),
    .X(_02546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10983_ (.A(_06542_),
    .X(_06545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10984_ (.A1(\design_top.IADDR[31] ),
    .A2(_06545_),
    .B1(\design_top.core0.NXPC[31] ),
    .B2(_06544_),
    .X(_02545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10985_ (.A1(\design_top.IADDR[30] ),
    .A2(_06545_),
    .B1(\design_top.core0.NXPC[30] ),
    .B2(_06544_),
    .X(_02544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10986_ (.A1(\design_top.IADDR[29] ),
    .A2(_06545_),
    .B1(\design_top.core0.NXPC[29] ),
    .B2(_06544_),
    .X(_02543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10987_ (.A1(\design_top.IADDR[28] ),
    .A2(_06545_),
    .B1(\design_top.core0.NXPC[28] ),
    .B2(_06544_),
    .X(_02542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10988_ (.A(_06540_),
    .X(_06546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10989_ (.A1(\design_top.IADDR[27] ),
    .A2(_06545_),
    .B1(\design_top.core0.NXPC[27] ),
    .B2(_06546_),
    .X(_02541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10990_ (.A(_06542_),
    .X(_06547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10991_ (.A1(\design_top.IADDR[26] ),
    .A2(_06547_),
    .B1(\design_top.core0.NXPC[26] ),
    .B2(_06546_),
    .X(_02540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10992_ (.A1(\design_top.IADDR[25] ),
    .A2(_06547_),
    .B1(\design_top.core0.NXPC[25] ),
    .B2(_06546_),
    .X(_02539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10993_ (.A1(\design_top.IADDR[24] ),
    .A2(_06547_),
    .B1(\design_top.core0.NXPC[24] ),
    .B2(_06546_),
    .X(_02538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10994_ (.A1(\design_top.IADDR[23] ),
    .A2(_06547_),
    .B1(\design_top.core0.NXPC[23] ),
    .B2(_06546_),
    .X(_02537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10995_ (.A(_06540_),
    .X(_06548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10996_ (.A1(\design_top.IADDR[22] ),
    .A2(_06547_),
    .B1(\design_top.core0.NXPC[22] ),
    .B2(_06548_),
    .X(_02536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10997_ (.A(_06542_),
    .X(_06549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10998_ (.A1(\design_top.IADDR[21] ),
    .A2(_06549_),
    .B1(\design_top.core0.NXPC[21] ),
    .B2(_06548_),
    .X(_02535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _10999_ (.A1(\design_top.IADDR[20] ),
    .A2(_06549_),
    .B1(\design_top.core0.NXPC[20] ),
    .B2(_06548_),
    .X(_02534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11000_ (.A1(\design_top.IADDR[19] ),
    .A2(_06549_),
    .B1(\design_top.core0.NXPC[19] ),
    .B2(_06548_),
    .X(_02533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11001_ (.A1(\design_top.IADDR[18] ),
    .A2(_06549_),
    .B1(\design_top.core0.NXPC[18] ),
    .B2(_06548_),
    .X(_02532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11002_ (.A(_06540_),
    .X(_06550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11003_ (.A1(\design_top.IADDR[17] ),
    .A2(_06549_),
    .B1(\design_top.core0.NXPC[17] ),
    .B2(_06550_),
    .X(_02531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11004_ (.A(_06542_),
    .X(_06551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11005_ (.A1(\design_top.IADDR[16] ),
    .A2(_06551_),
    .B1(\design_top.core0.NXPC[16] ),
    .B2(_06550_),
    .X(_02530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11006_ (.A1(\design_top.IADDR[15] ),
    .A2(_06551_),
    .B1(\design_top.core0.NXPC[15] ),
    .B2(_06550_),
    .X(_02529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11007_ (.A1(\design_top.IADDR[14] ),
    .A2(_06551_),
    .B1(\design_top.core0.NXPC[14] ),
    .B2(_06550_),
    .X(_02528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11008_ (.A1(\design_top.IADDR[13] ),
    .A2(_06551_),
    .B1(\design_top.core0.NXPC[13] ),
    .B2(_06550_),
    .X(_02527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11009_ (.A(_05302_),
    .X(_06552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11010_ (.A1(\design_top.IADDR[12] ),
    .A2(_06551_),
    .B1(\design_top.core0.NXPC[12] ),
    .B2(_06552_),
    .X(_02526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11011_ (.A(_05384_),
    .X(_06553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11012_ (.A1(\design_top.IADDR[11] ),
    .A2(_06553_),
    .B1(\design_top.core0.NXPC[11] ),
    .B2(_06552_),
    .X(_02525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11013_ (.A1(\design_top.IADDR[10] ),
    .A2(_06553_),
    .B1(\design_top.core0.NXPC[10] ),
    .B2(_06552_),
    .X(_02524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11014_ (.A1(\design_top.IADDR[9] ),
    .A2(_06553_),
    .B1(\design_top.core0.NXPC[9] ),
    .B2(_06552_),
    .X(_02523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11015_ (.A1(\design_top.IADDR[8] ),
    .A2(_06553_),
    .B1(\design_top.core0.NXPC[8] ),
    .B2(_06552_),
    .X(_02522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11016_ (.A(_05302_),
    .X(_06554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11017_ (.A1(\design_top.IADDR[7] ),
    .A2(_06553_),
    .B1(\design_top.core0.NXPC[7] ),
    .B2(_06554_),
    .X(_02521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11018_ (.A(_05384_),
    .X(_06555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11019_ (.A1(\design_top.IADDR[6] ),
    .A2(_06555_),
    .B1(\design_top.core0.NXPC[6] ),
    .B2(_06554_),
    .X(_02520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11020_ (.A1(\design_top.IADDR[5] ),
    .A2(_06555_),
    .B1(\design_top.core0.NXPC[5] ),
    .B2(_06554_),
    .X(_02519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11021_ (.A1(_05469_),
    .A2(_06555_),
    .B1(\design_top.core0.NXPC[4] ),
    .B2(_06554_),
    .X(_02518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11022_ (.A1(io_out[19]),
    .A2(_06555_),
    .B1(\design_top.core0.NXPC[3] ),
    .B2(_06554_),
    .X(_02517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11023_ (.A1(io_out[18]),
    .A2(_06555_),
    .B1(\design_top.core0.NXPC[2] ),
    .B2(_05434_),
    .X(_02516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11024_ (.A1(io_out[17]),
    .A2(_05379_),
    .B1(\design_top.core0.NXPC[1] ),
    .B2(_05434_),
    .X(_02515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11025_ (.A1(io_out[16]),
    .A2(_05379_),
    .B1(\design_top.core0.NXPC[0] ),
    .B2(_05434_),
    .X(_02514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11026_ (.A(_04758_),
    .X(_00714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11027_ (.A(_00720_),
    .B(_04682_),
    .Y(_00721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11028_ (.A(_04842_),
    .X(_00722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11029_ (.A(_04665_),
    .B(_00723_),
    .Y(_00724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11030_ (.A(_04775_),
    .X(_06556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11031_ (.A(_06556_),
    .X(_00726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11032_ (.A(_00482_),
    .B(_00732_),
    .Y(_00733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11033_ (.A(_04782_),
    .X(_00734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11034_ (.A(_04656_),
    .B(_00740_),
    .Y(_00741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11035_ (.A(_04785_),
    .X(_06557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11036_ (.A(_06557_),
    .X(_00743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11037_ (.A(_04658_),
    .B(_00749_),
    .Y(_00750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11038_ (.A(_04630_),
    .Y(_00757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11039_ (.A(_04791_),
    .X(_00759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11040_ (.A(\design_top.core0.REG1[13][31] ),
    .Y(_00377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11041_ (.A(\design_top.core0.REG1[14][31] ),
    .Y(_00378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11042_ (.A(\design_top.core0.REG1[15][31] ),
    .Y(_00379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11043_ (.A(_00772_),
    .B(_04632_),
    .Y(_00774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11044_ (.A(\design_top.core0.REG1[8][31] ),
    .Y(_00371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11045_ (.A(\design_top.core0.REG1[9][31] ),
    .Y(_00372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11046_ (.A(\design_top.core0.REG1[10][31] ),
    .Y(_00373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11047_ (.A(\design_top.core0.REG1[11][31] ),
    .Y(_00374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11048_ (.A(\design_top.core0.REG1[12][31] ),
    .Y(_00376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11049_ (.A(_04634_),
    .B(_00781_),
    .Y(_00782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11050_ (.A(_00524_),
    .B(_00783_),
    .Y(_00785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11051_ (.A(_04808_),
    .X(_00786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11052_ (.A(\design_top.core0.REG1[2][31] ),
    .Y(_00363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11053_ (.A(\design_top.core0.REG1[3][31] ),
    .Y(_00364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11054_ (.A(\design_top.core0.REG1[4][31] ),
    .Y(_00366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11055_ (.A(\design_top.core0.REG1[5][31] ),
    .Y(_00367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11056_ (.A(\design_top.core0.REG1[6][31] ),
    .Y(_00368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11057_ (.A(\design_top.core0.REG1[7][31] ),
    .Y(_00369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11058_ (.A(_00530_),
    .B(_00792_),
    .Y(_00793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11059_ (.A(_04720_),
    .Y(io_out[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11060_ (.A(\design_top.core0.REG1[1][31] ),
    .Y(_00362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11061_ (.A(_00799_),
    .B(_04642_),
    .Y(_00801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11062_ (.A(_04802_),
    .X(_00802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11063_ (.A(_00808_),
    .X(_06558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11064_ (.A(_06558_),
    .X(_06559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11065_ (.A(_04644_),
    .B(_06559_),
    .Y(_00809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11066_ (.A(_04650_),
    .Y(_00810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11067_ (.A(_00816_),
    .B(_00342_),
    .Y(_00818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11068_ (.A1(_00316_),
    .A2(_04626_),
    .B1(_00313_),
    .B2(_00304_),
    .X(_06560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11069_ (.A(_06560_),
    .Y(_00819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11070_ (.A(_00825_),
    .X(_06561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11071_ (.A(_06561_),
    .X(_06562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11072_ (.A(_06562_),
    .B(_06560_),
    .Y(_00826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11073_ (.A(_04627_),
    .Y(_00827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11074_ (.A(_04629_),
    .Y(_00834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11075_ (.A1_N(\design_top.IACK[7] ),
    .A2_N(\design_top.IREQ[7] ),
    .B1(\design_top.IACK[7] ),
    .B2(\design_top.IREQ[7] ),
    .X(_00346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11076_ (.A(_04806_),
    .X(_01389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11077_ (.A1(_00816_),
    .A2(_04650_),
    .B1(_00818_),
    .X(_06563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11078_ (.A(_04661_),
    .B(_00819_),
    .X(_06564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11079_ (.A(_06564_),
    .X(_01655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11080_ (.A1(_00825_),
    .A2(_06560_),
    .B1(_01655_),
    .X(_06565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11081_ (.A(_00840_),
    .Y(_06566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11082_ (.A(_06566_),
    .B(_00333_),
    .Y(_06567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11083_ (.A1(_00833_),
    .A2(_00827_),
    .B1(_04628_),
    .B2(_06567_),
    .X(_06568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11084_ (.A1(_00825_),
    .A2(_00819_),
    .B1(_06565_),
    .B2(_06568_),
    .X(_06569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11085_ (.A1(_00816_),
    .A2(_00810_),
    .B1(_06563_),
    .B2(_06569_),
    .X(_06570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11086_ (.A(_04647_),
    .X(_06571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11087_ (.A(_04804_),
    .X(_01391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _11088_ (.A1(_04802_),
    .A2(_00808_),
    .A3(_04643_),
    .B1(_00799_),
    .B2(_01391_),
    .X(_06572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11089_ (.A1(_04808_),
    .A2(_00792_),
    .B1(_04641_),
    .B2(_06572_),
    .X(_06573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11090_ (.A(_06571_),
    .B(_06573_),
    .X(_06574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11091_ (.A1(_01389_),
    .A2(_00783_),
    .B1(_04648_),
    .B2(_06570_),
    .C1(_06574_),
    .X(_06575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _11092_ (.A1(_00775_),
    .A2(_00781_),
    .A3(_04633_),
    .B1(_00772_),
    .B2(_01385_),
    .X(_06576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11093_ (.A1(_04791_),
    .A2(_00765_),
    .B1(_04638_),
    .B2(_06576_),
    .X(_06577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11094_ (.A(_04631_),
    .B(_06577_),
    .X(_06578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11095_ (.A1(_00756_),
    .A2(_01383_),
    .B1(_04639_),
    .B2(_06575_),
    .C1(_06578_),
    .X(_06579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11096_ (.A(_06579_),
    .X(_06580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11097_ (.A1(_00743_),
    .A2(_00749_),
    .B1(_04660_),
    .B2(_06580_),
    .X(_06581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11098_ (.A1(_00734_),
    .A2(_00740_),
    .B1(_04657_),
    .B2(_06581_),
    .X(_06582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11099_ (.A1(_00726_),
    .A2(_00732_),
    .B1(_04654_),
    .B2(_06582_),
    .X(_06583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11100_ (.A1(_00722_),
    .A2(_00723_),
    .B1(_04666_),
    .B2(_06583_),
    .X(_06584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11101_ (.A(_00591_),
    .Y(_06585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11102_ (.A(_04722_),
    .X(_00594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11103_ (.A(_04728_),
    .X(_06586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11104_ (.A(_04863_),
    .X(_00603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _11105_ (.A1(_06586_),
    .A2(_00618_),
    .A3(_04705_),
    .B1(_00603_),
    .B2(_00609_),
    .X(_06587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11106_ (.A1(_00594_),
    .A2(_00600_),
    .B1(_04700_),
    .B2(_06587_),
    .X(_06588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11107_ (.A(_04733_),
    .X(_06589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11108_ (.A(_06589_),
    .X(_00620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11109_ (.A(_04771_),
    .X(_00654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11110_ (.A(_04849_),
    .X(_00688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11111_ (.A(_04750_),
    .X(_00697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11112_ (.A(_04756_),
    .X(_00705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _11113_ (.A1(_00720_),
    .A2(_00714_),
    .A3(_04679_),
    .B1(_00705_),
    .B2(_00711_),
    .X(_06590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11114_ (.A1(_00697_),
    .A2(_00703_),
    .B1(_04686_),
    .B2(_06590_),
    .X(_06591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11115_ (.A1(_00688_),
    .A2(_00694_),
    .B1(_04681_),
    .B2(_06591_),
    .X(_06592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11116_ (.A(_04768_),
    .X(_06593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11117_ (.A(_04761_),
    .X(_00671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _11118_ (.A1(_04764_),
    .A2(_00686_),
    .A3(_04698_),
    .B1(_00671_),
    .B2(_00677_),
    .X(_06594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11119_ (.A1(_06593_),
    .A2(_00669_),
    .B1(_04690_),
    .B2(_06594_),
    .X(_06595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11120_ (.A(_04692_),
    .B(_06595_),
    .X(_06596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11121_ (.A1(_00654_),
    .A2(_00660_),
    .B1(_04699_),
    .B2(_06592_),
    .C1(_06596_),
    .X(_06597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11122_ (.A(_04735_),
    .X(_06598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11123_ (.A(_06598_),
    .X(_00629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11124_ (.A(_04746_),
    .X(_00646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11125_ (.A(_04743_),
    .X(_00637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _11126_ (.A1(_00646_),
    .A2(_00652_),
    .A3(_04673_),
    .B1(_00637_),
    .B2(_00643_),
    .X(_06599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11127_ (.A1(_00629_),
    .A2(_00635_),
    .B1(_04671_),
    .B2(_06599_),
    .X(_06600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11128_ (.A(_04669_),
    .B(_06600_),
    .X(_06601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11129_ (.A1(_00620_),
    .A2(_00626_),
    .B1(_04676_),
    .B2(_06597_),
    .C1(_06601_),
    .X(_06602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11130_ (.A1(_04702_),
    .A2(_06588_),
    .B1(_04706_),
    .B2(_06602_),
    .X(_06603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221ai_2 _11131_ (.A1(_04707_),
    .A2(_06584_),
    .B1(_04867_),
    .B2(_06585_),
    .C1(_06603_),
    .Y(_00841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11132_ (.A(_00582_),
    .Y(_06604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11133_ (.A(_00381_),
    .B(_00582_),
    .Y(_06605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11134_ (.A1(_00722_),
    .A2(_00576_),
    .B1(_06556_),
    .B2(_00731_),
    .X(_06606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11135_ (.A(_00739_),
    .Y(_06607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11136_ (.A(_00748_),
    .Y(_06608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11137_ (.A1(_01383_),
    .A2(_00755_),
    .B1(_00759_),
    .B2(_00764_),
    .X(_06609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11138_ (.A(_00764_),
    .Y(_06610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11139_ (.A(_00771_),
    .Y(_06611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11140_ (.A(_00780_),
    .Y(_06612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11141_ (.A1(_04634_),
    .A2(_06612_),
    .B1(_04632_),
    .B2(_06611_),
    .X(_06613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a221oi_2 _11142_ (.A1(_00506_),
    .A2(_06610_),
    .B1(_04632_),
    .B2(_06611_),
    .C1(_06613_),
    .Y(_06614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11143_ (.A1(_06557_),
    .A2(_00748_),
    .B1(_01383_),
    .B2(_00755_),
    .X(_06615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11144_ (.A1(_06609_),
    .A2(_06614_),
    .B1(_06615_),
    .Y(_06616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221ai_2 _11145_ (.A1(_04656_),
    .A2(_06607_),
    .B1(_04658_),
    .B2(_06608_),
    .C1(_06616_),
    .Y(_06617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11146_ (.A1(_00734_),
    .A2(_00739_),
    .B1(_00726_),
    .B2(_00731_),
    .C1(_06617_),
    .X(_06618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11147_ (.A1(_00722_),
    .A2(_00576_),
    .B1(_06606_),
    .B2(_06618_),
    .X(_06619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11148_ (.A1(_01389_),
    .A2(_00570_),
    .B1(_00786_),
    .B2(_00791_),
    .X(_06620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11149_ (.A1(_01391_),
    .A2(_00798_),
    .B1(_00802_),
    .B2(_00807_),
    .X(_06621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11150_ (.A1(_04825_),
    .A2(_00815_),
    .B1(_04663_),
    .B2(_00824_),
    .X(_06622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11151_ (.A(_00832_),
    .Y(_06623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11152_ (.A(_00324_),
    .B(_06623_),
    .X(_06624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11153_ (.A(_06624_),
    .Y(_06625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11154_ (.A1(_04821_),
    .A2(_00832_),
    .B1(_04819_),
    .B2(_00839_),
    .C1(_06624_),
    .X(_06626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11155_ (.A1(_06625_),
    .A2(_06626_),
    .B1(_04663_),
    .B2(_00824_),
    .X(_06627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11156_ (.A(_04825_),
    .B(_00815_),
    .X(_06628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11157_ (.A1(_00802_),
    .A2(_00807_),
    .B1(_06622_),
    .B2(_06627_),
    .C1(_06628_),
    .X(_06629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11158_ (.A(_01391_),
    .B(_00798_),
    .X(_06630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11159_ (.A1(_00786_),
    .A2(_00791_),
    .B1(_06621_),
    .B2(_06629_),
    .C1(_06630_),
    .X(_06631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221ai_2 _11160_ (.A1(_00759_),
    .A2(_00764_),
    .B1(_01385_),
    .B2(_00771_),
    .C1(_06613_),
    .Y(_06632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221ai_2 _11161_ (.A1(_00734_),
    .A2(_00739_),
    .B1(_06556_),
    .B2(_00731_),
    .C1(_06615_),
    .Y(_06633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11162_ (.A(_00576_),
    .Y(_06634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a221o_2 _11163_ (.A1(_04665_),
    .A2(_06634_),
    .B1(_04634_),
    .B2(_06612_),
    .C1(_06606_),
    .X(_06635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a221o_2 _11164_ (.A1(_00734_),
    .A2(_00739_),
    .B1(_00743_),
    .B2(_00748_),
    .C1(_06609_),
    .X(_06636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11165_ (.A(_06632_),
    .B(_06633_),
    .C(_06635_),
    .D(_06636_),
    .X(_06637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11166_ (.A(_06637_),
    .Y(_06638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11167_ (.A1(_01389_),
    .A2(_00570_),
    .B1(_06620_),
    .B2(_06631_),
    .C1(_06638_),
    .X(_06639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11168_ (.A(_06619_),
    .B(_06639_),
    .Y(_06640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11169_ (.A1(_00688_),
    .A2(_00693_),
    .B1(_00697_),
    .B2(_00702_),
    .X(_06641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11170_ (.A(_00671_),
    .B(_00676_),
    .X(_06642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11171_ (.A1(_00654_),
    .A2(_00659_),
    .B1(_06642_),
    .Y(_06643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11172_ (.A1(_00719_),
    .A2(_00714_),
    .B1(_00705_),
    .B2(_00710_),
    .X(_06644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11173_ (.A1(_00671_),
    .A2(_00676_),
    .B1(_00685_),
    .B2(_04764_),
    .X(_06645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11174_ (.A1(_00654_),
    .A2(_00659_),
    .B1(_06593_),
    .B2(_00668_),
    .X(_06646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11175_ (.A1(_00697_),
    .A2(_00702_),
    .B1(_00705_),
    .B2(_00710_),
    .X(_06647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4b_2 _11176_ (.A(_06644_),
    .B(_06645_),
    .C(_06646_),
    .D_N(_06647_),
    .X(_06648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11177_ (.A(_06593_),
    .X(_00663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11178_ (.A(_04764_),
    .X(_00680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11179_ (.A1(_00719_),
    .A2(_00714_),
    .B1(_00688_),
    .B2(_00693_),
    .X(_06649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11180_ (.A1(_00663_),
    .A2(_00668_),
    .B1(_00685_),
    .B2(_00680_),
    .C1(_06649_),
    .X(_06650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4b_2 _11181_ (.A(_06641_),
    .B(_06643_),
    .C(_06648_),
    .D_N(_06650_),
    .X(_06651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _11182_ (.A1(_06644_),
    .A2(_06647_),
    .B1(_06641_),
    .X(_06652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11183_ (.A1(_00688_),
    .A2(_00693_),
    .B1(_00685_),
    .B2(_00680_),
    .C1(_06652_),
    .X(_06653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11184_ (.A1(_00663_),
    .A2(_00668_),
    .B1(_06645_),
    .B2(_06653_),
    .C1(_06642_),
    .X(_06654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _11185_ (.A1(_00654_),
    .A2(_00659_),
    .B1(_06646_),
    .B2(_06654_),
    .Y(_06655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11186_ (.A1(_06640_),
    .A2(_06651_),
    .B1(_06655_),
    .X(_06656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11187_ (.A1(_06589_),
    .A2(_00625_),
    .B1(_06598_),
    .B2(_00634_),
    .X(_06657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11188_ (.A1(_00651_),
    .A2(_04746_),
    .B1(_04743_),
    .B2(_00642_),
    .X(_06658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11189_ (.A(_00599_),
    .Y(_06659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11190_ (.A(_04863_),
    .B(_00608_),
    .X(_06660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11191_ (.A(_06660_),
    .Y(_06661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11192_ (.A1(_00603_),
    .A2(_00608_),
    .B1(_06586_),
    .B2(_00617_),
    .X(_06662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _11193_ (.A1(_04721_),
    .A2(_06659_),
    .B1(_06661_),
    .C1(_06662_),
    .X(_06663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11194_ (.A(_04721_),
    .B(_06659_),
    .Y(_06664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11195_ (.A(_06586_),
    .B(_00617_),
    .X(_06665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11196_ (.A(_00381_),
    .X(_06666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _11197_ (.A1(_06666_),
    .A2(_00582_),
    .B1(_06605_),
    .Y(_06667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11198_ (.A1(_04743_),
    .A2(_00642_),
    .B1(_00651_),
    .B2(_04746_),
    .X(_06668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11199_ (.A1(_06589_),
    .A2(_00625_),
    .B1(_06598_),
    .B2(_00634_),
    .C1(_06668_),
    .X(_06669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and4b_2 _11200_ (.A_N(_06664_),
    .B(_06665_),
    .C(_06667_),
    .D(_06669_),
    .X(_06670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4b_2 _11201_ (.A(_06657_),
    .B(_06658_),
    .C(_06663_),
    .D_N(_06670_),
    .X(_06671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11202_ (.A1(_00637_),
    .A2(_00642_),
    .B1(_06598_),
    .B2(_00634_),
    .C1(_06658_),
    .X(_06672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11203_ (.A1(_00620_),
    .A2(_00625_),
    .B1(_06657_),
    .B2(_06672_),
    .C1(_06665_),
    .X(_06673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11204_ (.A1(_00594_),
    .A2(_00599_),
    .B1(_06662_),
    .B2(_06673_),
    .C1(_06660_),
    .X(_06674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21bai_2 _11205_ (.A1(_06664_),
    .A2(_06674_),
    .B1_N(_06605_),
    .Y(_06675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221ai_2 _11206_ (.A1(_04867_),
    .A2(_06604_),
    .B1(_06656_),
    .B2(_06671_),
    .C1(_06675_),
    .Y(_06676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11207_ (.A(_00839_),
    .Y(_06677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11208_ (.A1(_00802_),
    .A2(_00807_),
    .B1(_04663_),
    .B2(_00824_),
    .X(_06678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11209_ (.A1(_01389_),
    .A2(_00570_),
    .B1(_04808_),
    .B2(_00791_),
    .X(_06679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _11210_ (.A(_06628_),
    .B(_06630_),
    .C(_06679_),
    .X(_06680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2111a_2 _11211_ (.A1(_00333_),
    .A2(_06677_),
    .B1(_06678_),
    .C1(_06680_),
    .D1(_06626_),
    .X(_06681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4b_2 _11212_ (.A(_06620_),
    .B(_06621_),
    .C(_06622_),
    .D_N(_06681_),
    .X(_06682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11213_ (.A(_06651_),
    .B(_06671_),
    .C(_06637_),
    .D(_06682_),
    .X(_06683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11214_ (.A1(_04867_),
    .A2(_06604_),
    .B1(_06605_),
    .B2(_06676_),
    .C1(_06683_),
    .X(_00842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11215_ (.A(_06586_),
    .X(_00612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11216_ (.A(_00845_),
    .Y(_06684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11217_ (.A1(_00603_),
    .A2(_00845_),
    .B1(_04704_),
    .B2(_06684_),
    .X(_06685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11218_ (.A1_N(_00612_),
    .A2_N(_00846_),
    .B1(_00612_),
    .B2(_00846_),
    .X(_06686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11219_ (.A(_06686_),
    .Y(_06687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11220_ (.A(_00843_),
    .Y(_06688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11221_ (.A1(_06666_),
    .A2(_00843_),
    .B1(_04867_),
    .B2(_06688_),
    .X(_06689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11222_ (.A1_N(_04722_),
    .A2_N(_00844_),
    .B1(_04722_),
    .B2(_00844_),
    .X(_06690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11223_ (.A(_06689_),
    .B(_06690_),
    .X(_06691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11224_ (.A(_06691_),
    .Y(_06692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _11225_ (.A1(_00620_),
    .A2(_00847_),
    .B1(_00629_),
    .C1(_00848_),
    .X(_06693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11226_ (.A1_N(_06589_),
    .A2_N(_00847_),
    .B1(_06589_),
    .B2(_00847_),
    .X(_06694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11227_ (.A1_N(_06598_),
    .A2_N(_00848_),
    .B1(_04735_),
    .B2(_00848_),
    .X(_06695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11228_ (.A(_06694_),
    .B(_06695_),
    .X(_06696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11229_ (.A(_00849_),
    .Y(_06697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _11230_ (.A1(_00637_),
    .A2(_00849_),
    .B1(_04746_),
    .B2(_00850_),
    .Y(_06698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11231_ (.A1(_04672_),
    .A2(_06697_),
    .B1(_06698_),
    .Y(_06699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11232_ (.A(_06696_),
    .B(_06699_),
    .X(_06700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11233_ (.A1(_04672_),
    .A2(_06697_),
    .B1(_00637_),
    .B2(_00849_),
    .X(_06701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11234_ (.A1_N(_00646_),
    .A2_N(_00850_),
    .B1(_00646_),
    .B2(_00850_),
    .X(_06702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11235_ (.A(_00851_),
    .Y(_06703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11236_ (.A(_04691_),
    .B(_06703_),
    .Y(_06704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _11237_ (.A1(_04691_),
    .A2(_06703_),
    .B1(_06704_),
    .X(_06705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11238_ (.A1_N(_06593_),
    .A2_N(_00852_),
    .B1(_04768_),
    .B2(_00852_),
    .X(_06706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11239_ (.A(_06705_),
    .B(_06706_),
    .X(_06707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11240_ (.A(_00853_),
    .Y(_06708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11241_ (.A(_00854_),
    .Y(_06709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11242_ (.A1(_04697_),
    .A2(_06708_),
    .B1(_04693_),
    .B2(_06709_),
    .X(_06710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11243_ (.A1(_04697_),
    .A2(_06708_),
    .B1(_06710_),
    .Y(_06711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11244_ (.A1(_00671_),
    .A2(_00853_),
    .B1(_04697_),
    .B2(_06708_),
    .X(_06712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11245_ (.A1(_04693_),
    .A2(_06709_),
    .B1(_04764_),
    .B2(_00854_),
    .X(_06713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11246_ (.A(_06712_),
    .B(_06713_),
    .C(_06707_),
    .X(_06714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11247_ (.A(_00855_),
    .Y(_06715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11248_ (.A(_04680_),
    .B(_06715_),
    .Y(_06716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _11249_ (.A1(_04680_),
    .A2(_06715_),
    .B1(_06716_),
    .X(_06717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11250_ (.A1_N(_04750_),
    .A2_N(_00856_),
    .B1(_04750_),
    .B2(_00856_),
    .X(_06718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11251_ (.A(_06717_),
    .B(_06718_),
    .X(_06719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11252_ (.A(_00857_),
    .Y(_06720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11253_ (.A(_00858_),
    .Y(_06721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11254_ (.A1(_04678_),
    .A2(_06720_),
    .B1(_04682_),
    .B2(_06721_),
    .X(_06722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11255_ (.A1(_04678_),
    .A2(_06720_),
    .B1(_06722_),
    .Y(_06723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _11256_ (.A1(_04842_),
    .A2(_00859_),
    .B1(_06556_),
    .C1(_00860_),
    .X(_06724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11257_ (.A1_N(_04842_),
    .A2_N(_00859_),
    .B1(_04842_),
    .B2(_00859_),
    .X(_06725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11258_ (.A1_N(_06556_),
    .A2_N(_00860_),
    .B1(_04775_),
    .B2(_00860_),
    .X(_06726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11259_ (.A(_06725_),
    .B(_06726_),
    .X(_06727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11260_ (.A(_00861_),
    .Y(_06728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _11261_ (.A1(_04782_),
    .A2(_00861_),
    .B1(_06557_),
    .B2(_00862_),
    .Y(_06729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11262_ (.A1(_04656_),
    .A2(_06728_),
    .B1(_06729_),
    .Y(_06730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11263_ (.A(_06727_),
    .B(_06730_),
    .X(_06731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11264_ (.A1(_04656_),
    .A2(_06728_),
    .B1(_04782_),
    .B2(_00861_),
    .X(_06732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11265_ (.A1_N(_06557_),
    .A2_N(_00862_),
    .B1(_06557_),
    .B2(_00862_),
    .X(_06733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11266_ (.A(_06732_),
    .B(_06733_),
    .C(_06727_),
    .D(_06579_),
    .X(_06734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2111a_2 _11267_ (.A1(_00722_),
    .A2(_00859_),
    .B1(_06724_),
    .C1(_06731_),
    .D1(_06734_),
    .X(_06735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11268_ (.A1(_00705_),
    .A2(_00857_),
    .B1(_04678_),
    .B2(_06720_),
    .X(_06736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11269_ (.A1(_04682_),
    .A2(_06721_),
    .B1(_04758_),
    .B2(_00858_),
    .X(_06737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11270_ (.A(_06736_),
    .B(_06737_),
    .C(_06719_),
    .X(_06738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _11271_ (.A1(_04750_),
    .A2(_00856_),
    .A3(_06716_),
    .B1(_04849_),
    .B2(_00855_),
    .X(_06739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11272_ (.A1(_06719_),
    .A2(_06723_),
    .B1(_06735_),
    .B2(_06738_),
    .C1(_06739_),
    .X(_06740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _11273_ (.A1(_06593_),
    .A2(_00852_),
    .A3(_06704_),
    .B1(_04771_),
    .B2(_00851_),
    .X(_06741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11274_ (.A1(_06707_),
    .A2(_06711_),
    .B1(_06714_),
    .B2(_06740_),
    .C1(_06741_),
    .X(_06742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11275_ (.A(_06701_),
    .B(_06702_),
    .C(_06696_),
    .D(_06742_),
    .X(_06743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2111a_2 _11276_ (.A1(_00620_),
    .A2(_00847_),
    .B1(_06693_),
    .C1(_06700_),
    .D1(_06743_),
    .X(_06744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11277_ (.A(_06744_),
    .Y(_06745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _11278_ (.A1(_00603_),
    .A2(_00845_),
    .B1(_06586_),
    .B2(_00846_),
    .Y(_06746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11279_ (.A1(_04704_),
    .A2(_06684_),
    .B1(_06746_),
    .Y(_06747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _11280_ (.A1(_06666_),
    .A2(_00843_),
    .B1(_00594_),
    .C1(_00844_),
    .X(_06748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221ai_2 _11281_ (.A1(_06666_),
    .A2(_00843_),
    .B1(_06691_),
    .B2(_06747_),
    .C1(_06748_),
    .Y(_06749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a41o_2 _11282_ (.A1(_06685_),
    .A2(_06687_),
    .A3(_06692_),
    .A4(_06745_),
    .B1(_06749_),
    .X(_00863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11283_ (.A(\design_top.core0.FCT3[0] ),
    .Y(_06750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11284_ (.A(\design_top.core0.FCT3[2] ),
    .X(_06751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _11285_ (.A(_05446_),
    .B(_06750_),
    .C(_06751_),
    .X(_00864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11286_ (.A(_06676_),
    .B(_06683_),
    .X(_00865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _11287_ (.A(_05446_),
    .B(\design_top.core0.FCT3[0] ),
    .C(\design_top.core0.FCT3[2] ),
    .X(_00866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11288_ (.A(_06751_),
    .B(_00539_),
    .Y(_00537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11289_ (.A1(_00332_),
    .A2(_04626_),
    .B1(_00329_),
    .B2(_00304_),
    .X(_06752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11290_ (.A(_06752_),
    .Y(_00867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11291_ (.A(_06566_),
    .B(_00867_),
    .X(_06753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11292_ (.A(_06753_),
    .X(_01516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11293_ (.A(_01516_),
    .Y(_06754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11294_ (.A(_00840_),
    .B(_06752_),
    .Y(_01517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11295_ (.A(_06754_),
    .B(_01517_),
    .X(_00868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11296_ (.A(_04651_),
    .Y(_00869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11297_ (.A(_04645_),
    .X(_00870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11298_ (.A(_04643_),
    .Y(_00871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11299_ (.A(_06571_),
    .Y(_00872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11300_ (.A(_04633_),
    .Y(_00874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11301_ (.A(_04637_),
    .X(_00875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11302_ (.A(_04694_),
    .X(_00883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11303_ (.A(_04689_),
    .X(_00885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11304_ (.A(_04675_),
    .X(_00887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11305_ (.A(_04670_),
    .X(_00889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11306_ (.A(_04703_),
    .Y(_00891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11307_ (.A(_04702_),
    .Y(_00894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2b_2 _11308_ (.A_N(_04708_),
    .B(_00868_),
    .Y(_00895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11309_ (.A(_04624_),
    .B(_00539_),
    .Y(_00538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11310_ (.A(_05446_),
    .B(_06750_),
    .X(_06755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11311_ (.A(_06755_),
    .X(_00534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11312_ (.A(_04624_),
    .B(_00534_),
    .Y(_00533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11313_ (.A1(\design_top.core0.XJALR ),
    .A2(\design_top.core0.XJAL ),
    .B1(_00309_),
    .X(_00590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11314_ (.A(_05015_),
    .X(_06756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11315_ (.A(_06756_),
    .X(_00540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11316_ (.A(_06484_),
    .X(_06757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11317_ (.A(_06757_),
    .X(_00535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11318_ (.A(_06485_),
    .X(_06758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11319_ (.A(_06758_),
    .Y(_00907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11320_ (.A(io_out[19]),
    .B(io_out[18]),
    .Y(_06759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11321_ (.A(_06759_),
    .Y(_06760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _11322_ (.A(\design_top.IADDR[4] ),
    .B(_06760_),
    .C(\design_top.IADDR[5] ),
    .X(_06761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11323_ (.A(\design_top.IADDR[6] ),
    .B(_06761_),
    .Y(_06762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11324_ (.A(_06762_),
    .Y(_06763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11325_ (.A(\design_top.IADDR[7] ),
    .B(_06763_),
    .Y(_06764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11326_ (.A(_06764_),
    .Y(_06765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11327_ (.A(\design_top.IADDR[8] ),
    .B(_06765_),
    .Y(_06766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11328_ (.A(_06766_),
    .Y(_06767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11329_ (.A(\design_top.IADDR[9] ),
    .B(_06767_),
    .Y(_06768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11330_ (.A(_06768_),
    .Y(_06769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11331_ (.A(\design_top.IADDR[10] ),
    .B(_06769_),
    .Y(_06770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11332_ (.A(_06770_),
    .Y(_06771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11333_ (.A(\design_top.IADDR[11] ),
    .B(_06771_),
    .Y(_06772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11334_ (.A(_06772_),
    .Y(_06773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11335_ (.A(\design_top.IADDR[12] ),
    .B(_06773_),
    .Y(_06774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11336_ (.A(_06774_),
    .Y(_06775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11337_ (.A(\design_top.IADDR[13] ),
    .B(_06775_),
    .Y(_06776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11338_ (.A(_06776_),
    .Y(_06777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11339_ (.A(\design_top.IADDR[14] ),
    .B(_06777_),
    .Y(_06778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11340_ (.A(_06778_),
    .Y(_06779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11341_ (.A(\design_top.IADDR[15] ),
    .B(_06779_),
    .Y(_06780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11342_ (.A(\design_top.IADDR[16] ),
    .Y(_06781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _11343_ (.A(_06780_),
    .B(_06781_),
    .C_N(\design_top.IADDR[17] ),
    .X(_06782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3b_2 _11344_ (.A_N(_06782_),
    .B(\design_top.IADDR[18] ),
    .C(\design_top.IADDR[19] ),
    .X(_06783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11345_ (.A(\design_top.IADDR[20] ),
    .B(_06783_),
    .Y(_06784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11346_ (.A(_06784_),
    .Y(_06785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11347_ (.A(\design_top.IADDR[21] ),
    .B(_06785_),
    .Y(_06786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11348_ (.A(_06786_),
    .Y(_06787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11349_ (.A(\design_top.IADDR[22] ),
    .B(_06787_),
    .Y(_06788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11350_ (.A(_06788_),
    .Y(_06789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11351_ (.A(\design_top.IADDR[23] ),
    .B(_06789_),
    .Y(_06790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11352_ (.A(\design_top.IADDR[24] ),
    .Y(_06791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _11353_ (.A(_06790_),
    .B(_06791_),
    .C_N(\design_top.IADDR[25] ),
    .X(_06792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3b_2 _11354_ (.A_N(_06792_),
    .B(\design_top.IADDR[26] ),
    .C(\design_top.IADDR[27] ),
    .X(_06793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11355_ (.A(\design_top.IADDR[28] ),
    .B(_06793_),
    .Y(_06794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11356_ (.A(_06794_),
    .Y(_06795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11357_ (.A(\design_top.IADDR[29] ),
    .B(_06795_),
    .Y(_06796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11358_ (.A1(\design_top.IADDR[29] ),
    .A2(_06795_),
    .B1(_06796_),
    .X(_00908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11359_ (.A(_04729_),
    .B(\design_top.core0.PC[28] ),
    .Y(_06797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11360_ (.A(\design_top.core0.PC[27] ),
    .Y(_06798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11361_ (.A(_04734_),
    .X(_00411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11362_ (.A(\design_top.core0.PC[26] ),
    .Y(_06799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _11363_ (.A1(_00405_),
    .A2(_06798_),
    .B1(_00411_),
    .C1(_06799_),
    .X(_06800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11364_ (.A1(\design_top.core0.SIMM[27] ),
    .A2(\design_top.core0.PC[27] ),
    .B1(_00405_),
    .B2(_06798_),
    .X(_06801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11365_ (.A1(\design_top.core0.SIMM[26] ),
    .A2(\design_top.core0.PC[26] ),
    .B1(_00411_),
    .B2(_06799_),
    .X(_06802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11366_ (.A(_06801_),
    .B(_06802_),
    .X(_06803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11367_ (.A1(_05402_),
    .A2(\design_top.core0.PC[25] ),
    .B1(_05405_),
    .B2(\design_top.core0.PC[24] ),
    .X(_06804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11368_ (.A1(_05402_),
    .A2(\design_top.core0.PC[25] ),
    .B1(_06804_),
    .Y(_06805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11369_ (.A(_06803_),
    .B(_06805_),
    .X(_06806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11370_ (.A1_N(_05402_),
    .A2_N(\design_top.core0.PC[25] ),
    .B1(_05402_),
    .B2(\design_top.core0.PC[25] ),
    .X(_06807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11371_ (.A(_06807_),
    .Y(_06808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11372_ (.A1_N(_05405_),
    .A2_N(\design_top.core0.PC[24] ),
    .B1(\design_top.core0.SIMM[24] ),
    .B2(\design_top.core0.PC[24] ),
    .X(_06809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11373_ (.A(_06809_),
    .Y(_06810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11374_ (.A(_04753_),
    .B(\design_top.core0.PC[19] ),
    .X(_06811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11375_ (.A1(_04753_),
    .A2(\design_top.core0.PC[19] ),
    .B1_N(_06811_),
    .X(_06812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11376_ (.A(_06812_),
    .Y(_06813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11377_ (.A(\design_top.core0.PC[18] ),
    .Y(_06814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11378_ (.A1(_00459_),
    .A2(_06814_),
    .B1(_04751_),
    .B2(\design_top.core0.PC[18] ),
    .X(_06815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11379_ (.A1_N(_05411_),
    .A2_N(\design_top.core0.PC[17] ),
    .B1(_05411_),
    .B2(\design_top.core0.PC[17] ),
    .X(_06816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11380_ (.A1_N(_05414_),
    .A2_N(\design_top.core0.PC[16] ),
    .B1(_05414_),
    .B2(\design_top.core0.PC[16] ),
    .X(_06817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and4_2 _11381_ (.A(_06813_),
    .B(_06815_),
    .C(_06816_),
    .D(_06817_),
    .X(_06818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11382_ (.A1_N(_05408_),
    .A2_N(\design_top.core0.PC[21] ),
    .B1(_05408_),
    .B2(\design_top.core0.PC[21] ),
    .X(_06819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11383_ (.A(_06819_),
    .Y(_06820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11384_ (.A(\design_top.core0.PC[20] ),
    .Y(_06821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11385_ (.A1(_00447_),
    .A2(_06821_),
    .B1(_04765_),
    .B2(\design_top.core0.PC[20] ),
    .X(_06822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11386_ (.A(_06822_),
    .Y(_06823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11387_ (.A(\design_top.core0.PC[22] ),
    .Y(_06824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11388_ (.A1(_04769_),
    .A2(\design_top.core0.PC[22] ),
    .B1(_00435_),
    .B2(_06824_),
    .X(_06825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11389_ (.A(\design_top.core0.PC[23] ),
    .Y(_06826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11390_ (.A1(_04846_),
    .A2(\design_top.core0.PC[23] ),
    .B1(_00429_),
    .B2(_06826_),
    .X(_06827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor4_2 _11391_ (.A(_06820_),
    .B(_06823_),
    .C(_06825_),
    .D(_06827_),
    .Y(_06828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11392_ (.A(_04799_),
    .B(\design_top.core0.PC[11] ),
    .X(_06829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11393_ (.A1(_04799_),
    .A2(\design_top.core0.PC[11] ),
    .B1_N(_06829_),
    .X(_06830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11394_ (.A(_06830_),
    .Y(_06831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11395_ (.A(\design_top.core0.PC[10] ),
    .Y(_06832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11396_ (.A1(_00507_),
    .A2(_06832_),
    .B1(\design_top.core0.SIMM[10] ),
    .B2(\design_top.core0.PC[10] ),
    .X(_06833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11397_ (.A1_N(_05382_),
    .A2_N(\design_top.core0.PC[9] ),
    .B1(_05382_),
    .B2(\design_top.core0.PC[9] ),
    .X(_06834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11398_ (.A1_N(_05386_),
    .A2_N(\design_top.core0.PC[8] ),
    .B1(_05386_),
    .B2(\design_top.core0.PC[8] ),
    .X(_06835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and4_2 _11399_ (.A(_06831_),
    .B(_06833_),
    .C(_06834_),
    .D(_06835_),
    .X(_06836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11400_ (.A1_N(_05417_),
    .A2_N(\design_top.core0.PC[13] ),
    .B1(_05417_),
    .B2(\design_top.core0.PC[13] ),
    .X(_06837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11401_ (.A(_06837_),
    .Y(_06838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11402_ (.A(\design_top.core0.PC[12] ),
    .Y(_06839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11403_ (.A1(_00495_),
    .A2(_06839_),
    .B1(_04786_),
    .B2(\design_top.core0.PC[12] ),
    .X(_06840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11404_ (.A(_06840_),
    .Y(_06841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11405_ (.A(\design_top.core0.PC[14] ),
    .Y(_06842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11406_ (.A1(_04776_),
    .A2(\design_top.core0.PC[14] ),
    .B1(_00483_),
    .B2(_06842_),
    .X(_06843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11407_ (.A(\design_top.core0.PC[15] ),
    .Y(_06844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11408_ (.A1(_04841_),
    .A2(\design_top.core0.PC[15] ),
    .B1(_00477_),
    .B2(_06844_),
    .X(_06845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor4_2 _11409_ (.A(_06838_),
    .B(_06841_),
    .C(_06843_),
    .D(_06845_),
    .Y(_06846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11410_ (.A1_N(_05388_),
    .A2_N(\design_top.core0.PC[7] ),
    .B1(_05388_),
    .B2(\design_top.core0.PC[7] ),
    .X(_06847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11411_ (.A1_N(_05389_),
    .A2_N(\design_top.core0.PC[6] ),
    .B1(_05389_),
    .B2(\design_top.core0.PC[6] ),
    .X(_06848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11412_ (.A1_N(_05391_),
    .A2_N(\design_top.core0.PC[5] ),
    .B1(_05391_),
    .B2(\design_top.core0.PC[5] ),
    .X(_06849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11413_ (.A1_N(_05392_),
    .A2_N(\design_top.core0.PC[4] ),
    .B1(_05392_),
    .B2(\design_top.core0.PC[4] ),
    .X(_06850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11414_ (.A(_04811_),
    .B(\design_top.core0.PC[3] ),
    .Y(_06851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11415_ (.A(_04814_),
    .B(\design_top.core0.PC[2] ),
    .Y(_06852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11416_ (.A1_N(_04817_),
    .A2_N(\design_top.core0.PC[1] ),
    .B1(_04817_),
    .B2(\design_top.core0.PC[1] ),
    .X(_06853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11417_ (.A(\design_top.core0.PC[0] ),
    .Y(_06854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11418_ (.A(_04818_),
    .B(_06854_),
    .Y(_06855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11419_ (.A1(_04817_),
    .A2(\design_top.core0.PC[1] ),
    .B1(_06853_),
    .B2(_06855_),
    .X(_06856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11420_ (.A(_06856_),
    .Y(_06857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11421_ (.A1_N(_04814_),
    .A2_N(\design_top.core0.PC[2] ),
    .B1(_06852_),
    .B2(_06857_),
    .X(_06858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2ai_2 _11422_ (.A1_N(_04811_),
    .A2_N(\design_top.core0.PC[3] ),
    .B1(_06851_),
    .B2(_06858_),
    .Y(_06859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11423_ (.A(_05391_),
    .B(\design_top.core0.PC[5] ),
    .X(_06860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a32o_2 _11424_ (.A1(_05392_),
    .A2(\design_top.core0.PC[4] ),
    .A3(_06860_),
    .B1(_05391_),
    .B2(\design_top.core0.PC[5] ),
    .X(_06861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _11425_ (.A1(_06849_),
    .A2(_06850_),
    .A3(_06859_),
    .B1(_06861_),
    .X(_06862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11426_ (.A(_05388_),
    .B(\design_top.core0.PC[7] ),
    .X(_06863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a32o_2 _11427_ (.A1(_05389_),
    .A2(\design_top.core0.PC[6] ),
    .A3(_06863_),
    .B1(_05388_),
    .B2(\design_top.core0.PC[7] ),
    .X(_06864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _11428_ (.A1(_06847_),
    .A2(_06848_),
    .A3(_06862_),
    .B1(_06864_),
    .X(_06865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11429_ (.A1(_05382_),
    .A2(\design_top.core0.PC[9] ),
    .B1(_05386_),
    .B2(\design_top.core0.PC[8] ),
    .X(_06866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11430_ (.A1(_05382_),
    .A2(\design_top.core0.PC[9] ),
    .B1(_06866_),
    .X(_06867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a32o_2 _11431_ (.A1(\design_top.core0.SIMM[10] ),
    .A2(\design_top.core0.PC[10] ),
    .A3(_06829_),
    .B1(_04799_),
    .B2(\design_top.core0.PC[11] ),
    .X(_06868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _11432_ (.A1(_06831_),
    .A2(_06833_),
    .A3(_06867_),
    .B1(_06868_),
    .X(_06869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11433_ (.A1(_05417_),
    .A2(\design_top.core0.PC[13] ),
    .B1(_04786_),
    .B2(\design_top.core0.PC[12] ),
    .X(_06870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11434_ (.A1(_05417_),
    .A2(\design_top.core0.PC[13] ),
    .B1(_06870_),
    .X(_06871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _11435_ (.A1(_06837_),
    .A2(_06840_),
    .A3(_06869_),
    .B1(_06871_),
    .X(_06872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11436_ (.A1(_04776_),
    .A2(\design_top.core0.PC[14] ),
    .B1(_06872_),
    .X(_06873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11437_ (.A1(_04776_),
    .A2(\design_top.core0.PC[14] ),
    .B1(_04841_),
    .B2(\design_top.core0.PC[15] ),
    .X(_06874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11438_ (.A1(_04841_),
    .A2(\design_top.core0.PC[15] ),
    .B1(_06873_),
    .B2(_06874_),
    .X(_06875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _11439_ (.A1(_06836_),
    .A2(_06846_),
    .A3(_06865_),
    .B1(_06875_),
    .X(_06876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11440_ (.A1(_05411_),
    .A2(\design_top.core0.PC[17] ),
    .B1(\design_top.core0.SIMM[16] ),
    .B2(\design_top.core0.PC[16] ),
    .X(_06877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11441_ (.A1(_05411_),
    .A2(\design_top.core0.PC[17] ),
    .B1(_06877_),
    .X(_06878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a32o_2 _11442_ (.A1(_04751_),
    .A2(\design_top.core0.PC[18] ),
    .A3(_06811_),
    .B1(_04753_),
    .B2(\design_top.core0.PC[19] ),
    .X(_06879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _11443_ (.A1(_06813_),
    .A2(_06815_),
    .A3(_06878_),
    .B1(_06879_),
    .X(_06880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11444_ (.A1(_05408_),
    .A2(\design_top.core0.PC[21] ),
    .B1(_04765_),
    .B2(\design_top.core0.PC[20] ),
    .X(_06881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11445_ (.A1(_05408_),
    .A2(\design_top.core0.PC[21] ),
    .B1(_06881_),
    .X(_06882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _11446_ (.A1(_06819_),
    .A2(_06822_),
    .A3(_06880_),
    .B1(_06882_),
    .X(_06883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11447_ (.A1(_04769_),
    .A2(\design_top.core0.PC[22] ),
    .B1(_06883_),
    .X(_06884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11448_ (.A1(_04769_),
    .A2(\design_top.core0.PC[22] ),
    .B1(_04846_),
    .B2(\design_top.core0.PC[23] ),
    .X(_06885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11449_ (.A1(_04846_),
    .A2(\design_top.core0.PC[23] ),
    .B1(_06884_),
    .B2(_06885_),
    .X(_06886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _11450_ (.A1(_06818_),
    .A2(_06828_),
    .A3(_06876_),
    .B1(_06886_),
    .X(_06887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11451_ (.A(_06887_),
    .Y(_06888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11452_ (.A(_06808_),
    .B(_06810_),
    .C(_06803_),
    .D(_06888_),
    .X(_06889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2111a_2 _11453_ (.A1(_00405_),
    .A2(_06798_),
    .B1(_06800_),
    .C1(_06806_),
    .D1(_06889_),
    .X(_06890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11454_ (.A1_N(_04729_),
    .A2_N(\design_top.core0.PC[28] ),
    .B1(_06797_),
    .B2(_06890_),
    .X(_06891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11455_ (.A(_04724_),
    .B(\design_top.core0.PC[29] ),
    .Y(_06892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _11456_ (.A1(_04724_),
    .A2(\design_top.core0.PC[29] ),
    .B1(_06892_),
    .X(_06893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11457_ (.A1_N(_06891_),
    .A2_N(_06893_),
    .B1(_06891_),
    .B2(_06893_),
    .X(_00910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11458_ (.A(_00910_),
    .Y(_00909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11459_ (.A1(_00399_),
    .A2(_00612_),
    .B1(_04862_),
    .B2(_04731_),
    .X(_06894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11460_ (.A(_06894_),
    .Y(_06895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11461_ (.A1(_04727_),
    .A2(_06894_),
    .B1(_04726_),
    .B2(_06895_),
    .X(_00911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11462_ (.A(_06796_),
    .Y(_06896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11463_ (.A(\design_top.IADDR[30] ),
    .B(_06896_),
    .Y(_06897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11464_ (.A1(\design_top.IADDR[30] ),
    .A2(_06896_),
    .B1(_06897_),
    .X(_00913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11465_ (.A(\design_top.core0.PC[30] ),
    .Y(_06898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11466_ (.A1(\design_top.core0.SIMM[30] ),
    .A2(\design_top.core0.PC[30] ),
    .B1(_00387_),
    .B2(_06898_),
    .X(_06899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11467_ (.A1_N(_04724_),
    .A2_N(\design_top.core0.PC[29] ),
    .B1(_06891_),
    .B2(_06892_),
    .X(_06900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11468_ (.A1_N(_06899_),
    .A2_N(_06900_),
    .B1(_06899_),
    .B2(_06900_),
    .X(_00914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11469_ (.A(_00914_),
    .Y(_00915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _11470_ (.A1_N(_04723_),
    .A2_N(_04865_),
    .B1(_04723_),
    .B2(_04865_),
    .Y(_00916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11471_ (.A(\design_top.IADDR[31] ),
    .Y(_06901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a32o_2 _11472_ (.A1(\design_top.IADDR[30] ),
    .A2(_06896_),
    .A3(_06901_),
    .B1(\design_top.IADDR[31] ),
    .B2(_06897_),
    .X(_00918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _11473_ (.A1(_00387_),
    .A2(_06898_),
    .B1(_06899_),
    .B2(_06900_),
    .Y(_06902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11474_ (.A1_N(_01360_),
    .A2_N(\design_top.core0.PC[31] ),
    .B1(_01360_),
    .B2(\design_top.core0.PC[31] ),
    .X(_06903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11475_ (.A1_N(_06902_),
    .A2_N(_06903_),
    .B1(_06902_),
    .B2(_06903_),
    .X(_00919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11476_ (.A(_00919_),
    .Y(_00920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11477_ (.A(_05539_),
    .B(_05512_),
    .X(_00922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11478_ (.A(_04678_),
    .B(_00711_),
    .Y(_00712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11479_ (.A(_04680_),
    .B(_00694_),
    .Y(_00695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11480_ (.A(_04693_),
    .B(_00686_),
    .Y(_00687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11481_ (.A(_04697_),
    .B(_00677_),
    .Y(_00678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11482_ (.A(_04688_),
    .B(_00669_),
    .Y(_00670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11483_ (.A(_04691_),
    .B(_00660_),
    .Y(_00661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11484_ (.A(_04674_),
    .B(_00652_),
    .Y(_00653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11485_ (.A(_04672_),
    .B(_00643_),
    .Y(_00644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11486_ (.A(_00410_),
    .B(_00635_),
    .Y(_00636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11487_ (.A(_00404_),
    .B(_00626_),
    .Y(_00627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11488_ (.A(_04704_),
    .B(_00609_),
    .Y(_00610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11489_ (.A(_04721_),
    .B(_00600_),
    .Y(_00601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _11490_ (.A1(_00326_),
    .A2(_04819_),
    .B1(_04820_),
    .C1(_04822_),
    .X(_06904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11491_ (.A(_06904_),
    .X(_06905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11492_ (.A(_06905_),
    .Y(_00545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11493_ (.A(_05016_),
    .X(_00552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11494_ (.A(_06757_),
    .X(_06906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _11495_ (.A(_00839_),
    .B(_06906_),
    .C(_00540_),
    .X(_01055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11496_ (.A(_06751_),
    .B(_00534_),
    .Y(_00532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11497_ (.A(_06677_),
    .X(_06907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11498_ (.A(_05274_),
    .X(_06908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11499_ (.A(_06908_),
    .X(_06909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11500_ (.A(_06907_),
    .B(_06909_),
    .Y(_01056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _11501_ (.A(_00832_),
    .B(_06906_),
    .C(_00540_),
    .X(_01058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11502_ (.A(_06623_),
    .X(_06910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11503_ (.A(_06910_),
    .B(_06909_),
    .Y(_01059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11504_ (.A(_06484_),
    .X(_06911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _11505_ (.A(_00824_),
    .B(_06911_),
    .C(_00540_),
    .X(_01061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11506_ (.A(_00824_),
    .Y(_06912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11507_ (.A(_06912_),
    .B(_06909_),
    .Y(_01062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _11508_ (.A(_00815_),
    .B(_06911_),
    .C(_00540_),
    .X(_01064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11509_ (.A(_00815_),
    .Y(_06913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11510_ (.A(_06913_),
    .B(_06909_),
    .Y(_01065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _11511_ (.A(_00807_),
    .B(_06911_),
    .C(_06756_),
    .X(_01067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11512_ (.A(_00807_),
    .Y(_06914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11513_ (.A(_06914_),
    .B(_06909_),
    .Y(_01068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _11514_ (.A(_00798_),
    .B(_06911_),
    .C(_06756_),
    .X(_01070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11515_ (.A(_00798_),
    .Y(_06915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11516_ (.A(_06908_),
    .X(_06916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11517_ (.A(_06915_),
    .B(_06916_),
    .Y(_01071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _11518_ (.A(_00791_),
    .B(_06911_),
    .C(_06756_),
    .X(_01073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11519_ (.A(_00791_),
    .Y(_06917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11520_ (.A(_06917_),
    .B(_06916_),
    .Y(_01074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _11521_ (.A(_00570_),
    .B(_06757_),
    .C(_06756_),
    .X(_01076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11522_ (.A(_00570_),
    .Y(_06918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11523_ (.A(_06918_),
    .B(_06916_),
    .Y(_01077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11524_ (.A(\design_top.TIMER[0] ),
    .Y(_01079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11525_ (.A1(\design_top.TIMER[1] ),
    .A2(\design_top.TIMER[0] ),
    .B1_N(_05037_),
    .X(_01080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11526_ (.A1(\design_top.TIMER[2] ),
    .A2(_05037_),
    .B1_N(_05038_),
    .X(_01081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11527_ (.A1(\design_top.TIMER[3] ),
    .A2(_05038_),
    .B1_N(_05039_),
    .X(_01082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11528_ (.A1(\design_top.TIMER[4] ),
    .A2(_05039_),
    .B1_N(_05040_),
    .X(_01083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11529_ (.A1(\design_top.TIMER[5] ),
    .A2(_05040_),
    .B1_N(_05041_),
    .X(_01084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11530_ (.A1(\design_top.TIMER[6] ),
    .A2(_05041_),
    .B1_N(_05042_),
    .X(_01085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11531_ (.A1(\design_top.TIMER[7] ),
    .A2(_05042_),
    .B1_N(_05043_),
    .X(_01086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11532_ (.A1(\design_top.TIMER[8] ),
    .A2(_05043_),
    .B1_N(_05044_),
    .X(_01087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11533_ (.A1(\design_top.TIMER[9] ),
    .A2(_05044_),
    .B1_N(_05045_),
    .X(_01088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11534_ (.A1(\design_top.TIMER[10] ),
    .A2(_05045_),
    .B1_N(_05046_),
    .X(_01089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11535_ (.A1(\design_top.TIMER[11] ),
    .A2(_05046_),
    .B1_N(_05047_),
    .X(_01090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11536_ (.A1(\design_top.TIMER[12] ),
    .A2(_05047_),
    .B1_N(_05048_),
    .X(_01091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11537_ (.A1(\design_top.TIMER[13] ),
    .A2(_05048_),
    .B1_N(_05049_),
    .X(_01092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11538_ (.A1(\design_top.TIMER[14] ),
    .A2(_05049_),
    .B1_N(_05050_),
    .X(_01093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11539_ (.A1(\design_top.TIMER[15] ),
    .A2(_05050_),
    .B1_N(_05051_),
    .X(_01094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11540_ (.A(\design_top.TIMER[16] ),
    .B(_05051_),
    .X(_06919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11541_ (.A1(\design_top.TIMER[16] ),
    .A2(_05051_),
    .B1_N(_06919_),
    .X(_01095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11542_ (.A(\design_top.TIMER[17] ),
    .B(_06919_),
    .X(_06920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11543_ (.A1(\design_top.TIMER[17] ),
    .A2(_06919_),
    .B1_N(_06920_),
    .X(_01096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11544_ (.A(\design_top.TIMER[18] ),
    .B(_06920_),
    .X(_06921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11545_ (.A1(\design_top.TIMER[18] ),
    .A2(_06920_),
    .B1_N(_06921_),
    .X(_01097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11546_ (.A1(\design_top.TIMER[19] ),
    .A2(_06921_),
    .B1_N(_05052_),
    .X(_01098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11547_ (.A(\design_top.TIMER[20] ),
    .B(_05052_),
    .X(_06922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11548_ (.A1(\design_top.TIMER[20] ),
    .A2(_05052_),
    .B1_N(_06922_),
    .X(_01099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11549_ (.A1(\design_top.TIMER[21] ),
    .A2(_06922_),
    .B1_N(_05053_),
    .X(_01100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11550_ (.A(\design_top.TIMER[22] ),
    .B(_05053_),
    .X(_06923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11551_ (.A1(\design_top.TIMER[22] ),
    .A2(_05053_),
    .B1_N(_06923_),
    .X(_01101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11552_ (.A1(\design_top.TIMER[23] ),
    .A2(_06923_),
    .B1_N(_05054_),
    .X(_01102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11553_ (.A(\design_top.TIMER[24] ),
    .B(_05054_),
    .Y(_06924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _11554_ (.A1(\design_top.TIMER[24] ),
    .A2(_05054_),
    .B1(_06924_),
    .X(_01103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11555_ (.A(\design_top.TIMER[25] ),
    .Y(_06925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11556_ (.A1(_06925_),
    .A2(_06924_),
    .B1(_05055_),
    .Y(_01104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11557_ (.A1(\design_top.TIMER[26] ),
    .A2(_05055_),
    .B1_N(_05056_),
    .X(_01105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11558_ (.A1(\design_top.TIMER[27] ),
    .A2(_05056_),
    .B1_N(_05057_),
    .X(_01106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11559_ (.A(\design_top.TIMER[28] ),
    .B(_05057_),
    .X(_06926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11560_ (.A1(\design_top.TIMER[28] ),
    .A2(_05057_),
    .B1_N(_06926_),
    .X(_01107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11561_ (.A(\design_top.TIMER[29] ),
    .B(_06926_),
    .X(_06927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _11562_ (.A1(\design_top.TIMER[29] ),
    .A2(_06926_),
    .B1_N(_06927_),
    .X(_01108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11563_ (.A1_N(\design_top.TIMER[30] ),
    .A2_N(_06927_),
    .B1(\design_top.TIMER[30] ),
    .B2(_06927_),
    .X(_01109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11564_ (.A1(\design_top.TIMER[30] ),
    .A2(_06927_),
    .B1(\design_top.TIMER[31] ),
    .X(_06928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11565_ (.A(_00345_),
    .B(_06928_),
    .X(_01110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11566_ (.A(_06666_),
    .B(_06585_),
    .X(_00593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11567_ (.A(_04621_),
    .B(_04711_),
    .Y(_00589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11568_ (.A(\design_top.DACK[0] ),
    .B(\design_top.DACK[1] ),
    .Y(_00588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11569_ (.A(\design_top.uart0.UART_XSTATE[0] ),
    .B(_05512_),
    .Y(_00586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11570_ (.A(_06634_),
    .B(_00535_),
    .Y(_00577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11571_ (.A(_05016_),
    .X(_06929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11572_ (.A(_06929_),
    .Y(_00551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11573_ (.A(_06918_),
    .B(_00552_),
    .Y(_00571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11574_ (.A(_06906_),
    .B(_00534_),
    .Y(_00544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11575_ (.A(_06904_),
    .X(_00546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11576_ (.A(\design_top.IDATA[20] ),
    .Y(_06930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11577_ (.A(_05311_),
    .X(_06931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor4_2 _11578_ (.A(_06930_),
    .B(_00009_),
    .C(_00008_),
    .D(_06931_),
    .Y(_01305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11579_ (.A(_05311_),
    .X(_06932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11580_ (.A(_05350_),
    .B(_06932_),
    .Y(_01306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11581_ (.A(_05345_),
    .B(_06932_),
    .Y(_01309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11582_ (.A(_05342_),
    .B(_06932_),
    .Y(_01312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11583_ (.A(_05340_),
    .B(_06932_),
    .Y(_01316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11584_ (.A(_05338_),
    .B(_06932_),
    .Y(_01319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11585_ (.A(_05311_),
    .X(_06933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11586_ (.A(_05336_),
    .B(_06933_),
    .Y(_01322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11587_ (.A(_05331_),
    .B(_06933_),
    .Y(_01325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11588_ (.A(_05329_),
    .B(_06933_),
    .Y(_01328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11589_ (.A(_05325_),
    .B(_06933_),
    .Y(_01331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11590_ (.A(_05320_),
    .B(_06933_),
    .Y(_01334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11591_ (.A(_05311_),
    .X(_06934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11592_ (.A(_05300_),
    .B(_06934_),
    .Y(_01337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11593_ (.A(\design_top.IDATA[12] ),
    .B(_06934_),
    .X(_01340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11594_ (.A(\design_top.IDATA[13] ),
    .B(_06934_),
    .X(_01343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11595_ (.A(\design_top.IDATA[14] ),
    .B(_06934_),
    .X(_01345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11596_ (.A(\design_top.IDATA[15] ),
    .B(_06934_),
    .X(_01347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11597_ (.A(\design_top.IDATA[16] ),
    .B(_06931_),
    .X(_01349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11598_ (.A(\design_top.IDATA[17] ),
    .B(_06931_),
    .X(_01351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11599_ (.A(\design_top.IDATA[18] ),
    .B(_06931_),
    .X(_01353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11600_ (.A(_01262_),
    .B(_06931_),
    .X(_01355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11601_ (.A(_06930_),
    .B(_01240_),
    .Y(_01357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11602_ (.A(\design_top.core0.NXPC[31] ),
    .Y(_01359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11603_ (.A(_00833_),
    .X(_06935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11604_ (.A(_06935_),
    .B(_00324_),
    .Y(_01361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11605_ (.A(_00883_),
    .B(_00884_),
    .C(_00885_),
    .D(_00886_),
    .X(_06936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11606_ (.A(_04685_),
    .X(_02137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11607_ (.A(_00881_),
    .B(_00880_),
    .C(_00882_),
    .D(_02137_),
    .X(_06937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11608_ (.A(_00878_),
    .B(_04659_),
    .C(_04653_),
    .D(_00879_),
    .X(_06938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11609_ (.A(_00874_),
    .B(_00873_),
    .C(_00876_),
    .D(_00875_),
    .X(_06939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11610_ (.A(_04664_),
    .Y(_01656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11611_ (.A1(_00834_),
    .A2(_01516_),
    .B1(_01361_),
    .X(_06940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11612_ (.A1(_01656_),
    .A2(_06940_),
    .B1(_01655_),
    .X(_06941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11613_ (.A1(_00869_),
    .A2(_06941_),
    .B1(_00818_),
    .Y(_06942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11614_ (.A(_06942_),
    .Y(_06943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11615_ (.A(_04640_),
    .X(_01846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11616_ (.A(_00871_),
    .B(_00870_),
    .C(_01846_),
    .D(_00872_),
    .X(_06944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _11617_ (.A1(_00801_),
    .A2(_01758_),
    .B1(_00800_),
    .X(_06945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _11618_ (.A1(_01845_),
    .A2(_06945_),
    .B1(_00793_),
    .C1(_00784_),
    .X(_06946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _11619_ (.A1(_06943_),
    .A2(_06944_),
    .B1(_00785_),
    .C1(_06946_),
    .X(_06947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _11620_ (.A1(_00774_),
    .A2(_01914_),
    .B1(_00773_),
    .Y(_06948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11621_ (.A(_04636_),
    .B(_06948_),
    .Y(_06949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _11622_ (.A1(_00757_),
    .A2(_00766_),
    .A3(_06949_),
    .B1(_00758_),
    .X(_06950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _11623_ (.A1(_00742_),
    .A2(_02005_),
    .B1(_00741_),
    .X(_06951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _11624_ (.A1(_02053_),
    .A2(_06951_),
    .B1(_00733_),
    .C1(_00724_),
    .X(_06952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _11625_ (.A1(_06938_),
    .A2(_06950_),
    .B1(_00725_),
    .C1(_06952_),
    .X(_06953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _11626_ (.A1(_06938_),
    .A2(_06939_),
    .A3(_06947_),
    .B1(_06953_),
    .X(_06954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _11627_ (.A1(_00713_),
    .A2(_02094_),
    .B1(_00712_),
    .Y(_06955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11628_ (.A(_04684_),
    .B(_06955_),
    .Y(_06956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _11629_ (.A1(_00695_),
    .A2(_00704_),
    .A3(_06956_),
    .B1(_00696_),
    .X(_06957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _11630_ (.A1(_02178_),
    .A2(_00679_),
    .B1(_00678_),
    .X(_06958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _11631_ (.A1(_02220_),
    .A2(_06958_),
    .B1(_00670_),
    .C1(_00661_),
    .X(_06959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _11632_ (.A1(_06936_),
    .A2(_06957_),
    .B1(_00662_),
    .C1(_06959_),
    .X(_06960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _11633_ (.A1(_06936_),
    .A2(_06937_),
    .A3(_06954_),
    .B1(_06960_),
    .X(_06961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11634_ (.A(_04675_),
    .B(_00888_),
    .C(_00890_),
    .D(_00889_),
    .X(_06962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _11635_ (.A1(_02260_),
    .A2(_00645_),
    .B1(_00644_),
    .X(_06963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _11636_ (.A1(_00636_),
    .A2(_06963_),
    .B1(_00628_),
    .C1(_02302_),
    .X(_06964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11637_ (.A1(_06961_),
    .A2(_06962_),
    .B1(_00627_),
    .B2(_06964_),
    .X(_06965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11638_ (.A(_00398_),
    .B(_00618_),
    .Y(_02343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11639_ (.A1(_00619_),
    .A2(_06965_),
    .B1(_02343_),
    .Y(_06966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11640_ (.A(_06966_),
    .Y(_06967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11641_ (.A1(_00610_),
    .A2(_06967_),
    .B1(_00611_),
    .X(_06968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11642_ (.A1(_00893_),
    .A2(_06968_),
    .B1(_00602_),
    .X(_06969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11643_ (.A1_N(_00894_),
    .A2_N(_06969_),
    .B1(_00894_),
    .B2(_06969_),
    .X(_01362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11644_ (.A(_05421_),
    .B(_05436_),
    .Y(_01363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11645_ (.A(_06685_),
    .Y(_06970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _11646_ (.A1(_06970_),
    .A2(_06686_),
    .A3(_06744_),
    .B1(_06747_),
    .X(_06971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11647_ (.A1(_00594_),
    .A2(_00844_),
    .B1(_06690_),
    .B2(_06971_),
    .X(_06972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11648_ (.A1_N(_06689_),
    .A2_N(_06972_),
    .B1(_06689_),
    .B2(_06972_),
    .X(_01364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11649_ (.A(_00381_),
    .B(_00840_),
    .X(_01400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11650_ (.A(_06935_),
    .B(_01400_),
    .X(_01401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11651_ (.A(_06562_),
    .B(_01401_),
    .X(_01402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11652_ (.A(_04649_),
    .X(_06973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11653_ (.A(_06973_),
    .B(_01402_),
    .X(_01403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11654_ (.A(_06559_),
    .B(_01403_),
    .X(_01404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _11655_ (.A(\design_top.core0.FCT3[1] ),
    .B(_06750_),
    .C(_04624_),
    .X(_06974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11656_ (.A(_06974_),
    .X(_06975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11657_ (.A(_06975_),
    .X(_01407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _11658_ (.A(_05446_),
    .B(\design_top.core0.FCT3[0] ),
    .C(_04624_),
    .X(_06976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11659_ (.A(_06976_),
    .X(_06977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11660_ (.A(_06977_),
    .X(_01408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11661_ (.A(_01406_),
    .B(_01407_),
    .C(_01408_),
    .X(_01409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11662_ (.A(\design_top.RAMFF[31] ),
    .Y(_01412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11663_ (.A(\design_top.XADDR[2] ),
    .B(\design_top.XADDR[3] ),
    .Y(_01413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11664_ (.A(\design_top.IOMUX[3][31] ),
    .Y(_06978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11665_ (.A(\design_top.XADDR[2] ),
    .Y(_01571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11666_ (.A(\design_top.XADDR[3] ),
    .Y(_06979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11667_ (.A(_01571_),
    .B(_06979_),
    .X(_06980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11668_ (.A(_06980_),
    .X(_06981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11669_ (.A(_06981_),
    .X(_06982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11670_ (.A(\design_top.GPIOFF[15] ),
    .Y(_06983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11671_ (.A(\design_top.XADDR[2] ),
    .B(_06979_),
    .X(_06984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11672_ (.A(_06984_),
    .X(_06985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11673_ (.A(_06985_),
    .X(_06986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11674_ (.A1(_06978_),
    .A2(_06982_),
    .B1(_06983_),
    .B2(_06986_),
    .X(_01414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11675_ (.A(\design_top.RAMFF[15] ),
    .Y(_01417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11676_ (.A(\design_top.IOMUX[3][15] ),
    .Y(_06987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11677_ (.A(_06980_),
    .X(_06988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11678_ (.A(\design_top.LEDFF[15] ),
    .Y(_06989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11679_ (.A(_06984_),
    .X(_06990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11680_ (.A(_01571_),
    .B(\design_top.XADDR[3] ),
    .Y(_06991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11681_ (.A(_06991_),
    .X(_06992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11682_ (.A(\design_top.uart0.UART_RFIFO[7] ),
    .B(_06992_),
    .Y(_06993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11683_ (.A1(_06987_),
    .A2(_06988_),
    .B1(_06989_),
    .B2(_06990_),
    .C1(_06993_),
    .X(_01418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11684_ (.A(_06751_),
    .B(_06755_),
    .C(_01420_),
    .X(_01421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11685_ (.A(\design_top.RAMFF[23] ),
    .Y(_01423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11686_ (.A(\design_top.IOMUX[3][23] ),
    .Y(_06994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11687_ (.A(\design_top.GPIOFF[7] ),
    .Y(_06995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11688_ (.A1(_06994_),
    .A2(_06982_),
    .B1(_06995_),
    .B2(_06986_),
    .X(_01424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11689_ (.A(\design_top.RAMFF[7] ),
    .Y(_01426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11690_ (.A(\design_top.IOMUX[3][7] ),
    .Y(_06996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11691_ (.A(\design_top.LEDFF[7] ),
    .Y(_06997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11692_ (.A1(_06996_),
    .A2(_06982_),
    .B1(_06997_),
    .B2(_06986_),
    .X(_01427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11693_ (.A(_06751_),
    .B(_00539_),
    .C(_01431_),
    .X(_01432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _11694_ (.A(_04615_),
    .B(_04616_),
    .C(\design_top.core0.XLUI ),
    .X(_01434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _11695_ (.A(_04615_),
    .B(_04616_),
    .C(\design_top.core0.XAUIPC ),
    .X(_01437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11696_ (.A(_06907_),
    .B(_00546_),
    .Y(_01443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11697_ (.A(_06612_),
    .B(_06916_),
    .Y(_01444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11698_ (.A(_06910_),
    .B(_00546_),
    .Y(_01446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11699_ (.A(_06611_),
    .B(_06916_),
    .Y(_01447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11700_ (.A(_06912_),
    .B(_00546_),
    .Y(_01449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11701_ (.A(_06908_),
    .X(_06998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11702_ (.A(_06610_),
    .B(_06998_),
    .Y(_01450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11703_ (.A(_06913_),
    .B(_00546_),
    .Y(_01452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11704_ (.A(_00755_),
    .Y(_06999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11705_ (.A(_06999_),
    .B(_06998_),
    .Y(_01453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11706_ (.A(_06914_),
    .B(_06905_),
    .Y(_01455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11707_ (.A(_06608_),
    .B(_06998_),
    .Y(_01456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11708_ (.A(_06915_),
    .B(_06905_),
    .Y(_01458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11709_ (.A(_06607_),
    .B(_06998_),
    .Y(_01459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11710_ (.A(_06917_),
    .B(_06905_),
    .Y(_01461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11711_ (.A(_00731_),
    .Y(_07000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11712_ (.A(_07000_),
    .B(_06998_),
    .Y(_01462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11713_ (.A(_06918_),
    .B(_06905_),
    .Y(_01464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11714_ (.A(_06634_),
    .B(_06908_),
    .Y(_01465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11715_ (.A(_06485_),
    .X(_00541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11716_ (.A(_06907_),
    .B(_00541_),
    .Y(_01467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11717_ (.A(_06907_),
    .B(_00535_),
    .Y(_01468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11718_ (.A(_06910_),
    .B(_00541_),
    .Y(_01470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11719_ (.A(_06910_),
    .B(_00535_),
    .Y(_01471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11720_ (.A(_06912_),
    .B(_00541_),
    .Y(_01473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11721_ (.A(_06912_),
    .B(_00535_),
    .Y(_01474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11722_ (.A(_06913_),
    .B(_00541_),
    .Y(_01476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11723_ (.A(_06757_),
    .X(_07001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11724_ (.A(_06913_),
    .B(_07001_),
    .Y(_01477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11725_ (.A(_06914_),
    .B(_06758_),
    .Y(_01479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11726_ (.A(_06914_),
    .B(_07001_),
    .Y(_01480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11727_ (.A(_06915_),
    .B(_06758_),
    .Y(_01482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11728_ (.A(_06915_),
    .B(_07001_),
    .Y(_01483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11729_ (.A(_06917_),
    .B(_06758_),
    .Y(_01485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11730_ (.A(_06917_),
    .B(_07001_),
    .Y(_01486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11731_ (.A(_06918_),
    .B(_06758_),
    .Y(_01488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11732_ (.A(_06918_),
    .B(_07001_),
    .Y(_01489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11733_ (.A(_06907_),
    .B(_00552_),
    .Y(_01491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11734_ (.A(_06757_),
    .X(_07002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11735_ (.A(_06612_),
    .B(_07002_),
    .Y(_01492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11736_ (.A(_06910_),
    .B(_00552_),
    .Y(_01494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11737_ (.A(_06611_),
    .B(_07002_),
    .Y(_01495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11738_ (.A(_06912_),
    .B(_00552_),
    .Y(_01497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11739_ (.A(_06610_),
    .B(_07002_),
    .Y(_01498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11740_ (.A(_06913_),
    .B(_06929_),
    .Y(_01500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11741_ (.A(_06999_),
    .B(_07002_),
    .Y(_01501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11742_ (.A(_06914_),
    .B(_06929_),
    .Y(_01503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11743_ (.A(_06608_),
    .B(_07002_),
    .Y(_01504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11744_ (.A(_06915_),
    .B(_06929_),
    .Y(_01506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11745_ (.A(_06607_),
    .B(_06906_),
    .Y(_01507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11746_ (.A(_06917_),
    .B(_06929_),
    .Y(_01509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11747_ (.A(_07000_),
    .B(_06906_),
    .Y(_01510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11748_ (.A(\design_top.core0.RESMODE[1] ),
    .Y(_07003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11749_ (.A(_05578_),
    .B(_07003_),
    .Y(_01512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11750_ (.A(_00901_),
    .Y(_01513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11751_ (.A(_04615_),
    .B(_04616_),
    .Y(_01514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11752_ (.A(\design_top.core0.NXPC[0] ),
    .Y(_01515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11753_ (.A(_00840_),
    .B(_00867_),
    .X(_01518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11754_ (.A(_06935_),
    .B(_01518_),
    .X(_01519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11755_ (.A(_06562_),
    .B(_01519_),
    .X(_01520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11756_ (.A(_06973_),
    .B(_01520_),
    .X(_01521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11757_ (.A(_06559_),
    .B(_01521_),
    .X(_01522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11758_ (.A(_01553_),
    .X(_01554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11759_ (.A(\design_top.RAMFF[0] ),
    .Y(_01561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11760_ (.A1_N(\design_top.uart0.UART_XREQ ),
    .A2_N(_05699_),
    .B1(\design_top.uart0.UART_XREQ ),
    .B2(_05699_),
    .X(_01562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11761_ (.A(\design_top.IOMUX[3][0] ),
    .Y(_07004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11762_ (.A(io_out[8]),
    .Y(_07005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11763_ (.A(_01571_),
    .B(\design_top.XADDR[3] ),
    .C(_01562_),
    .X(_07006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11764_ (.A1(_07004_),
    .A2(_06988_),
    .B1(_07005_),
    .B2(_06990_),
    .C1(_07006_),
    .X(_01563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11765_ (.A(\design_top.RAMFF[16] ),
    .Y(_01565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11766_ (.A(\design_top.IOMUX[3][16] ),
    .Y(_07007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11767_ (.A(io_out[15]),
    .Y(_07008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11768_ (.A1(_07007_),
    .A2(_06982_),
    .B1(_07008_),
    .B2(_06986_),
    .X(_01566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11769_ (.A(\design_top.RAMFF[24] ),
    .Y(_01570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11770_ (.A(\design_top.IOMUX[3][24] ),
    .Y(_07009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11771_ (.A(\design_top.GPIOFF[8] ),
    .Y(_07010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11772_ (.A1(_07009_),
    .A2(_06982_),
    .B1(_07010_),
    .B2(_06986_),
    .X(_01572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11773_ (.A(\design_top.RAMFF[8] ),
    .Y(_01575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11774_ (.A(\design_top.IOMUX[3][8] ),
    .Y(_07011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11775_ (.A(\design_top.LEDFF[8] ),
    .Y(_07012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11776_ (.A(\design_top.uart0.UART_RFIFO[0] ),
    .B(_06992_),
    .Y(_07013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11777_ (.A1(_07011_),
    .A2(_06988_),
    .B1(_07012_),
    .B2(_06990_),
    .C1(_07013_),
    .X(_01576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _11778_ (.A1(_00326_),
    .A2(_06854_),
    .B1(_06855_),
    .X(_01584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11779_ (.A(\design_top.core0.NXPC[1] ),
    .Y(_01586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11780_ (.A1(_04629_),
    .A2(_06754_),
    .B1(_00834_),
    .B2(_01516_),
    .X(_01588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11781_ (.A1_N(_04629_),
    .A2_N(_06567_),
    .B1(_04629_),
    .B2(_06567_),
    .X(_01589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11782_ (.A(_06935_),
    .B(_01395_),
    .X(_01590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11783_ (.A(_06562_),
    .B(_01590_),
    .X(_01591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11784_ (.A(_06973_),
    .B(_01591_),
    .X(_01592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11785_ (.A(_06559_),
    .B(_01592_),
    .X(_01593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11786_ (.A(_01627_),
    .B(_01407_),
    .C(_01408_),
    .X(_01628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11787_ (.A(\design_top.RAMFF[1] ),
    .Y(_01631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11788_ (.A(\design_top.IOMUX[3][1] ),
    .Y(_07014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11789_ (.A(_06980_),
    .X(_07015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11790_ (.A(io_out[9]),
    .Y(_07016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11791_ (.A(_06984_),
    .X(_07017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11792_ (.A1(\design_top.uart0.UART_RACK ),
    .A2(\design_top.uart0.UART_RREQ ),
    .B1(_06991_),
    .Y(_07018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _11793_ (.A1(\design_top.uart0.UART_RACK ),
    .A2(\design_top.uart0.UART_RREQ ),
    .B1(_07018_),
    .X(_07019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11794_ (.A1(_07014_),
    .A2(_07015_),
    .B1(_07016_),
    .B2(_07017_),
    .C1(_07019_),
    .X(_01632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11795_ (.A(\design_top.RAMFF[17] ),
    .Y(_01634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11796_ (.A(\design_top.IOMUX[3][17] ),
    .Y(_07020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11797_ (.A(_06981_),
    .X(_07021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11798_ (.A(\design_top.GPIOFF[1] ),
    .Y(_07022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11799_ (.A(_06985_),
    .X(_07023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11800_ (.A1(_07020_),
    .A2(_07021_),
    .B1(_07022_),
    .B2(_07023_),
    .X(_01635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11801_ (.A(\design_top.RAMFF[25] ),
    .Y(_01639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11802_ (.A(\design_top.IOMUX[3][25] ),
    .Y(_07024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11803_ (.A(\design_top.GPIOFF[9] ),
    .Y(_07025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11804_ (.A1(_07024_),
    .A2(_07021_),
    .B1(_07025_),
    .B2(_07023_),
    .X(_01640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11805_ (.A(\design_top.RAMFF[9] ),
    .Y(_01643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11806_ (.A(\design_top.IOMUX[3][9] ),
    .Y(_07026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11807_ (.A(\design_top.LEDFF[9] ),
    .Y(_07027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11808_ (.A(\design_top.uart0.UART_RFIFO[1] ),
    .B(_06992_),
    .Y(_07028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11809_ (.A1(_07026_),
    .A2(_07015_),
    .B1(_07027_),
    .B2(_07017_),
    .C1(_07028_),
    .X(_01644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2ai_2 _11810_ (.A1_N(_06853_),
    .A2_N(_06855_),
    .B1(_06853_),
    .B2(_06855_),
    .Y(_01652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11811_ (.A(\design_top.core0.NXPC[2] ),
    .Y(_01654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11812_ (.A1_N(_01656_),
    .A2_N(_06940_),
    .B1(_01656_),
    .B2(_06940_),
    .X(_01657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11813_ (.A1_N(_06565_),
    .A2_N(_06568_),
    .B1(_06565_),
    .B2(_06568_),
    .X(_01658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11814_ (.A(_06562_),
    .B(_01660_),
    .X(_01661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11815_ (.A(_06973_),
    .B(_01661_),
    .X(_01662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11816_ (.A(_06559_),
    .B(_01662_),
    .X(_01663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11817_ (.A(_06935_),
    .B(_01549_),
    .X(_01675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11818_ (.A(_01682_),
    .B(_01407_),
    .C(_01408_),
    .X(_01683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11819_ (.A(\design_top.RAMFF[2] ),
    .Y(_01686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11820_ (.A(\design_top.IOMUX[3][2] ),
    .Y(_07029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11821_ (.A(io_out[10]),
    .Y(_07030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11822_ (.A1(_07029_),
    .A2(_07021_),
    .B1(_07030_),
    .B2(_07023_),
    .X(_01687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11823_ (.A(\design_top.RAMFF[18] ),
    .Y(_01689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11824_ (.A(\design_top.IOMUX[3][18] ),
    .Y(_07031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11825_ (.A(\design_top.GPIOFF[2] ),
    .Y(_07032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11826_ (.A1(_07031_),
    .A2(_07021_),
    .B1(_07032_),
    .B2(_07023_),
    .X(_01690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11827_ (.A(\design_top.RAMFF[26] ),
    .Y(_01695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11828_ (.A(\design_top.IOMUX[3][26] ),
    .Y(_07033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11829_ (.A(\design_top.GPIOFF[10] ),
    .Y(_07034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11830_ (.A1(_07033_),
    .A2(_07021_),
    .B1(_07034_),
    .B2(_07023_),
    .X(_01696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11831_ (.A(\design_top.RAMFF[10] ),
    .Y(_01698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11832_ (.A(\design_top.IOMUX[3][10] ),
    .Y(_04438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11833_ (.A(\design_top.LEDFF[10] ),
    .Y(_04439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _11834_ (.A1(\design_top.uart0.UART_RFIFO[2] ),
    .A2(_06991_),
    .B1(_01413_),
    .Y(_04440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11835_ (.A1(_04438_),
    .A2(_07015_),
    .B1(_04439_),
    .B2(_07017_),
    .C1(_04440_),
    .X(_01699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _11836_ (.A1(_04814_),
    .A2(\design_top.core0.PC[2] ),
    .B1(_06852_),
    .Y(_04441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11837_ (.A1_N(_06856_),
    .A2_N(_04441_),
    .B1(_06856_),
    .B2(_04441_),
    .X(_01707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11838_ (.A(\design_top.core0.NXPC[3] ),
    .Y(_01709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11839_ (.A1_N(_00869_),
    .A2_N(_06941_),
    .B1(_00869_),
    .B2(_06941_),
    .X(_01710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11840_ (.A1_N(_06563_),
    .A2_N(_06569_),
    .B1(_06563_),
    .B2(_06569_),
    .X(_01711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11841_ (.A(_06561_),
    .B(_01396_),
    .X(_01712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11842_ (.A(_06973_),
    .B(_01712_),
    .X(_01713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11843_ (.A(_06558_),
    .X(_04442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11844_ (.A(_04442_),
    .X(_04443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11845_ (.A(_04443_),
    .B(_01713_),
    .X(_01714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11846_ (.A(_01731_),
    .B(_01407_),
    .C(_01408_),
    .X(_01732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11847_ (.A(\design_top.RAMFF[3] ),
    .Y(_01735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11848_ (.A(\design_top.IOMUX[3][3] ),
    .Y(_04444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11849_ (.A(_06981_),
    .X(_04445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11850_ (.A(io_out[11]),
    .Y(_04446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11851_ (.A(_06985_),
    .X(_04447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11852_ (.A1(_04444_),
    .A2(_04445_),
    .B1(_04446_),
    .B2(_04447_),
    .X(_01736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11853_ (.A(\design_top.RAMFF[19] ),
    .Y(_01738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11854_ (.A(\design_top.IOMUX[3][19] ),
    .Y(_04448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11855_ (.A(\design_top.GPIOFF[3] ),
    .Y(_04449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11856_ (.A1(_04448_),
    .A2(_04445_),
    .B1(_04449_),
    .B2(_04447_),
    .X(_01739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11857_ (.A(\design_top.RAMFF[27] ),
    .Y(_01743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11858_ (.A(\design_top.IOMUX[3][27] ),
    .Y(_04450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11859_ (.A(\design_top.GPIOFF[11] ),
    .Y(_04451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11860_ (.A1(_04450_),
    .A2(_04445_),
    .B1(_04451_),
    .B2(_04447_),
    .X(_01744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11861_ (.A(\design_top.RAMFF[11] ),
    .Y(_01746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11862_ (.A(\design_top.IOMUX[3][11] ),
    .Y(_04452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11863_ (.A(\design_top.LEDFF[11] ),
    .Y(_04453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11864_ (.A(\design_top.uart0.UART_RFIFO[3] ),
    .B(_06992_),
    .Y(_04454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11865_ (.A1(_04452_),
    .A2(_07015_),
    .B1(_04453_),
    .B2(_07017_),
    .C1(_04454_),
    .X(_01747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _11866_ (.A1(_04811_),
    .A2(\design_top.core0.PC[3] ),
    .B1(_06851_),
    .X(_04455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11867_ (.A1_N(_06858_),
    .A2_N(_04455_),
    .B1(_06858_),
    .B2(_04455_),
    .X(_02409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11868_ (.A(_02409_),
    .Y(_01755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11869_ (.A(\design_top.core0.NXPC[4] ),
    .Y(_01757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11870_ (.A1(_04646_),
    .A2(_06942_),
    .B1(_00870_),
    .B2(_06943_),
    .X(_01759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11871_ (.A1_N(_04646_),
    .A2_N(_06570_),
    .B1(_04646_),
    .B2(_06570_),
    .X(_01760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11872_ (.A(_04649_),
    .X(_04456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11873_ (.A(_04456_),
    .B(_01763_),
    .X(_01764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11874_ (.A(_04443_),
    .B(_01764_),
    .X(_01765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11875_ (.A(_06561_),
    .B(_01550_),
    .X(_01770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11876_ (.A(_06975_),
    .X(_04457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11877_ (.A(_06977_),
    .X(_04458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11878_ (.A(_01775_),
    .B(_04457_),
    .C(_04458_),
    .X(_01776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11879_ (.A(\design_top.RAMFF[4] ),
    .Y(_01779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11880_ (.A(\design_top.IOMUX[3][4] ),
    .Y(_04459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11881_ (.A(\design_top.LEDFF[4] ),
    .Y(_04460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11882_ (.A1(_04459_),
    .A2(_04445_),
    .B1(_04460_),
    .B2(_04447_),
    .X(_01780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11883_ (.A(\design_top.RAMFF[20] ),
    .Y(_01782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11884_ (.A(\design_top.IOMUX[3][20] ),
    .Y(_04461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11885_ (.A(\design_top.GPIOFF[4] ),
    .Y(_04462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11886_ (.A1(_04461_),
    .A2(_04445_),
    .B1(_04462_),
    .B2(_04447_),
    .X(_01783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11887_ (.A(\design_top.RAMFF[28] ),
    .Y(_01787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11888_ (.A(\design_top.IOMUX[3][28] ),
    .Y(_04463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11889_ (.A(_06980_),
    .X(_04464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11890_ (.A(\design_top.GPIOFF[12] ),
    .Y(_04465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11891_ (.A(_06984_),
    .X(_04466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11892_ (.A1(_04463_),
    .A2(_04464_),
    .B1(_04465_),
    .B2(_04466_),
    .X(_01788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11893_ (.A(\design_top.RAMFF[12] ),
    .Y(_01790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11894_ (.A(\design_top.IOMUX[3][12] ),
    .Y(_04467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11895_ (.A(\design_top.LEDFF[12] ),
    .Y(_04468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11896_ (.A(\design_top.uart0.UART_RFIFO[4] ),
    .B(_06992_),
    .Y(_04469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11897_ (.A1(_04467_),
    .A2(_07015_),
    .B1(_04468_),
    .B2(_07017_),
    .C1(_04469_),
    .X(_01791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11898_ (.A1_N(_06859_),
    .A2_N(_06850_),
    .B1(_06859_),
    .B2(_06850_),
    .X(_02412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11899_ (.A(_02412_),
    .Y(_01799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11900_ (.A(\design_top.core0.NXPC[5] ),
    .Y(_01801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11901_ (.A(_04643_),
    .X(_04470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11902_ (.A1(_00870_),
    .A2(_06943_),
    .B1(_01758_),
    .Y(_04471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11903_ (.A1_N(_04470_),
    .A2_N(_04471_),
    .B1(_04470_),
    .B2(_04471_),
    .X(_01802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11904_ (.A1(_00802_),
    .A2(_00808_),
    .B1(_04646_),
    .B2(_06570_),
    .X(_04472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11905_ (.A1_N(_04470_),
    .A2_N(_04472_),
    .B1(_04470_),
    .B2(_04472_),
    .X(_01803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11906_ (.A(_04456_),
    .B(_01805_),
    .X(_01806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11907_ (.A(_04443_),
    .B(_01806_),
    .X(_01807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11908_ (.A(_06561_),
    .B(_01620_),
    .X(_01812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11909_ (.A(_01817_),
    .B(_04457_),
    .C(_04458_),
    .X(_01818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11910_ (.A(\design_top.RAMFF[5] ),
    .Y(_01821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11911_ (.A(\design_top.IOMUX[3][5] ),
    .Y(_04473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11912_ (.A(\design_top.LEDFF[5] ),
    .Y(_04474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11913_ (.A1(_04473_),
    .A2(_04464_),
    .B1(_04474_),
    .B2(_04466_),
    .X(_01822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11914_ (.A(\design_top.RAMFF[21] ),
    .Y(_01824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11915_ (.A(\design_top.IOMUX[3][21] ),
    .Y(_04475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11916_ (.A(\design_top.GPIOFF[5] ),
    .Y(_04476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11917_ (.A1(_04475_),
    .A2(_04464_),
    .B1(_04476_),
    .B2(_04466_),
    .X(_01825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11918_ (.A(\design_top.RAMFF[29] ),
    .Y(_01830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11919_ (.A(\design_top.IOMUX[3][29] ),
    .Y(_04477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11920_ (.A(\design_top.GPIOFF[13] ),
    .Y(_04478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11921_ (.A1(_04477_),
    .A2(_04464_),
    .B1(_04478_),
    .B2(_04466_),
    .X(_01831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11922_ (.A(\design_top.RAMFF[13] ),
    .Y(_01833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11923_ (.A(\design_top.IOMUX[3][13] ),
    .Y(_04479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11924_ (.A(\design_top.LEDFF[13] ),
    .Y(_04480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _11925_ (.A1(\design_top.uart0.UART_RFIFO[5] ),
    .A2(_06991_),
    .B1(_01413_),
    .Y(_04481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11926_ (.A1(_04479_),
    .A2(_06981_),
    .B1(_04480_),
    .B2(_06985_),
    .C1(_04481_),
    .X(_01834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11927_ (.A1(_05392_),
    .A2(\design_top.core0.PC[4] ),
    .B1(_06859_),
    .B2(_06850_),
    .X(_04482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11928_ (.A1_N(_06849_),
    .A2_N(_04482_),
    .B1(_06849_),
    .B2(_04482_),
    .X(_02416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11929_ (.A(_02416_),
    .Y(_01842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11930_ (.A(\design_top.core0.NXPC[6] ),
    .Y(_01844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _11931_ (.A1(_00871_),
    .A2(_00870_),
    .A3(_06943_),
    .B1(_06945_),
    .X(_04483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11932_ (.A1_N(_01846_),
    .A2_N(_04483_),
    .B1(_01846_),
    .B2(_04483_),
    .X(_01847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11933_ (.A1(_00799_),
    .A2(_01391_),
    .B1(_04470_),
    .B2(_04472_),
    .X(_04484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11934_ (.A1_N(_04641_),
    .A2_N(_04484_),
    .B1(_04641_),
    .B2(_04484_),
    .X(_01848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11935_ (.A(_04456_),
    .B(_01851_),
    .X(_01852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11936_ (.A(_04443_),
    .B(_01852_),
    .X(_01853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11937_ (.A(_06561_),
    .B(_01675_),
    .X(_01858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11938_ (.A(_01863_),
    .B(_04457_),
    .C(_04458_),
    .X(_01864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11939_ (.A(\design_top.RAMFF[6] ),
    .Y(_01867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11940_ (.A(\design_top.IOMUX[3][6] ),
    .Y(_04485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11941_ (.A(\design_top.LEDFF[6] ),
    .Y(_04486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11942_ (.A1(_04485_),
    .A2(_04464_),
    .B1(_04486_),
    .B2(_04466_),
    .X(_01868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11943_ (.A(\design_top.RAMFF[22] ),
    .Y(_01870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11944_ (.A(\design_top.IOMUX[3][22] ),
    .Y(_04487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11945_ (.A(\design_top.GPIOFF[6] ),
    .Y(_04488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11946_ (.A1(_04487_),
    .A2(_06988_),
    .B1(_04488_),
    .B2(_06990_),
    .X(_01871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11947_ (.A(\design_top.RAMFF[30] ),
    .Y(_01876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11948_ (.A(\design_top.IOMUX[3][30] ),
    .Y(_04489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11949_ (.A(\design_top.GPIOFF[14] ),
    .Y(_04490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11950_ (.A1(_04489_),
    .A2(_06988_),
    .B1(_04490_),
    .B2(_06990_),
    .X(_01877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11951_ (.A(\design_top.RAMFF[14] ),
    .Y(_01879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11952_ (.A(\design_top.IOMUX[3][14] ),
    .Y(_04491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11953_ (.A(\design_top.LEDFF[14] ),
    .Y(_04492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _11954_ (.A1(\design_top.uart0.UART_RFIFO[6] ),
    .A2(_06991_),
    .B1(_01413_),
    .Y(_04493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11955_ (.A1(_04491_),
    .A2(_06981_),
    .B1(_04492_),
    .B2(_06985_),
    .C1(_04493_),
    .X(_01880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11956_ (.A1_N(_06862_),
    .A2_N(_06848_),
    .B1(_06862_),
    .B2(_06848_),
    .X(_02419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11957_ (.A(_02419_),
    .Y(_01888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11958_ (.A(\design_top.core0.NXPC[7] ),
    .Y(_01890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11959_ (.A1(_01846_),
    .A2(_04483_),
    .B1(_01845_),
    .Y(_04494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11960_ (.A1_N(_06571_),
    .A2_N(_04494_),
    .B1(_06571_),
    .B2(_04494_),
    .X(_01891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11961_ (.A1(_00786_),
    .A2(_00792_),
    .B1(_04641_),
    .B2(_04484_),
    .X(_04495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11962_ (.A(_04495_),
    .Y(_04496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11963_ (.A1(_00872_),
    .A2(_04495_),
    .B1(_06571_),
    .B2(_04496_),
    .X(_01892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11964_ (.A(_04456_),
    .B(_01397_),
    .X(_01893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11965_ (.A(_04443_),
    .B(_01893_),
    .X(_01894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11966_ (.A(_01902_),
    .B(_04457_),
    .C(_04458_),
    .X(_01903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11967_ (.A1(_05389_),
    .A2(\design_top.core0.PC[6] ),
    .B1(_06862_),
    .B2(_06848_),
    .X(_04497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11968_ (.A1_N(_06847_),
    .A2_N(_04497_),
    .B1(_06847_),
    .B2(_04497_),
    .X(_02423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11969_ (.A(_02423_),
    .Y(_01911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11970_ (.A(\design_top.core0.NXPC[8] ),
    .Y(_01913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11971_ (.A(_04635_),
    .X(_04498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11972_ (.A(_06947_),
    .Y(_04499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11973_ (.A1(_04498_),
    .A2(_04499_),
    .B1(_00873_),
    .B2(_06947_),
    .X(_01915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11974_ (.A1_N(_04498_),
    .A2_N(_06575_),
    .B1(_04498_),
    .B2(_06575_),
    .X(_01916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11975_ (.A(_04442_),
    .X(_04500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11976_ (.A(_04500_),
    .B(_01920_),
    .X(_01921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11977_ (.A(_04456_),
    .B(_01551_),
    .X(_01923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11978_ (.A(_01926_),
    .B(_04457_),
    .C(_04458_),
    .X(_01927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11979_ (.A(_06865_),
    .X(_04501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11980_ (.A1_N(_04501_),
    .A2_N(_06835_),
    .B1(_04501_),
    .B2(_06835_),
    .X(_02427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11981_ (.A(_02427_),
    .Y(_01935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11982_ (.A(\design_top.core0.NXPC[9] ),
    .Y(_01937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11983_ (.A(_04633_),
    .X(_04502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11984_ (.A1(_00873_),
    .A2(_06947_),
    .B1(_01914_),
    .Y(_04503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11985_ (.A1_N(_04502_),
    .A2_N(_04503_),
    .B1(_04502_),
    .B2(_04503_),
    .X(_01938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11986_ (.A1(_00775_),
    .A2(_00781_),
    .B1(_04498_),
    .B2(_06575_),
    .X(_04504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11987_ (.A1_N(_04502_),
    .A2_N(_04504_),
    .B1(_04502_),
    .B2(_04504_),
    .X(_01939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11988_ (.A(_04500_),
    .B(_01942_),
    .X(_01943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11989_ (.A(_04649_),
    .X(_04505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11990_ (.A(_04505_),
    .B(_01621_),
    .X(_01945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11991_ (.A(_06975_),
    .X(_04506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11992_ (.A(_06977_),
    .X(_04507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11993_ (.A(_01948_),
    .B(_04506_),
    .C(_04507_),
    .X(_01949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11994_ (.A1(_05386_),
    .A2(\design_top.core0.PC[8] ),
    .B1(_04501_),
    .B2(_06835_),
    .X(_04508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11995_ (.A1_N(_06834_),
    .A2_N(_04508_),
    .B1(_06834_),
    .B2(_04508_),
    .X(_02431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11996_ (.A(_02431_),
    .Y(_01957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11997_ (.A(\design_top.core0.NXPC[10] ),
    .Y(_01959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31oi_2 _11998_ (.A1(_04502_),
    .A2(_04498_),
    .A3(_04499_),
    .B1(_06948_),
    .Y(_04509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11999_ (.A1_N(_00875_),
    .A2_N(_04509_),
    .B1(_00875_),
    .B2(_04509_),
    .X(_01961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12000_ (.A1(_00772_),
    .A2(_01385_),
    .B1(_04633_),
    .B2(_04504_),
    .X(_04510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12001_ (.A1_N(_04638_),
    .A2_N(_04510_),
    .B1(_04638_),
    .B2(_04510_),
    .X(_01962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12002_ (.A(_04500_),
    .B(_01966_),
    .X(_01967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12003_ (.A(_04505_),
    .B(_01676_),
    .X(_01969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12004_ (.A(_01972_),
    .B(_04506_),
    .C(_04507_),
    .X(_01973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12005_ (.A(_06833_),
    .Y(_04511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31oi_2 _12006_ (.A1(_06834_),
    .A2(_06835_),
    .A3(_04501_),
    .B1(_06867_),
    .Y(_04512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12007_ (.A1_N(_04511_),
    .A2_N(_04512_),
    .B1(_04511_),
    .B2(_04512_),
    .X(_01981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12008_ (.A(\design_top.core0.NXPC[11] ),
    .Y(_01983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _12009_ (.A1(_00875_),
    .A2(_04509_),
    .B1(_01960_),
    .Y(_04513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12010_ (.A1_N(_04631_),
    .A2_N(_04513_),
    .B1(_04631_),
    .B2(_04513_),
    .X(_01984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12011_ (.A1(_00759_),
    .A2(_00765_),
    .B1(_04638_),
    .B2(_04510_),
    .X(_04514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12012_ (.A(_04514_),
    .Y(_04515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12013_ (.A1(_00876_),
    .A2(_04514_),
    .B1(_04631_),
    .B2(_04515_),
    .X(_01985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12014_ (.A(_04500_),
    .B(_01987_),
    .X(_01988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12015_ (.A(_04505_),
    .B(_01726_),
    .X(_01990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12016_ (.A(_01993_),
    .B(_04506_),
    .C(_04507_),
    .X(_01994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12017_ (.A1(_00507_),
    .A2(_06832_),
    .B1(_04511_),
    .B2(_04512_),
    .X(_04516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12018_ (.A1_N(_06830_),
    .A2_N(_04516_),
    .B1(_06830_),
    .B2(_04516_),
    .X(_02002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12019_ (.A(\design_top.core0.NXPC[12] ),
    .Y(_02004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _12020_ (.A1(_06947_),
    .A2(_06939_),
    .B1(_06950_),
    .Y(_04517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12021_ (.A(_04517_),
    .Y(_04518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12022_ (.A1(_04660_),
    .A2(_04517_),
    .B1(_00877_),
    .B2(_04518_),
    .X(_02006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12023_ (.A1_N(_06580_),
    .A2_N(_06733_),
    .B1(_06580_),
    .B2(_06733_),
    .X(_02007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12024_ (.A(_04500_),
    .B(_02011_),
    .X(_02012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12025_ (.A(_04505_),
    .B(_01770_),
    .X(_02014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12026_ (.A(_02017_),
    .B(_04506_),
    .C(_04507_),
    .X(_02018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _12027_ (.A1(_04501_),
    .A2(_06836_),
    .B1(_06869_),
    .Y(_04519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12028_ (.A(_04519_),
    .Y(_04520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12029_ (.A1(_06841_),
    .A2(_04519_),
    .B1(_06840_),
    .B2(_04520_),
    .X(_02443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12030_ (.A(_02443_),
    .Y(_02026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12031_ (.A(\design_top.core0.NXPC[13] ),
    .Y(_02028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _12032_ (.A1(_00877_),
    .A2(_04518_),
    .B1(_02005_),
    .Y(_04521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12033_ (.A1_N(_04657_),
    .A2_N(_04521_),
    .B1(_04657_),
    .B2(_04521_),
    .X(_02029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12034_ (.A1(_00743_),
    .A2(_00862_),
    .B1(_06580_),
    .B2(_06733_),
    .X(_04522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12035_ (.A1_N(_06732_),
    .A2_N(_04522_),
    .B1(_06732_),
    .B2(_04522_),
    .X(_02030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12036_ (.A(_06558_),
    .X(_04523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12037_ (.A(_04523_),
    .B(_02033_),
    .X(_02034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12038_ (.A(_04505_),
    .B(_01812_),
    .X(_02036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12039_ (.A(_02039_),
    .B(_04506_),
    .C(_04507_),
    .X(_02040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12040_ (.A1(_00495_),
    .A2(_06839_),
    .B1(_06841_),
    .B2(_04519_),
    .X(_04524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12041_ (.A1_N(_06838_),
    .A2_N(_04524_),
    .B1(_06838_),
    .B2(_04524_),
    .X(_02048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _12042_ (.A(_02049_),
    .B(_05604_),
    .Y(_02050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _12043_ (.A(\design_top.core0.RESMODE[0] ),
    .B(_07003_),
    .C(_00903_),
    .Y(_02051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12044_ (.A(\design_top.core0.NXPC[14] ),
    .Y(_02052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _12045_ (.A1(_00878_),
    .A2(_00877_),
    .A3(_04518_),
    .B1(_06951_),
    .X(_04525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12046_ (.A1_N(_02054_),
    .A2_N(_04525_),
    .B1(_02054_),
    .B2(_04525_),
    .X(_02055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _12047_ (.A1(_06732_),
    .A2(_06733_),
    .A3(_06580_),
    .B1(_06730_),
    .X(_04526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12048_ (.A1_N(_06726_),
    .A2_N(_04526_),
    .B1(_06726_),
    .B2(_04526_),
    .X(_02056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12049_ (.A(_04523_),
    .B(_02060_),
    .X(_02061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12050_ (.A(_04649_),
    .B(_01858_),
    .X(_02063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12051_ (.A(_06974_),
    .X(_04527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12052_ (.A(_06976_),
    .X(_04528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12053_ (.A(_02066_),
    .B(_04527_),
    .C(_04528_),
    .X(_02067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31oi_2 _12054_ (.A1(_06837_),
    .A2(_06840_),
    .A3(_04520_),
    .B1(_06871_),
    .Y(_04529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12055_ (.A1_N(_06843_),
    .A2_N(_04529_),
    .B1(_06843_),
    .B2(_04529_),
    .X(_02075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12056_ (.A(\design_top.core0.NXPC[15] ),
    .Y(_02077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _12057_ (.A1(_02054_),
    .A2(_04525_),
    .B1(_02053_),
    .Y(_04530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12058_ (.A1_N(_04666_),
    .A2_N(_04530_),
    .B1(_04666_),
    .B2(_04530_),
    .X(_02078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12059_ (.A1(_00726_),
    .A2(_00860_),
    .B1(_06726_),
    .B2(_04526_),
    .X(_04531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12060_ (.A1_N(_06725_),
    .A2_N(_04531_),
    .B1(_06725_),
    .B2(_04531_),
    .X(_02079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12061_ (.A(_04523_),
    .B(_01398_),
    .X(_02080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12062_ (.A(_02083_),
    .B(_04527_),
    .C(_04528_),
    .X(_02084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12063_ (.A1(_00483_),
    .A2(_06842_),
    .B1(_06843_),
    .B2(_04529_),
    .X(_04532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12064_ (.A1_N(_06845_),
    .A2_N(_04532_),
    .B1(_06845_),
    .B2(_04532_),
    .X(_02091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12065_ (.A(\design_top.core0.NXPC[16] ),
    .Y(_02093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12066_ (.A(_06954_),
    .Y(_04533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12067_ (.A1(_04683_),
    .A2(_04533_),
    .B1(_00880_),
    .B2(_06954_),
    .X(_02095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12068_ (.A1_N(_06735_),
    .A2_N(_06737_),
    .B1(_06735_),
    .B2(_06737_),
    .X(_02096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12069_ (.A(_04523_),
    .B(_01552_),
    .X(_02102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12070_ (.A(_02105_),
    .B(_04527_),
    .C(_04528_),
    .X(_02106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12071_ (.A(_06876_),
    .X(_04534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _12072_ (.A1_N(_04534_),
    .A2_N(_06817_),
    .B1(_04534_),
    .B2(_06817_),
    .X(_02459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12073_ (.A(_02459_),
    .Y(_02113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12074_ (.A(\design_top.core0.NXPC[17] ),
    .Y(_02115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _12075_ (.A1(_00880_),
    .A2(_06954_),
    .B1(_02094_),
    .Y(_04535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12076_ (.A1_N(_04679_),
    .A2_N(_04535_),
    .B1(_04679_),
    .B2(_04535_),
    .X(_02116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12077_ (.A1(_00714_),
    .A2(_00858_),
    .B1(_06735_),
    .B2(_06737_),
    .X(_04536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12078_ (.A1_N(_06736_),
    .A2_N(_04536_),
    .B1(_06736_),
    .B2(_04536_),
    .X(_02117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12079_ (.A(_04523_),
    .B(_01622_),
    .X(_02122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12080_ (.A(_02125_),
    .B(_04527_),
    .C(_04528_),
    .X(_02126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12081_ (.A1(_05414_),
    .A2(\design_top.core0.PC[16] ),
    .B1(_04534_),
    .B2(_06817_),
    .X(_04537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _12082_ (.A1_N(_06816_),
    .A2_N(_04537_),
    .B1(_06816_),
    .B2(_04537_),
    .X(_02463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12083_ (.A(_02463_),
    .Y(_02133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12084_ (.A(\design_top.core0.NXPC[18] ),
    .Y(_02135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31oi_2 _12085_ (.A1(_04679_),
    .A2(_04683_),
    .A3(_04533_),
    .B1(_06955_),
    .Y(_04538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12086_ (.A1_N(_02137_),
    .A2_N(_04538_),
    .B1(_02137_),
    .B2(_04538_),
    .X(_02138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _12087_ (.A1(_06736_),
    .A2(_06737_),
    .A3(_06735_),
    .B1(_06723_),
    .X(_04539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12088_ (.A1_N(_06718_),
    .A2_N(_04539_),
    .B1(_06718_),
    .B2(_04539_),
    .X(_02139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12089_ (.A(_06558_),
    .X(_04540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12090_ (.A(_04540_),
    .B(_01677_),
    .X(_02145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12091_ (.A(_02148_),
    .B(_04527_),
    .C(_04528_),
    .X(_02149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12092_ (.A(_06815_),
    .Y(_04541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31oi_2 _12093_ (.A1(_06816_),
    .A2(_06817_),
    .A3(_04534_),
    .B1(_06878_),
    .Y(_04542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12094_ (.A1_N(_04541_),
    .A2_N(_04542_),
    .B1(_04541_),
    .B2(_04542_),
    .X(_02156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12095_ (.A(\design_top.core0.NXPC[19] ),
    .Y(_02158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _12096_ (.A1(_02137_),
    .A2(_04538_),
    .B1(_02136_),
    .Y(_04543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12097_ (.A1_N(_04681_),
    .A2_N(_04543_),
    .B1(_04681_),
    .B2(_04543_),
    .X(_02159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12098_ (.A1(_00697_),
    .A2(_00856_),
    .B1(_06718_),
    .B2(_04539_),
    .X(_04544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12099_ (.A1_N(_06717_),
    .A2_N(_04544_),
    .B1(_06717_),
    .B2(_04544_),
    .X(_02160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12100_ (.A(_04540_),
    .B(_01727_),
    .X(_02164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12101_ (.A(_06974_),
    .X(_04545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12102_ (.A(_06976_),
    .X(_04546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12103_ (.A(_02167_),
    .B(_04545_),
    .C(_04546_),
    .X(_02168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12104_ (.A1(_00459_),
    .A2(_06814_),
    .B1(_04541_),
    .B2(_04542_),
    .X(_04547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12105_ (.A1_N(_06812_),
    .A2_N(_04547_),
    .B1(_06812_),
    .B2(_04547_),
    .X(_02175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12106_ (.A(\design_top.core0.NXPC[20] ),
    .Y(_02177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _12107_ (.A1(_06954_),
    .A2(_06937_),
    .B1(_06957_),
    .Y(_04548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12108_ (.A(_04548_),
    .Y(_04549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12109_ (.A1(_04695_),
    .A2(_04548_),
    .B1(_00883_),
    .B2(_04549_),
    .X(_02179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12110_ (.A1_N(_06713_),
    .A2_N(_06740_),
    .B1(_06713_),
    .B2(_06740_),
    .X(_02180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12111_ (.A(_04540_),
    .B(_01771_),
    .X(_02186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12112_ (.A(_02189_),
    .B(_04545_),
    .C(_04546_),
    .X(_02190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _12113_ (.A1(_04534_),
    .A2(_06818_),
    .B1(_06880_),
    .Y(_04550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12114_ (.A(_04550_),
    .Y(_04551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12115_ (.A1(_06823_),
    .A2(_04550_),
    .B1(_06822_),
    .B2(_04551_),
    .X(_02475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12116_ (.A(_02475_),
    .Y(_02197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12117_ (.A(\design_top.core0.NXPC[21] ),
    .Y(_02199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _12118_ (.A1(_00883_),
    .A2(_04549_),
    .B1(_02178_),
    .Y(_04552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12119_ (.A1_N(_04698_),
    .A2_N(_04552_),
    .B1(_04698_),
    .B2(_04552_),
    .X(_02200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12120_ (.A1(_00680_),
    .A2(_00854_),
    .B1(_06713_),
    .B2(_06740_),
    .X(_04553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12121_ (.A1_N(_06712_),
    .A2_N(_04553_),
    .B1(_06712_),
    .B2(_04553_),
    .X(_02201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12122_ (.A(_04540_),
    .B(_01813_),
    .X(_02206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12123_ (.A(_02209_),
    .B(_04545_),
    .C(_04546_),
    .X(_02210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12124_ (.A1(_00447_),
    .A2(_06821_),
    .B1(_06823_),
    .B2(_04550_),
    .X(_04554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12125_ (.A1_N(_06820_),
    .A2_N(_04554_),
    .B1(_06820_),
    .B2(_04554_),
    .X(_02217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12126_ (.A(\design_top.core0.NXPC[22] ),
    .Y(_02219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _12127_ (.A1(_00883_),
    .A2(_00884_),
    .A3(_04549_),
    .B1(_06958_),
    .X(_04555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12128_ (.A1_N(_00885_),
    .A2_N(_04555_),
    .B1(_00885_),
    .B2(_04555_),
    .X(_02221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _12129_ (.A1(_06712_),
    .A2(_06713_),
    .A3(_06740_),
    .B1(_06711_),
    .X(_04556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12130_ (.A1_N(_06706_),
    .A2_N(_04556_),
    .B1(_06706_),
    .B2(_04556_),
    .X(_02222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12131_ (.A(_04540_),
    .B(_01859_),
    .X(_02228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12132_ (.A(_02231_),
    .B(_04545_),
    .C(_04546_),
    .X(_02232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31oi_2 _12133_ (.A1(_06819_),
    .A2(_06822_),
    .A3(_04551_),
    .B1(_06882_),
    .Y(_04557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12134_ (.A1_N(_06825_),
    .A2_N(_04557_),
    .B1(_06825_),
    .B2(_04557_),
    .X(_02239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12135_ (.A(\design_top.core0.NXPC[23] ),
    .Y(_02241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _12136_ (.A1(_00885_),
    .A2(_04555_),
    .B1(_02220_),
    .Y(_04558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12137_ (.A1_N(_04692_),
    .A2_N(_04558_),
    .B1(_04692_),
    .B2(_04558_),
    .X(_02242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12138_ (.A1(_00663_),
    .A2(_00852_),
    .B1(_06706_),
    .B2(_04556_),
    .X(_04559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12139_ (.A1_N(_06705_),
    .A2_N(_04559_),
    .B1(_06705_),
    .B2(_04559_),
    .X(_02243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12140_ (.A(_06558_),
    .X(_04560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12141_ (.A(_04560_),
    .B(_01899_),
    .X(_02246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12142_ (.A(_02249_),
    .B(_04545_),
    .C(_04546_),
    .X(_02250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12143_ (.A1(_00435_),
    .A2(_06824_),
    .B1(_06825_),
    .B2(_04557_),
    .X(_04561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12144_ (.A1_N(_06827_),
    .A2_N(_04561_),
    .B1(_06827_),
    .B2(_04561_),
    .X(_02257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _12145_ (.A(_06908_),
    .B(_00534_),
    .Y(_00536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12146_ (.A(\design_top.core0.NXPC[24] ),
    .Y(_02259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12147_ (.A1_N(_00887_),
    .A2_N(_06961_),
    .B1(_00887_),
    .B2(_06961_),
    .X(_02261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12148_ (.A1_N(_06702_),
    .A2_N(_06742_),
    .B1(_06702_),
    .B2(_06742_),
    .X(_02262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12149_ (.A(_04560_),
    .B(_01923_),
    .X(_02268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12150_ (.A(_06974_),
    .X(_04562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12151_ (.A(_06976_),
    .X(_04563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12152_ (.A(_02271_),
    .B(_04562_),
    .C(_04563_),
    .X(_02272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12153_ (.A1(_06888_),
    .A2(_06810_),
    .B1(_06887_),
    .B2(_06809_),
    .X(_02491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12154_ (.A(_02491_),
    .Y(_02279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12155_ (.A(\design_top.core0.NXPC[25] ),
    .Y(_02281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _12156_ (.A1(_00887_),
    .A2(_06961_),
    .B1(_02260_),
    .Y(_04564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12157_ (.A1_N(_04673_),
    .A2_N(_04564_),
    .B1(_04673_),
    .B2(_04564_),
    .X(_02282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12158_ (.A1(_00646_),
    .A2(_00850_),
    .B1(_06702_),
    .B2(_06742_),
    .X(_04565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12159_ (.A1_N(_06701_),
    .A2_N(_04565_),
    .B1(_06701_),
    .B2(_04565_),
    .X(_02283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12160_ (.A(_04560_),
    .B(_01945_),
    .X(_02288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12161_ (.A(_02291_),
    .B(_04562_),
    .C(_04563_),
    .X(_02292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12162_ (.A1(_05405_),
    .A2(\design_top.core0.PC[24] ),
    .B1(_06887_),
    .B2(_06809_),
    .X(_04566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _12163_ (.A1_N(_06807_),
    .A2_N(_04566_),
    .B1(_06807_),
    .B2(_04566_),
    .X(_02495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12164_ (.A(_02495_),
    .Y(_02299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12165_ (.A(\design_top.core0.NXPC[26] ),
    .Y(_02301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _12166_ (.A1(_00887_),
    .A2(_00888_),
    .A3(_06961_),
    .B1(_06963_),
    .X(_04567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12167_ (.A1_N(_00889_),
    .A2_N(_04567_),
    .B1(_00889_),
    .B2(_04567_),
    .X(_02303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _12168_ (.A1(_06701_),
    .A2(_06702_),
    .A3(_06742_),
    .B1(_06699_),
    .X(_04568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12169_ (.A1_N(_06695_),
    .A2_N(_04568_),
    .B1(_06695_),
    .B2(_04568_),
    .X(_02304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12170_ (.A(_04560_),
    .B(_01969_),
    .X(_02310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12171_ (.A(_02313_),
    .B(_04562_),
    .C(_04563_),
    .X(_02314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _12172_ (.A1(_06808_),
    .A2(_06810_),
    .A3(_06888_),
    .B1(_06805_),
    .X(_04569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12173_ (.A1_N(_06802_),
    .A2_N(_04569_),
    .B1(_06802_),
    .B2(_04569_),
    .X(_02321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12174_ (.A(\design_top.core0.NXPC[27] ),
    .Y(_02323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _12175_ (.A1(_00889_),
    .A2(_04567_),
    .B1(_02302_),
    .Y(_04570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12176_ (.A1_N(_04669_),
    .A2_N(_04570_),
    .B1(_04669_),
    .B2(_04570_),
    .X(_02324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12177_ (.A1(_00629_),
    .A2(_00848_),
    .B1(_06695_),
    .B2(_04568_),
    .X(_04571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12178_ (.A1_N(_06694_),
    .A2_N(_04571_),
    .B1(_06694_),
    .B2(_04571_),
    .X(_02325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12179_ (.A(_04560_),
    .B(_01990_),
    .X(_02329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12180_ (.A(_02332_),
    .B(_04562_),
    .C(_04563_),
    .X(_02333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12181_ (.A1(_00411_),
    .A2(_06799_),
    .B1(_06802_),
    .B2(_04569_),
    .X(_04572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12182_ (.A1_N(_06801_),
    .A2_N(_04572_),
    .B1(_06801_),
    .B2(_04572_),
    .X(_02340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12183_ (.A(\design_top.core0.NXPC[28] ),
    .Y(_02342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12184_ (.A1_N(_00891_),
    .A2_N(_06965_),
    .B1(_00891_),
    .B2(_06965_),
    .X(_02344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12185_ (.A1(_06745_),
    .A2(_06687_),
    .B1(_06744_),
    .B2(_06686_),
    .X(_02345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12186_ (.A(_04442_),
    .B(_02014_),
    .X(_02351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12187_ (.A(_02354_),
    .B(_04562_),
    .C(_04563_),
    .X(_02355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _12188_ (.A1(_04729_),
    .A2(\design_top.core0.PC[28] ),
    .B1(_06797_),
    .X(_04573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _12189_ (.A1_N(_06890_),
    .A2_N(_04573_),
    .B1(_06890_),
    .B2(_04573_),
    .X(_02507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12190_ (.A(_02507_),
    .Y(_02362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12191_ (.A(\design_top.core0.NXPC[29] ),
    .Y(_02364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12192_ (.A1(_00892_),
    .A2(_06967_),
    .B1(_04705_),
    .B2(_06966_),
    .X(_02365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12193_ (.A1(_00612_),
    .A2(_00846_),
    .B1(_06744_),
    .B2(_06686_),
    .X(_04574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12194_ (.A1_N(_06970_),
    .A2_N(_04574_),
    .B1(_06970_),
    .B2(_04574_),
    .X(_02366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12195_ (.A(_04442_),
    .B(_02036_),
    .X(_02371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12196_ (.A(_02374_),
    .B(_06975_),
    .C(_06977_),
    .X(_02375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12197_ (.A(\design_top.core0.NXPC[30] ),
    .Y(_02383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12198_ (.A1_N(_00893_),
    .A2_N(_06968_),
    .B1(_00893_),
    .B2(_06968_),
    .X(_02384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12199_ (.A1_N(_06690_),
    .A2_N(_06971_),
    .B1(_06690_),
    .B2(_06971_),
    .X(_02385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12200_ (.A(_04442_),
    .B(_02063_),
    .X(_02391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _12201_ (.A(_02394_),
    .B(_06975_),
    .C(_06977_),
    .X(_02395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12202_ (.A(io_out[18]),
    .Y(_02405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12203_ (.A(_01707_),
    .Y(_02406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12204_ (.A1(io_out[19]),
    .A2(io_out[18]),
    .B1(_06759_),
    .X(_02408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _12205_ (.A1_N(_05469_),
    .A2_N(_06760_),
    .B1(_05469_),
    .B2(_06760_),
    .X(_02411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _12206_ (.A1(_05469_),
    .A2(_06760_),
    .B1(\design_top.IADDR[5] ),
    .Y(_04575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _12207_ (.A(_06761_),
    .B(_04575_),
    .Y(_02414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12208_ (.A1(\design_top.IADDR[6] ),
    .A2(_06761_),
    .B1(_06762_),
    .X(_02418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _12209_ (.A1(_04803_),
    .A2(_04805_),
    .A3(_04827_),
    .B1(_04829_),
    .X(_04576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _12210_ (.A1_N(_04809_),
    .A2_N(_04576_),
    .B1(_04809_),
    .B2(_04576_),
    .Y(_02420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12211_ (.A1(\design_top.IADDR[7] ),
    .A2(_06763_),
    .B1(_06764_),
    .X(_02422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12212_ (.A1(_00531_),
    .A2(_00786_),
    .B1(_04809_),
    .B2(_04576_),
    .X(_04577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _12213_ (.A1_N(_04807_),
    .A2_N(_04577_),
    .B1(_04807_),
    .B2(_04577_),
    .Y(_02424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12214_ (.A1(\design_top.IADDR[8] ),
    .A2(_06765_),
    .B1(_06766_),
    .X(_02426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12215_ (.A(_04832_),
    .X(_04578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12216_ (.A(_04578_),
    .Y(_04579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12217_ (.A1(_04578_),
    .A2(_04836_),
    .B1(_04579_),
    .B2(_04835_),
    .X(_02428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12218_ (.A1(\design_top.IADDR[9] ),
    .A2(_06767_),
    .B1(_06768_),
    .X(_02430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12219_ (.A1(_00519_),
    .A2(_00775_),
    .B1(_04578_),
    .B2(_04836_),
    .X(_04580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12220_ (.A(_04580_),
    .Y(_04581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12221_ (.A1(_04834_),
    .A2(_04580_),
    .B1(_04833_),
    .B2(_04581_),
    .X(_02432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12222_ (.A1(\design_top.IADDR[10] ),
    .A2(_06769_),
    .B1(_06770_),
    .X(_02434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12223_ (.A(_01981_),
    .Y(_02435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _12224_ (.A1(_04834_),
    .A2(_04836_),
    .A3(_04578_),
    .B1(_04798_),
    .X(_04582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12225_ (.A(_04582_),
    .Y(_04583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12226_ (.A1(_04793_),
    .A2(_04582_),
    .B1(_04792_),
    .B2(_04583_),
    .X(_02436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12227_ (.A1(\design_top.IADDR[11] ),
    .A2(_06771_),
    .B1(_06772_),
    .X(_02438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12228_ (.A(_02002_),
    .Y(_02439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12229_ (.A1(_00507_),
    .A2(_00759_),
    .B1(_04793_),
    .B2(_04582_),
    .X(_04584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12230_ (.A(_04584_),
    .Y(_04585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12231_ (.A1(_04796_),
    .A2(_04584_),
    .B1(_04795_),
    .B2(_04585_),
    .X(_02440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12232_ (.A1(\design_top.IADDR[12] ),
    .A2(_06773_),
    .B1(_06774_),
    .X(_02442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _12233_ (.A1(_04578_),
    .A2(_04837_),
    .B1(_04801_),
    .Y(_04586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12234_ (.A(_04586_),
    .Y(_04587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12235_ (.A1(_04788_),
    .A2(_04587_),
    .B1(_04787_),
    .B2(_04586_),
    .X(_02444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12236_ (.A1(\design_top.IADDR[13] ),
    .A2(_06775_),
    .B1(_06776_),
    .X(_02446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12237_ (.A(_02048_),
    .Y(_02447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12238_ (.A1(_00495_),
    .A2(_00743_),
    .B1(_04788_),
    .B2(_04587_),
    .X(_04588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12239_ (.A(_04588_),
    .Y(_04589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12240_ (.A1(_04784_),
    .A2(_04588_),
    .B1(_04783_),
    .B2(_04589_),
    .X(_02448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12241_ (.A1(\design_top.IADDR[14] ),
    .A2(_06777_),
    .B1(_06778_),
    .X(_02450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12242_ (.A(_02075_),
    .Y(_02451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _12243_ (.A1(_04784_),
    .A2(_04788_),
    .A3(_04587_),
    .B1(_04840_),
    .X(_04590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12244_ (.A(_04590_),
    .Y(_04591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12245_ (.A1(_04778_),
    .A2(_04590_),
    .B1(_04777_),
    .B2(_04591_),
    .X(_02452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12246_ (.A1(\design_top.IADDR[15] ),
    .A2(_06779_),
    .B1(_06780_),
    .X(_02454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12247_ (.A(_02091_),
    .Y(_02455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12248_ (.A1(_00483_),
    .A2(_00726_),
    .B1(_04778_),
    .B2(_04590_),
    .X(_04592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12249_ (.A(_04592_),
    .Y(_04593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12250_ (.A1(_04781_),
    .A2(_04592_),
    .B1(_04780_),
    .B2(_04593_),
    .X(_02456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _12251_ (.A(_06781_),
    .B(_06780_),
    .Y(_04594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _12252_ (.A1(_06781_),
    .A2(_06780_),
    .B1(_04594_),
    .Y(_02458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12253_ (.A(_04845_),
    .X(_04595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _12254_ (.A1_N(_04595_),
    .A2_N(_04759_),
    .B1(_04595_),
    .B2(_04759_),
    .X(_02460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12255_ (.A1(\design_top.IADDR[17] ),
    .A2(_04594_),
    .B1(_06782_),
    .X(_02462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12256_ (.A1(_05414_),
    .A2(_04682_),
    .B1(_04595_),
    .B2(_04759_),
    .X(_04596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _12257_ (.A1_N(_04757_),
    .A2_N(_04596_),
    .B1(_04757_),
    .B2(_04596_),
    .X(_02464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12258_ (.A(\design_top.IADDR[18] ),
    .Y(_04597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _12259_ (.A(_04597_),
    .B(_06782_),
    .Y(_04598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _12260_ (.A1(_04597_),
    .A2(_06782_),
    .B1(_04598_),
    .Y(_02466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12261_ (.A(_02156_),
    .Y(_02467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _12262_ (.A1(_04757_),
    .A2(_04759_),
    .A3(_04595_),
    .B1(_04848_),
    .X(_04599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _12263_ (.A1_N(_04752_),
    .A2_N(_04599_),
    .B1(_04752_),
    .B2(_04599_),
    .X(_02468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ba_2 _12264_ (.A1(\design_top.IADDR[19] ),
    .A2(_04598_),
    .B1_N(_06783_),
    .X(_02470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12265_ (.A(_02175_),
    .Y(_02471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12266_ (.A1(_04751_),
    .A2(_00458_),
    .B1(_04752_),
    .B2(_04599_),
    .X(_04600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _12267_ (.A1_N(_04755_),
    .A2_N(_04600_),
    .B1(_04755_),
    .B2(_04600_),
    .X(_02472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12268_ (.A1(\design_top.IADDR[20] ),
    .A2(_06783_),
    .B1(_06784_),
    .X(_02474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _12269_ (.A1(_04595_),
    .A2(_04760_),
    .B1(_04852_),
    .Y(_04601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12270_ (.A(_04601_),
    .Y(_04602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12271_ (.A1(_04767_),
    .A2(_04601_),
    .B1(_04766_),
    .B2(_04602_),
    .X(_02476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12272_ (.A1(\design_top.IADDR[21] ),
    .A2(_06785_),
    .B1(_06786_),
    .X(_02478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12273_ (.A(_02217_),
    .Y(_02479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12274_ (.A1(_00447_),
    .A2(_00680_),
    .B1(_04767_),
    .B2(_04601_),
    .X(_04603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12275_ (.A(_04603_),
    .Y(_04604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12276_ (.A1(_04763_),
    .A2(_04603_),
    .B1(_04762_),
    .B2(_04604_),
    .X(_02480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12277_ (.A1(\design_top.IADDR[22] ),
    .A2(_06787_),
    .B1(_06788_),
    .X(_02482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12278_ (.A(_02239_),
    .Y(_02483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31oi_2 _12279_ (.A1(_04762_),
    .A2(_04766_),
    .A3(_04602_),
    .B1(_04854_),
    .Y(_04605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _12280_ (.A1_N(_04770_),
    .A2_N(_04605_),
    .B1(_04770_),
    .B2(_04605_),
    .Y(_02484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12281_ (.A1(\design_top.IADDR[23] ),
    .A2(_06789_),
    .B1(_06790_),
    .X(_02486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12282_ (.A(_02257_),
    .Y(_02487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12283_ (.A1(_00435_),
    .A2(_00663_),
    .B1(_04770_),
    .B2(_04605_),
    .X(_04606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _12284_ (.A1_N(_04772_),
    .A2_N(_04606_),
    .B1(_04772_),
    .B2(_04606_),
    .Y(_02488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _12285_ (.A(_06791_),
    .B(_06790_),
    .Y(_04607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _12286_ (.A1(_06791_),
    .A2(_06790_),
    .B1(_04607_),
    .Y(_02490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12287_ (.A1(_04860_),
    .A2(_04748_),
    .B1(_04859_),
    .B2(_04747_),
    .X(_02492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12288_ (.A1(\design_top.IADDR[25] ),
    .A2(_04607_),
    .B1(_06792_),
    .X(_02494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12289_ (.A1(_05405_),
    .A2(_04674_),
    .B1(_04859_),
    .B2(_04747_),
    .X(_04608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _12290_ (.A1_N(_04744_),
    .A2_N(_04608_),
    .B1(_04744_),
    .B2(_04608_),
    .X(_02496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12291_ (.A(\design_top.IADDR[26] ),
    .Y(_04609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _12292_ (.A(_04609_),
    .B(_06792_),
    .Y(_04610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _12293_ (.A1(_04609_),
    .A2(_06792_),
    .B1(_04610_),
    .Y(_02498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12294_ (.A(_02321_),
    .Y(_02499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _12295_ (.A1(_04745_),
    .A2(_04748_),
    .A3(_04860_),
    .B1(_04741_),
    .X(_04611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _12296_ (.A1_N(_04738_),
    .A2_N(_04611_),
    .B1(_04738_),
    .B2(_04611_),
    .Y(_02500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ba_2 _12297_ (.A1(\design_top.IADDR[27] ),
    .A2(_04610_),
    .B1_N(_06793_),
    .X(_02502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12298_ (.A(_02340_),
    .Y(_02503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12299_ (.A1(_00411_),
    .A2(_00629_),
    .B1(_04738_),
    .B2(_04611_),
    .X(_04612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _12300_ (.A1_N(_04737_),
    .A2_N(_04612_),
    .B1(_04737_),
    .B2(_04612_),
    .Y(_02504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12301_ (.A1(\design_top.IADDR[28] ),
    .A2(_06793_),
    .B1(_06794_),
    .X(_02506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12302_ (.A(_04862_),
    .Y(_04613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12303_ (.A1(_04862_),
    .A2(_04731_),
    .B1(_04613_),
    .B2(_04730_),
    .X(_02508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2b_2 _12304_ (.A_N(\design_top.uart0.UART_RXDFF[1] ),
    .B(_06518_),
    .Y(_02512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12305_ (.A(_02404_),
    .Y(_04614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _12306_ (.A1(io_out[17]),
    .A2(_04713_),
    .B1(_04614_),
    .B2(_04712_),
    .C1(_05426_),
    .X(_04437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12307_ (.LO(io_oeb[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12308_ (.LO(io_oeb[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12309_ (.LO(io_oeb[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12310_ (.LO(io_oeb[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12311_ (.LO(io_oeb[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12312_ (.LO(io_oeb[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12313_ (.LO(io_oeb[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12314_ (.LO(io_oeb[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12315_ (.LO(io_oeb[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12316_ (.LO(io_oeb[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12317_ (.LO(io_oeb[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12318_ (.LO(io_oeb[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12319_ (.LO(io_oeb[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12320_ (.LO(io_oeb[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12321_ (.LO(io_oeb[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12322_ (.LO(io_oeb[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12323_ (.LO(io_oeb[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12324_ (.LO(io_oeb[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12325_ (.LO(io_oeb[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12326_ (.LO(io_oeb[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12327_ (.LO(io_oeb[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12328_ (.LO(io_oeb[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12329_ (.LO(io_oeb[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12330_ (.LO(io_oeb[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12331_ (.LO(io_oeb[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12332_ (.LO(io_oeb[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12333_ (.LO(io_oeb[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12334_ (.LO(io_oeb[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12335_ (.LO(io_oeb[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12336_ (.LO(io_oeb[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12337_ (.LO(io_oeb[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12338_ (.LO(io_oeb[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12339_ (.LO(io_oeb[32]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12340_ (.LO(io_oeb[33]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12341_ (.LO(io_oeb[34]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12342_ (.LO(io_oeb[35]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12343_ (.LO(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12344_ (.LO(io_oeb[37]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12345_ (.LO(io_out[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12346_ (.LO(io_out[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12347_ (.LO(io_out[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12348_ (.LO(io_out[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12349_ (.LO(io_out[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12350_ (.LO(io_out[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12351_ (.LO(io_out[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12352_ (.LO(io_out[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12353_ (.LO(io_out[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12354_ (.LO(io_out[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12355_ (.LO(io_out[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12356_ (.LO(io_out[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12357_ (.LO(io_out[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12358_ (.LO(io_out[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12359_ (.LO(io_out[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12360_ (.LO(io_out[32]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12361_ (.LO(io_out[33]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12362_ (.LO(io_out[34]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12363_ (.LO(io_out[35]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12364_ (.LO(io_out[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12365_ (.LO(io_out[37]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12366_ (.LO(la_data_out[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12367_ (.LO(la_data_out[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12368_ (.LO(la_data_out[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12369_ (.LO(la_data_out[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12370_ (.LO(la_data_out[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12371_ (.LO(la_data_out[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12372_ (.LO(la_data_out[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12373_ (.LO(la_data_out[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12374_ (.LO(la_data_out[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12375_ (.LO(la_data_out[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12376_ (.LO(la_data_out[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12377_ (.LO(la_data_out[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12378_ (.LO(la_data_out[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12379_ (.LO(la_data_out[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12380_ (.LO(la_data_out[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12381_ (.LO(la_data_out[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12382_ (.LO(la_data_out[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12383_ (.LO(la_data_out[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12384_ (.LO(la_data_out[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12385_ (.LO(la_data_out[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12386_ (.LO(la_data_out[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12387_ (.LO(la_data_out[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12388_ (.LO(la_data_out[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12389_ (.LO(la_data_out[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12390_ (.LO(la_data_out[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12391_ (.LO(la_data_out[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12392_ (.LO(la_data_out[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12393_ (.LO(la_data_out[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12394_ (.LO(la_data_out[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12395_ (.LO(la_data_out[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12396_ (.LO(la_data_out[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12397_ (.LO(la_data_out[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12398_ (.LO(la_data_out[32]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12399_ (.LO(la_data_out[33]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12400_ (.LO(la_data_out[34]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12401_ (.LO(la_data_out[35]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12402_ (.LO(la_data_out[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12403_ (.LO(la_data_out[37]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12404_ (.LO(la_data_out[38]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12405_ (.LO(la_data_out[39]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12406_ (.LO(la_data_out[40]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12407_ (.LO(la_data_out[41]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12408_ (.LO(la_data_out[42]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12409_ (.LO(la_data_out[43]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12410_ (.LO(la_data_out[44]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12411_ (.LO(la_data_out[45]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12412_ (.LO(la_data_out[46]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12413_ (.LO(la_data_out[47]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12414_ (.LO(la_data_out[48]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12415_ (.LO(la_data_out[49]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12416_ (.LO(la_data_out[50]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12417_ (.LO(la_data_out[51]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12418_ (.LO(la_data_out[52]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12419_ (.LO(la_data_out[53]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12420_ (.LO(la_data_out[54]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12421_ (.LO(la_data_out[55]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12422_ (.LO(la_data_out[56]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12423_ (.LO(la_data_out[57]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12424_ (.LO(la_data_out[58]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12425_ (.LO(la_data_out[59]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12426_ (.LO(la_data_out[60]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12427_ (.LO(la_data_out[61]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12428_ (.LO(la_data_out[62]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12429_ (.LO(la_data_out[63]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12430_ (.LO(la_data_out[64]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12431_ (.LO(la_data_out[65]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12432_ (.LO(la_data_out[66]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12433_ (.LO(la_data_out[67]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12434_ (.LO(la_data_out[68]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12435_ (.LO(la_data_out[69]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12436_ (.LO(la_data_out[70]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12437_ (.LO(la_data_out[71]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12438_ (.LO(la_data_out[72]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12439_ (.LO(la_data_out[73]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12440_ (.LO(la_data_out[74]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12441_ (.LO(la_data_out[75]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12442_ (.LO(la_data_out[76]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12443_ (.LO(la_data_out[77]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12444_ (.LO(la_data_out[78]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12445_ (.LO(la_data_out[79]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12446_ (.LO(la_data_out[80]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12447_ (.LO(la_data_out[81]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12448_ (.LO(la_data_out[82]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12449_ (.LO(la_data_out[83]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12450_ (.LO(la_data_out[84]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12451_ (.LO(la_data_out[85]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12452_ (.LO(la_data_out[86]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12453_ (.LO(la_data_out[87]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12454_ (.LO(la_data_out[88]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12455_ (.LO(la_data_out[89]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12456_ (.LO(la_data_out[90]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12457_ (.LO(la_data_out[91]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12458_ (.LO(la_data_out[92]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12459_ (.LO(la_data_out[93]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12460_ (.LO(la_data_out[94]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12461_ (.LO(la_data_out[95]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12462_ (.LO(la_data_out[96]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12463_ (.LO(la_data_out[97]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12464_ (.LO(la_data_out[98]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12465_ (.LO(la_data_out[99]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12466_ (.LO(la_data_out[100]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12467_ (.LO(la_data_out[101]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12468_ (.LO(la_data_out[102]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12469_ (.LO(la_data_out[103]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12470_ (.LO(la_data_out[104]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12471_ (.LO(la_data_out[105]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12472_ (.LO(la_data_out[106]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12473_ (.LO(la_data_out[107]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12474_ (.LO(la_data_out[108]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12475_ (.LO(la_data_out[109]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12476_ (.LO(la_data_out[110]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12477_ (.LO(la_data_out[111]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12478_ (.LO(la_data_out[112]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12479_ (.LO(la_data_out[113]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12480_ (.LO(la_data_out[114]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12481_ (.LO(la_data_out[115]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12482_ (.LO(la_data_out[116]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12483_ (.LO(la_data_out[117]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12484_ (.LO(la_data_out[118]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12485_ (.LO(la_data_out[119]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12486_ (.LO(la_data_out[120]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12487_ (.LO(la_data_out[121]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12488_ (.LO(la_data_out[122]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12489_ (.LO(la_data_out[123]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12490_ (.LO(la_data_out[124]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12491_ (.LO(la_data_out[125]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12492_ (.LO(la_data_out[126]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12493_ (.LO(la_data_out[127]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12494_ (.LO(user_irq[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12495_ (.LO(user_irq[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12496_ (.LO(user_irq[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12497_ (.LO(wbs_ack_o),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12498_ (.LO(wbs_dat_o[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12499_ (.LO(wbs_dat_o[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12500_ (.LO(wbs_dat_o[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12501_ (.LO(wbs_dat_o[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12502_ (.LO(wbs_dat_o[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12503_ (.LO(wbs_dat_o[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12504_ (.LO(wbs_dat_o[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12505_ (.LO(wbs_dat_o[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12506_ (.LO(wbs_dat_o[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12507_ (.LO(wbs_dat_o[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12508_ (.LO(wbs_dat_o[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12509_ (.LO(wbs_dat_o[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12510_ (.LO(wbs_dat_o[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12511_ (.LO(wbs_dat_o[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12512_ (.LO(wbs_dat_o[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12513_ (.LO(wbs_dat_o[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12514_ (.LO(wbs_dat_o[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12515_ (.LO(wbs_dat_o[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12516_ (.LO(wbs_dat_o[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12517_ (.LO(wbs_dat_o[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12518_ (.LO(wbs_dat_o[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12519_ (.LO(wbs_dat_o[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12520_ (.LO(wbs_dat_o[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12521_ (.LO(wbs_dat_o[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12522_ (.LO(wbs_dat_o[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12523_ (.LO(wbs_dat_o[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12524_ (.LO(wbs_dat_o[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12525_ (.LO(wbs_dat_o[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12526_ (.LO(wbs_dat_o[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12527_ (.LO(wbs_dat_o[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12528_ (.LO(wbs_dat_o[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _12529_ (.LO(wbs_dat_o[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _12530_ (.A(io_out[15]),
    .X(\design_top.GPIOFF[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _12531_ (.A(io_out[8]),
    .X(\design_top.LEDFF[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _12532_ (.A(io_out[9]),
    .X(\design_top.LEDFF[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _12533_ (.A(io_out[10]),
    .X(\design_top.LEDFF[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _12534_ (.A(io_out[11]),
    .X(\design_top.LEDFF[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _12535_ (.A(io_out[14]),
    .X(\design_top.XTIMER ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12536_ (.A0(_00866_),
    .A1(_00539_),
    .S(io_out[12]),
    .X(_07035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12537_ (.A0(_00532_),
    .A1(_01363_),
    .S(_00537_),
    .X(_07036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12538_ (.A0(\design_top.ROMFF[0] ),
    .A1(\design_top.ROMFF2[0] ),
    .S(\design_top.HLT2 ),
    .X(io_out[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12539_ (.A0(\design_top.ROMFF[1] ),
    .A1(\design_top.ROMFF2[1] ),
    .S(\design_top.HLT2 ),
    .X(io_out[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12540_ (.A0(\design_top.ROMFF[2] ),
    .A1(\design_top.ROMFF2[2] ),
    .S(\design_top.HLT2 ),
    .X(io_out[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12541_ (.A0(\design_top.ROMFF[3] ),
    .A1(\design_top.ROMFF2[3] ),
    .S(\design_top.HLT2 ),
    .X(io_out[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12542_ (.A0(_00839_),
    .A1(_01056_),
    .S(_00532_),
    .X(_01057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12543_ (.A0(_01057_),
    .A1(_01055_),
    .S(_00537_),
    .X(\design_top.DATAO[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12544_ (.A0(_00832_),
    .A1(_01059_),
    .S(_00532_),
    .X(_01060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12545_ (.A0(_01060_),
    .A1(_01058_),
    .S(_00537_),
    .X(\design_top.DATAO[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12546_ (.A0(_00824_),
    .A1(_01062_),
    .S(_00532_),
    .X(_01063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12547_ (.A0(_01063_),
    .A1(_01061_),
    .S(_00537_),
    .X(\design_top.DATAO[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12548_ (.A0(_00815_),
    .A1(_01065_),
    .S(_00532_),
    .X(_01066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12549_ (.A0(_01066_),
    .A1(_01064_),
    .S(_00537_),
    .X(\design_top.DATAO[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12550_ (.A0(_00807_),
    .A1(_01068_),
    .S(_00532_),
    .X(_01069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12551_ (.A0(_01069_),
    .A1(_01067_),
    .S(_00537_),
    .X(\design_top.DATAO[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12552_ (.A0(_00798_),
    .A1(_01071_),
    .S(_00532_),
    .X(_01072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12553_ (.A0(_01072_),
    .A1(_01070_),
    .S(_00537_),
    .X(\design_top.DATAO[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12554_ (.A0(_00791_),
    .A1(_01074_),
    .S(_00532_),
    .X(_01075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12555_ (.A0(_01075_),
    .A1(_01073_),
    .S(_00537_),
    .X(\design_top.DATAO[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12556_ (.A0(_00570_),
    .A1(_01077_),
    .S(_00532_),
    .X(_01078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12557_ (.A0(_01078_),
    .A1(_01076_),
    .S(_00537_),
    .X(\design_top.DATAO[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12558_ (.A0(_00780_),
    .A1(_01444_),
    .S(_00532_),
    .X(_01445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12559_ (.A0(_01445_),
    .A1(_01443_),
    .S(_00537_),
    .X(\design_top.DATAO[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12560_ (.A0(_00771_),
    .A1(_01447_),
    .S(_00532_),
    .X(_01448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12561_ (.A0(_01448_),
    .A1(_01446_),
    .S(_00537_),
    .X(\design_top.DATAO[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12562_ (.A0(_00764_),
    .A1(_01450_),
    .S(_00532_),
    .X(_01451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12563_ (.A0(_01451_),
    .A1(_01449_),
    .S(_00537_),
    .X(\design_top.DATAO[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12564_ (.A0(_00755_),
    .A1(_01453_),
    .S(_00532_),
    .X(_01454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12565_ (.A0(_01454_),
    .A1(_01452_),
    .S(_00537_),
    .X(\design_top.DATAO[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12566_ (.A0(_00748_),
    .A1(_01456_),
    .S(_00532_),
    .X(_01457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12567_ (.A0(_01457_),
    .A1(_01455_),
    .S(_00537_),
    .X(\design_top.DATAO[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12568_ (.A0(_00739_),
    .A1(_01459_),
    .S(_00532_),
    .X(_01460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12569_ (.A0(_01460_),
    .A1(_01458_),
    .S(_00537_),
    .X(\design_top.DATAO[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12570_ (.A0(_00731_),
    .A1(_01462_),
    .S(_00532_),
    .X(_01463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12571_ (.A0(_01463_),
    .A1(_01461_),
    .S(_00537_),
    .X(\design_top.DATAO[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12572_ (.A0(_00576_),
    .A1(_01465_),
    .S(_00532_),
    .X(_01466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12573_ (.A0(_01466_),
    .A1(_01464_),
    .S(_00537_),
    .X(\design_top.DATAO[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12574_ (.A0(_00719_),
    .A1(_01468_),
    .S(_00532_),
    .X(_01469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12575_ (.A0(_01469_),
    .A1(_01467_),
    .S(_00537_),
    .X(\design_top.DATAO[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12576_ (.A0(_00710_),
    .A1(_01471_),
    .S(_00532_),
    .X(_01472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12577_ (.A0(_01472_),
    .A1(_01470_),
    .S(_00537_),
    .X(\design_top.DATAO[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12578_ (.A0(_00702_),
    .A1(_01474_),
    .S(_00532_),
    .X(_01475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12579_ (.A0(_01475_),
    .A1(_01473_),
    .S(_00537_),
    .X(\design_top.DATAO[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12580_ (.A0(_00693_),
    .A1(_01477_),
    .S(_00532_),
    .X(_01478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12581_ (.A0(_01478_),
    .A1(_01476_),
    .S(_00537_),
    .X(\design_top.DATAO[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12582_ (.A0(_00685_),
    .A1(_01480_),
    .S(_00532_),
    .X(_01481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12583_ (.A0(_01481_),
    .A1(_01479_),
    .S(_00537_),
    .X(\design_top.DATAO[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12584_ (.A0(_00676_),
    .A1(_01483_),
    .S(_00532_),
    .X(_01484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12585_ (.A0(_01484_),
    .A1(_01482_),
    .S(_00537_),
    .X(\design_top.DATAO[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12586_ (.A0(_00668_),
    .A1(_01486_),
    .S(_00532_),
    .X(_01487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12587_ (.A0(_01487_),
    .A1(_01485_),
    .S(_00537_),
    .X(\design_top.DATAO[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12588_ (.A0(_00659_),
    .A1(_01489_),
    .S(_00532_),
    .X(_01490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12589_ (.A0(_01490_),
    .A1(_01488_),
    .S(_00537_),
    .X(\design_top.DATAO[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12590_ (.A0(_00651_),
    .A1(_01492_),
    .S(_00532_),
    .X(_01493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12591_ (.A0(_01493_),
    .A1(_01491_),
    .S(_00537_),
    .X(\design_top.DATAO[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12592_ (.A0(_00642_),
    .A1(_01495_),
    .S(_00532_),
    .X(_01496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12593_ (.A0(_01496_),
    .A1(_01494_),
    .S(_00537_),
    .X(\design_top.DATAO[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12594_ (.A0(_00634_),
    .A1(_01498_),
    .S(_00532_),
    .X(_01499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12595_ (.A0(_01499_),
    .A1(_01497_),
    .S(_00537_),
    .X(\design_top.DATAO[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12596_ (.A0(_00625_),
    .A1(_01501_),
    .S(_00532_),
    .X(_01502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12597_ (.A0(_01502_),
    .A1(_01500_),
    .S(_00537_),
    .X(\design_top.DATAO[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12598_ (.A0(_00617_),
    .A1(_01504_),
    .S(_00532_),
    .X(_01505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12599_ (.A0(_01505_),
    .A1(_01503_),
    .S(_00537_),
    .X(\design_top.DATAO[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12600_ (.A0(_00608_),
    .A1(_01507_),
    .S(_00532_),
    .X(_01508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12601_ (.A0(_01508_),
    .A1(_01506_),
    .S(_00537_),
    .X(\design_top.DATAO[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12602_ (.A0(_00599_),
    .A1(_01510_),
    .S(_00532_),
    .X(_01511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12603_ (.A0(_01511_),
    .A1(_01509_),
    .S(_00537_),
    .X(\design_top.DATAO[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12604_ (.A0(_00582_),
    .A1(_00577_),
    .S(_00532_),
    .X(_00583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12605_ (.A0(_00583_),
    .A1(_00571_),
    .S(_00537_),
    .X(\design_top.DATAO[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12606_ (.A0(\design_top.ROMFF[7] ),
    .A1(\design_top.ROMFF2[7] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12607_ (.A0(\design_top.ROMFF[8] ),
    .A1(\design_top.ROMFF2[8] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12608_ (.A0(\design_top.ROMFF[9] ),
    .A1(\design_top.ROMFF2[9] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12609_ (.A0(\design_top.ROMFF[10] ),
    .A1(\design_top.ROMFF2[10] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12610_ (.A0(\design_top.ROMFF[12] ),
    .A1(\design_top.ROMFF2[12] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12611_ (.A0(\design_top.ROMFF[13] ),
    .A1(\design_top.ROMFF2[13] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12612_ (.A0(\design_top.ROMFF[14] ),
    .A1(\design_top.ROMFF2[14] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12613_ (.A0(\design_top.ROMFF[15] ),
    .A1(\design_top.ROMFF2[15] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12614_ (.A0(\design_top.ROMFF[16] ),
    .A1(\design_top.ROMFF2[16] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12615_ (.A0(\design_top.ROMFF[17] ),
    .A1(\design_top.ROMFF2[17] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12616_ (.A0(\design_top.ROMFF[18] ),
    .A1(\design_top.ROMFF2[18] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12617_ (.A0(\design_top.ROMFF[20] ),
    .A1(\design_top.ROMFF2[20] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12618_ (.A0(\design_top.ROMFF[21] ),
    .A1(\design_top.ROMFF2[21] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12619_ (.A0(\design_top.ROMFF[22] ),
    .A1(\design_top.ROMFF2[22] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12620_ (.A0(\design_top.ROMFF[23] ),
    .A1(\design_top.ROMFF2[23] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12621_ (.A0(\design_top.ROMFF[30] ),
    .A1(\design_top.ROMFF2[30] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12622_ (.A0(\design_top.ROMFF[31] ),
    .A1(\design_top.ROMFF2[31] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12623_ (.A0(_00923_),
    .A1(_00924_),
    .S(\design_top.uart0.UART_XSTATE[2] ),
    .X(_00925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12624_ (.A0(_00922_),
    .A1(_00925_),
    .S(\design_top.uart0.UART_XSTATE[3] ),
    .X(io_out[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12625_ (.A0(_00926_),
    .A1(_02512_),
    .S(_00344_),
    .X(_02513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12626_ (.A0(_02510_),
    .A1(_01562_),
    .S(_00586_),
    .X(_02511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12627_ (.A0(_01652_),
    .A1(_00535_),
    .S(_00589_),
    .X(_02404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12628_ (.A0(_01584_),
    .A1(_00540_),
    .S(_00589_),
    .X(_02403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12629_ (.A0(_02395_),
    .A1(_00893_),
    .S(_00538_),
    .X(_02396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12630_ (.A0(_02396_),
    .A1(_00601_),
    .S(_00864_),
    .X(_02397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12631_ (.A0(_01421_),
    .A1(_01878_),
    .S(_00534_),
    .X(_02398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12632_ (.A0(_02399_),
    .A1(_00387_),
    .S(_01434_),
    .X(_02400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12633_ (.A0(_02400_),
    .A1(_02383_),
    .S(_00590_),
    .X(_02401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12634_ (.A0(_02401_),
    .A1(_00914_),
    .S(_01437_),
    .X(_02402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12635_ (.A0(_02064_),
    .A1(_00381_),
    .S(_00808_),
    .X(_02392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12636_ (.A0(_02391_),
    .A1(_02392_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12637_ (.A0(_00594_),
    .A1(_00603_),
    .S(_00840_),
    .X(_02386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12638_ (.A0(_02386_),
    .A1(_02346_),
    .S(_00833_),
    .X(_02387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12639_ (.A0(_02387_),
    .A1(_02306_),
    .S(_00825_),
    .X(_02388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12640_ (.A0(_02388_),
    .A1(_02225_),
    .S(_00816_),
    .X(_02389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12641_ (.A0(_02389_),
    .A1(_02060_),
    .S(_00808_),
    .X(_02390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12642_ (.A0(_02375_),
    .A1(_00892_),
    .S(_00538_),
    .X(_02376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12643_ (.A0(_02376_),
    .A1(_00610_),
    .S(_00864_),
    .X(_02377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12644_ (.A0(_01421_),
    .A1(_01832_),
    .S(_00534_),
    .X(_02378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12645_ (.A0(_02379_),
    .A1(_00393_),
    .S(_01434_),
    .X(_02380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12646_ (.A0(_02380_),
    .A1(_02364_),
    .S(_00590_),
    .X(_02381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12647_ (.A0(_02381_),
    .A1(_00909_),
    .S(_01437_),
    .X(_02382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12648_ (.A0(_02037_),
    .A1(_00381_),
    .S(_00808_),
    .X(_02372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12649_ (.A0(_02371_),
    .A1(_02372_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12650_ (.A0(_01366_),
    .A1(_01368_),
    .S(_00833_),
    .X(_02367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12651_ (.A0(_02367_),
    .A1(_02284_),
    .S(_00825_),
    .X(_02368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12652_ (.A0(_02368_),
    .A1(_02203_),
    .S(_00816_),
    .X(_02369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12653_ (.A0(_02369_),
    .A1(_02033_),
    .S(_00808_),
    .X(_02370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12654_ (.A0(_02355_),
    .A1(_00891_),
    .S(_00538_),
    .X(_02356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12655_ (.A0(_02356_),
    .A1(_00619_),
    .S(_00864_),
    .X(_02357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12656_ (.A0(_01421_),
    .A1(_01789_),
    .S(_00534_),
    .X(_02358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12657_ (.A0(_02359_),
    .A1(_00399_),
    .S(_01434_),
    .X(_02360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12658_ (.A0(_02360_),
    .A1(_02342_),
    .S(_00590_),
    .X(_02361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12659_ (.A0(_02361_),
    .A1(_02362_),
    .S(_01437_),
    .X(_02363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12660_ (.A0(_02015_),
    .A1(_00381_),
    .S(_00808_),
    .X(_02352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12661_ (.A0(_02351_),
    .A1(_02352_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12662_ (.A0(_02346_),
    .A1(_02305_),
    .S(_00833_),
    .X(_02347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12663_ (.A0(_02347_),
    .A1(_02264_),
    .S(_00825_),
    .X(_02348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12664_ (.A0(_02348_),
    .A1(_02183_),
    .S(_00816_),
    .X(_02349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12665_ (.A0(_02349_),
    .A1(_02011_),
    .S(_00808_),
    .X(_02350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12666_ (.A0(_00612_),
    .A1(_00620_),
    .S(_00840_),
    .X(_02346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12667_ (.A0(_02333_),
    .A1(_00890_),
    .S(_00538_),
    .X(_02334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12668_ (.A0(_02334_),
    .A1(_00627_),
    .S(_00864_),
    .X(_02335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12669_ (.A0(_01421_),
    .A1(_01745_),
    .S(_00534_),
    .X(_02336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12670_ (.A0(_02337_),
    .A1(_00405_),
    .S(_01434_),
    .X(_02338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12671_ (.A0(_02338_),
    .A1(_02323_),
    .S(_00590_),
    .X(_02339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12672_ (.A0(_02339_),
    .A1(_02340_),
    .S(_01437_),
    .X(_02341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12673_ (.A0(_01991_),
    .A1(_00381_),
    .S(_00808_),
    .X(_02330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12674_ (.A0(_02329_),
    .A1(_02330_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12675_ (.A0(_01370_),
    .A1(_01374_),
    .S(_00825_),
    .X(_02326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12676_ (.A0(_02326_),
    .A1(_02161_),
    .S(_00816_),
    .X(_02327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12677_ (.A0(_02327_),
    .A1(_01987_),
    .S(_00808_),
    .X(_02328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12678_ (.A0(_02314_),
    .A1(_00889_),
    .S(_00538_),
    .X(_02315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12679_ (.A0(_02315_),
    .A1(_00636_),
    .S(_00864_),
    .X(_02316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12680_ (.A0(_01421_),
    .A1(_01697_),
    .S(_00534_),
    .X(_02317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12681_ (.A0(_02318_),
    .A1(_00411_),
    .S(_01434_),
    .X(_02319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12682_ (.A0(_02319_),
    .A1(_02301_),
    .S(_00590_),
    .X(_02320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12683_ (.A0(_02320_),
    .A1(_02321_),
    .S(_01437_),
    .X(_02322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12684_ (.A0(_01970_),
    .A1(_00381_),
    .S(_00808_),
    .X(_02311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12685_ (.A0(_02310_),
    .A1(_02311_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12686_ (.A0(_02306_),
    .A1(_02224_),
    .S(_00825_),
    .X(_02307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12687_ (.A0(_02307_),
    .A1(_02142_),
    .S(_00816_),
    .X(_02308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12688_ (.A0(_02308_),
    .A1(_01966_),
    .S(_00808_),
    .X(_02309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12689_ (.A0(_02305_),
    .A1(_02263_),
    .S(_00833_),
    .X(_02306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12690_ (.A0(_00629_),
    .A1(_00637_),
    .S(_00840_),
    .X(_02305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12691_ (.A0(_02292_),
    .A1(_00888_),
    .S(_00538_),
    .X(_02293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12692_ (.A0(_02293_),
    .A1(_00644_),
    .S(_00864_),
    .X(_02294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12693_ (.A0(_01421_),
    .A1(_01642_),
    .S(_00534_),
    .X(_02295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12694_ (.A0(_02296_),
    .A1(_00417_),
    .S(_01434_),
    .X(_02297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12695_ (.A0(_02297_),
    .A1(_02281_),
    .S(_00590_),
    .X(_02298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12696_ (.A0(_02298_),
    .A1(_02299_),
    .S(_01437_),
    .X(_02300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12697_ (.A0(_01946_),
    .A1(_00381_),
    .S(_00808_),
    .X(_02289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12698_ (.A0(_02288_),
    .A1(_02289_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12699_ (.A0(_02284_),
    .A1(_02202_),
    .S(_00825_),
    .X(_02285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12700_ (.A0(_02285_),
    .A1(_02119_),
    .S(_00816_),
    .X(_02286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12701_ (.A0(_02286_),
    .A1(_01942_),
    .S(_00808_),
    .X(_02287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12702_ (.A0(_01369_),
    .A1(_01372_),
    .S(_00833_),
    .X(_02284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12703_ (.A0(_02272_),
    .A1(_00887_),
    .S(_00538_),
    .X(_02273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12704_ (.A0(_02273_),
    .A1(_00653_),
    .S(_00864_),
    .X(_02274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12705_ (.A0(_01421_),
    .A1(_01574_),
    .S(_00534_),
    .X(_02275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12706_ (.A0(_02276_),
    .A1(_00423_),
    .S(_01434_),
    .X(_02277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12707_ (.A0(_02277_),
    .A1(_02259_),
    .S(_00590_),
    .X(_02278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12708_ (.A0(_02278_),
    .A1(_02279_),
    .S(_01437_),
    .X(_02280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12709_ (.A0(_01924_),
    .A1(_00381_),
    .S(_00808_),
    .X(_02269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12710_ (.A0(_02268_),
    .A1(_02269_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12711_ (.A0(_02264_),
    .A1(_02182_),
    .S(_00825_),
    .X(_02265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12712_ (.A0(_02265_),
    .A1(_02099_),
    .S(_00816_),
    .X(_02266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12713_ (.A0(_02266_),
    .A1(_01920_),
    .S(_00808_),
    .X(_02267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12714_ (.A0(_02263_),
    .A1(_02223_),
    .S(_00833_),
    .X(_02264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12715_ (.A0(_00646_),
    .A1(_00654_),
    .S(_00840_),
    .X(_02263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12716_ (.A0(_02250_),
    .A1(_00886_),
    .S(_00538_),
    .X(_02251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12717_ (.A0(_02251_),
    .A1(_00661_),
    .S(_00864_),
    .X(_02252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12718_ (.A0(_01421_),
    .A1(_01425_),
    .S(_00534_),
    .X(_02253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12719_ (.A0(_02254_),
    .A1(_00429_),
    .S(_01434_),
    .X(_02255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12720_ (.A0(_02255_),
    .A1(_02241_),
    .S(_00590_),
    .X(_02256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12721_ (.A0(_02256_),
    .A1(_02257_),
    .S(_01437_),
    .X(_02258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12722_ (.A0(_01900_),
    .A1(_00381_),
    .S(_00808_),
    .X(_02247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12723_ (.A0(_02246_),
    .A1(_02247_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12724_ (.A0(_01378_),
    .A1(_01388_),
    .S(_00816_),
    .X(_02244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12725_ (.A0(_02244_),
    .A1(_01893_),
    .S(_00808_),
    .X(_02245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12726_ (.A0(_02232_),
    .A1(_00885_),
    .S(_00538_),
    .X(_02233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12727_ (.A0(_02233_),
    .A1(_00670_),
    .S(_00864_),
    .X(_02234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12728_ (.A0(_01421_),
    .A1(_01873_),
    .S(_00534_),
    .X(_02235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12729_ (.A0(_02236_),
    .A1(_00435_),
    .S(_01434_),
    .X(_02237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12730_ (.A0(_02237_),
    .A1(_02219_),
    .S(_00590_),
    .X(_02238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12731_ (.A0(_02238_),
    .A1(_02239_),
    .S(_01437_),
    .X(_02240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12732_ (.A0(_01861_),
    .A1(_00381_),
    .S(_00808_),
    .X(_02229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12733_ (.A0(_02228_),
    .A1(_02229_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12734_ (.A0(_02225_),
    .A1(_02059_),
    .S(_00816_),
    .X(_02226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12735_ (.A0(_02226_),
    .A1(_01852_),
    .S(_00808_),
    .X(_02227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12736_ (.A0(_02224_),
    .A1(_02141_),
    .S(_00825_),
    .X(_02225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12737_ (.A0(_02223_),
    .A1(_02181_),
    .S(_00833_),
    .X(_02224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12738_ (.A0(_00663_),
    .A1(_00671_),
    .S(_00840_),
    .X(_02223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12739_ (.A0(_02210_),
    .A1(_00884_),
    .S(_00538_),
    .X(_02211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12740_ (.A0(_02211_),
    .A1(_00678_),
    .S(_00864_),
    .X(_02212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12741_ (.A0(_01421_),
    .A1(_01827_),
    .S(_00534_),
    .X(_02213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12742_ (.A0(_02214_),
    .A1(_00441_),
    .S(_01434_),
    .X(_02215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12743_ (.A0(_02215_),
    .A1(_02199_),
    .S(_00590_),
    .X(_02216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12744_ (.A0(_02216_),
    .A1(_02217_),
    .S(_01437_),
    .X(_02218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12745_ (.A0(_01815_),
    .A1(_00381_),
    .S(_00808_),
    .X(_02207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12746_ (.A0(_02206_),
    .A1(_02207_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12747_ (.A0(_02203_),
    .A1(_02032_),
    .S(_00816_),
    .X(_02204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12748_ (.A0(_02204_),
    .A1(_01806_),
    .S(_00808_),
    .X(_02205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12749_ (.A0(_02202_),
    .A1(_02118_),
    .S(_00825_),
    .X(_02203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12750_ (.A0(_01373_),
    .A1(_01375_),
    .S(_00833_),
    .X(_02202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12751_ (.A0(_02190_),
    .A1(_00883_),
    .S(_00538_),
    .X(_02191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12752_ (.A0(_02191_),
    .A1(_00687_),
    .S(_00864_),
    .X(_02192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12753_ (.A0(_01421_),
    .A1(_01784_),
    .S(_00534_),
    .X(_02193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12754_ (.A0(_02194_),
    .A1(_00447_),
    .S(_01434_),
    .X(_02195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12755_ (.A0(_02195_),
    .A1(_02177_),
    .S(_00590_),
    .X(_02196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12756_ (.A0(_02196_),
    .A1(_02197_),
    .S(_01437_),
    .X(_02198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12757_ (.A0(_01773_),
    .A1(_00381_),
    .S(_00808_),
    .X(_02187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12758_ (.A0(_02186_),
    .A1(_02187_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12759_ (.A0(_02183_),
    .A1(_02010_),
    .S(_00816_),
    .X(_02184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12760_ (.A0(_02184_),
    .A1(_01764_),
    .S(_00808_),
    .X(_02185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12761_ (.A0(_02182_),
    .A1(_02098_),
    .S(_00825_),
    .X(_02183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12762_ (.A0(_02181_),
    .A1(_02140_),
    .S(_00833_),
    .X(_02182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12763_ (.A0(_00680_),
    .A1(_00688_),
    .S(_00840_),
    .X(_02181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12764_ (.A0(_02168_),
    .A1(_00882_),
    .S(_00538_),
    .X(_02169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12765_ (.A0(_02169_),
    .A1(_00695_),
    .S(_00864_),
    .X(_02170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12766_ (.A0(_01421_),
    .A1(_01740_),
    .S(_00534_),
    .X(_02171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12767_ (.A0(_02172_),
    .A1(_00453_),
    .S(_01434_),
    .X(_02173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12768_ (.A0(_02173_),
    .A1(_02158_),
    .S(_00590_),
    .X(_02174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12769_ (.A0(_02174_),
    .A1(_02175_),
    .S(_01437_),
    .X(_02176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12770_ (.A0(_01729_),
    .A1(_00381_),
    .S(_00808_),
    .X(_02165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12771_ (.A0(_02164_),
    .A1(_02165_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12772_ (.A0(_02161_),
    .A1(_01986_),
    .S(_00816_),
    .X(_02162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12773_ (.A0(_02162_),
    .A1(_01713_),
    .S(_00808_),
    .X(_02163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12774_ (.A0(_01377_),
    .A1(_01382_),
    .S(_00825_),
    .X(_02161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12775_ (.A0(_02149_),
    .A1(_02137_),
    .S(_00538_),
    .X(_02150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12776_ (.A0(_02150_),
    .A1(_00704_),
    .S(_00864_),
    .X(_02151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12777_ (.A0(_01421_),
    .A1(_01692_),
    .S(_00534_),
    .X(_02152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12778_ (.A0(_02153_),
    .A1(_00459_),
    .S(_01434_),
    .X(_02154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12779_ (.A0(_02154_),
    .A1(_02135_),
    .S(_00590_),
    .X(_02155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12780_ (.A0(_02155_),
    .A1(_02156_),
    .S(_01437_),
    .X(_02157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12781_ (.A0(_01680_),
    .A1(_00381_),
    .S(_00808_),
    .X(_02146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12782_ (.A0(_02145_),
    .A1(_02146_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12783_ (.A0(_02142_),
    .A1(_01965_),
    .S(_00816_),
    .X(_02143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12784_ (.A0(_02143_),
    .A1(_01662_),
    .S(_00808_),
    .X(_02144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12785_ (.A0(_02141_),
    .A1(_02058_),
    .S(_00825_),
    .X(_02142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12786_ (.A0(_02140_),
    .A1(_02097_),
    .S(_00833_),
    .X(_02141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12787_ (.A0(_00697_),
    .A1(_00705_),
    .S(_00840_),
    .X(_02140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12788_ (.A0(_02126_),
    .A1(_00881_),
    .S(_00538_),
    .X(_02127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12789_ (.A0(_02127_),
    .A1(_00712_),
    .S(_00864_),
    .X(_02128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12790_ (.A0(_01421_),
    .A1(_01636_),
    .S(_00534_),
    .X(_02129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12791_ (.A0(_02130_),
    .A1(_00465_),
    .S(_01434_),
    .X(_02131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12792_ (.A0(_02131_),
    .A1(_02115_),
    .S(_00590_),
    .X(_02132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12793_ (.A0(_02132_),
    .A1(_02133_),
    .S(_01437_),
    .X(_02134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12794_ (.A0(_01625_),
    .A1(_00381_),
    .S(_00808_),
    .X(_02123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12795_ (.A0(_02122_),
    .A1(_02123_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12796_ (.A0(_02119_),
    .A1(_01941_),
    .S(_00816_),
    .X(_02120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12797_ (.A0(_02120_),
    .A1(_01592_),
    .S(_00808_),
    .X(_02121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12798_ (.A0(_02118_),
    .A1(_02031_),
    .S(_00825_),
    .X(_02119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12799_ (.A0(_01376_),
    .A1(_01380_),
    .S(_00833_),
    .X(_02118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12800_ (.A0(_02106_),
    .A1(_00880_),
    .S(_00538_),
    .X(_02107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12801_ (.A0(_02107_),
    .A1(_00721_),
    .S(_00864_),
    .X(_02108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12802_ (.A0(_01421_),
    .A1(_01567_),
    .S(_00534_),
    .X(_02109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12803_ (.A0(_02110_),
    .A1(_00471_),
    .S(_01434_),
    .X(_02111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12804_ (.A0(_02111_),
    .A1(_02093_),
    .S(_00590_),
    .X(_02112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12805_ (.A0(_02112_),
    .A1(_02113_),
    .S(_01437_),
    .X(_02114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12806_ (.A0(_01552_),
    .A1(_00381_),
    .S(_00808_),
    .X(_02103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12807_ (.A0(_02102_),
    .A1(_02103_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12808_ (.A0(_02099_),
    .A1(_01919_),
    .S(_00816_),
    .X(_02100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12809_ (.A0(_02100_),
    .A1(_01521_),
    .S(_00808_),
    .X(_02101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12810_ (.A0(_02098_),
    .A1(_02009_),
    .S(_00825_),
    .X(_02099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12811_ (.A0(_02097_),
    .A1(_02057_),
    .S(_00833_),
    .X(_02098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12812_ (.A0(_00714_),
    .A1(_00722_),
    .S(_00840_),
    .X(_02097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12813_ (.A0(_02084_),
    .A1(_00879_),
    .S(_00538_),
    .X(_02085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12814_ (.A0(_02085_),
    .A1(_00724_),
    .S(_00864_),
    .X(_02086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12815_ (.A0(_01420_),
    .A1(_01419_),
    .S(_00534_),
    .X(_02087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12816_ (.A0(_02088_),
    .A1(_00477_),
    .S(_01434_),
    .X(_02089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12817_ (.A0(_02089_),
    .A1(_02077_),
    .S(_00590_),
    .X(_02090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12818_ (.A0(_02090_),
    .A1(_02091_),
    .S(_01437_),
    .X(_02092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12819_ (.A0(_01896_),
    .A1(_01898_),
    .S(_00816_),
    .X(_02081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12820_ (.A0(_02067_),
    .A1(_02054_),
    .S(_00538_),
    .X(_02068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12821_ (.A0(_02068_),
    .A1(_00733_),
    .S(_00864_),
    .X(_02069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12822_ (.A0(_01878_),
    .A1(_01881_),
    .S(_00535_),
    .X(_02070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12823_ (.A0(_02070_),
    .A1(_01881_),
    .S(_00534_),
    .X(_02071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12824_ (.A0(_02072_),
    .A1(_00483_),
    .S(_01434_),
    .X(_02073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12825_ (.A0(_02073_),
    .A1(_02052_),
    .S(_00590_),
    .X(_02074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12826_ (.A0(_02074_),
    .A1(_02075_),
    .S(_01437_),
    .X(_02076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12827_ (.A0(_01860_),
    .A1(_00381_),
    .S(_00816_),
    .X(_02064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12828_ (.A0(_01855_),
    .A1(_01857_),
    .S(_00816_),
    .X(_02062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12829_ (.A0(_02059_),
    .A1(_01851_),
    .S(_00816_),
    .X(_02060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12830_ (.A0(_02058_),
    .A1(_01964_),
    .S(_00825_),
    .X(_02059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12831_ (.A0(_02057_),
    .A1(_02008_),
    .S(_00833_),
    .X(_02058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12832_ (.A0(_00726_),
    .A1(_00734_),
    .S(_00840_),
    .X(_02057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12833_ (.A0(_02040_),
    .A1(_00878_),
    .S(_00538_),
    .X(_02041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12834_ (.A0(_02041_),
    .A1(_00741_),
    .S(_00864_),
    .X(_02042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12835_ (.A0(_01832_),
    .A1(_01835_),
    .S(_00535_),
    .X(_02043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12836_ (.A0(_02043_),
    .A1(_01835_),
    .S(_00534_),
    .X(_02044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12837_ (.A0(_02045_),
    .A1(_00489_),
    .S(_01434_),
    .X(_02046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12838_ (.A0(_02046_),
    .A1(_02028_),
    .S(_00590_),
    .X(_02047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12839_ (.A0(_02047_),
    .A1(_02048_),
    .S(_01437_),
    .X(_02049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12840_ (.A0(_01814_),
    .A1(_00381_),
    .S(_00816_),
    .X(_02037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12841_ (.A0(_01809_),
    .A1(_01811_),
    .S(_00816_),
    .X(_02035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12842_ (.A0(_02032_),
    .A1(_01805_),
    .S(_00816_),
    .X(_02033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12843_ (.A0(_02031_),
    .A1(_01940_),
    .S(_00825_),
    .X(_02032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12844_ (.A0(_01381_),
    .A1(_01384_),
    .S(_00833_),
    .X(_02031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12845_ (.A0(_02018_),
    .A1(_00877_),
    .S(_00538_),
    .X(_02019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12846_ (.A0(_02019_),
    .A1(_00750_),
    .S(_00864_),
    .X(_02020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12847_ (.A0(_01789_),
    .A1(_01792_),
    .S(_00535_),
    .X(_02021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12848_ (.A0(_02021_),
    .A1(_01792_),
    .S(_00534_),
    .X(_02022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12849_ (.A0(_02023_),
    .A1(_00495_),
    .S(_01434_),
    .X(_02024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12850_ (.A0(_02024_),
    .A1(_02004_),
    .S(_00590_),
    .X(_02025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12851_ (.A0(_02025_),
    .A1(_02026_),
    .S(_01437_),
    .X(_02027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12852_ (.A0(_01772_),
    .A1(_00381_),
    .S(_00816_),
    .X(_02015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12853_ (.A0(_01767_),
    .A1(_01769_),
    .S(_00816_),
    .X(_02013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12854_ (.A0(_02010_),
    .A1(_01763_),
    .S(_00816_),
    .X(_02011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12855_ (.A0(_02009_),
    .A1(_01918_),
    .S(_00825_),
    .X(_02010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12856_ (.A0(_02008_),
    .A1(_01963_),
    .S(_00833_),
    .X(_02009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12857_ (.A0(_00743_),
    .A1(_01383_),
    .S(_00840_),
    .X(_02008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12858_ (.A0(_01994_),
    .A1(_00876_),
    .S(_00538_),
    .X(_01995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12859_ (.A0(_01995_),
    .A1(_00757_),
    .S(_00864_),
    .X(_01996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12860_ (.A0(_01745_),
    .A1(_01748_),
    .S(_00535_),
    .X(_01997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12861_ (.A0(_01997_),
    .A1(_01748_),
    .S(_00534_),
    .X(_01998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12862_ (.A0(_01999_),
    .A1(_00501_),
    .S(_01434_),
    .X(_02000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12863_ (.A0(_02000_),
    .A1(_01983_),
    .S(_00590_),
    .X(_02001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12864_ (.A0(_02001_),
    .A1(_02002_),
    .S(_01437_),
    .X(_02003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12865_ (.A0(_01728_),
    .A1(_00381_),
    .S(_00816_),
    .X(_01991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12866_ (.A0(_01720_),
    .A1(_01724_),
    .S(_00816_),
    .X(_01989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12867_ (.A0(_01986_),
    .A1(_01712_),
    .S(_00816_),
    .X(_01987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12868_ (.A0(_01387_),
    .A1(_01393_),
    .S(_00825_),
    .X(_01986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12869_ (.A0(_01973_),
    .A1(_00875_),
    .S(_00538_),
    .X(_01974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12870_ (.A0(_01974_),
    .A1(_00766_),
    .S(_00864_),
    .X(_01975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12871_ (.A0(_01697_),
    .A1(_01700_),
    .S(_00535_),
    .X(_01976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12872_ (.A0(_01976_),
    .A1(_01700_),
    .S(_00534_),
    .X(_01977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12873_ (.A0(_01978_),
    .A1(_00507_),
    .S(_01434_),
    .X(_01979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12874_ (.A0(_01979_),
    .A1(_01959_),
    .S(_00590_),
    .X(_01980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12875_ (.A0(_01980_),
    .A1(_01981_),
    .S(_01437_),
    .X(_01982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12876_ (.A0(_01679_),
    .A1(_00381_),
    .S(_00816_),
    .X(_01970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12877_ (.A0(_01669_),
    .A1(_01673_),
    .S(_00816_),
    .X(_01968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12878_ (.A0(_01965_),
    .A1(_01661_),
    .S(_00816_),
    .X(_01966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12879_ (.A0(_01964_),
    .A1(_01850_),
    .S(_00825_),
    .X(_01965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12880_ (.A0(_01963_),
    .A1(_01917_),
    .S(_00833_),
    .X(_01964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12881_ (.A0(_00759_),
    .A1(_01385_),
    .S(_00840_),
    .X(_01963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12882_ (.A0(_01949_),
    .A1(_00874_),
    .S(_00538_),
    .X(_01950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12883_ (.A0(_01950_),
    .A1(_00773_),
    .S(_00864_),
    .X(_01951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12884_ (.A0(_01642_),
    .A1(_01645_),
    .S(_00535_),
    .X(_01952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12885_ (.A0(_01952_),
    .A1(_01645_),
    .S(_00534_),
    .X(_01953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12886_ (.A0(_01954_),
    .A1(_00513_),
    .S(_01434_),
    .X(_01955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12887_ (.A0(_01955_),
    .A1(_01937_),
    .S(_00590_),
    .X(_01956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12888_ (.A0(_01956_),
    .A1(_01957_),
    .S(_01437_),
    .X(_01958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12889_ (.A0(_01624_),
    .A1(_00381_),
    .S(_00816_),
    .X(_01946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12890_ (.A0(_01607_),
    .A1(_01615_),
    .S(_00816_),
    .X(_01944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12891_ (.A0(_01941_),
    .A1(_01591_),
    .S(_00816_),
    .X(_01942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12892_ (.A0(_01940_),
    .A1(_01804_),
    .S(_00825_),
    .X(_01941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12893_ (.A0(_01386_),
    .A1(_01390_),
    .S(_00833_),
    .X(_01940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12894_ (.A0(_01927_),
    .A1(_00873_),
    .S(_00538_),
    .X(_01928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12895_ (.A0(_01928_),
    .A1(_00782_),
    .S(_00864_),
    .X(_01929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12896_ (.A0(_01574_),
    .A1(_01577_),
    .S(_00535_),
    .X(_01930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12897_ (.A0(_01930_),
    .A1(_01577_),
    .S(_00534_),
    .X(_01931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12898_ (.A0(_01932_),
    .A1(_00519_),
    .S(_01434_),
    .X(_01933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12899_ (.A0(_01933_),
    .A1(_01913_),
    .S(_00590_),
    .X(_01934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12900_ (.A0(_01934_),
    .A1(_01935_),
    .S(_01437_),
    .X(_01936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12901_ (.A0(_01551_),
    .A1(_00381_),
    .S(_00816_),
    .X(_01924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12902_ (.A0(_01536_),
    .A1(_01544_),
    .S(_00816_),
    .X(_01922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12903_ (.A0(_01919_),
    .A1(_01520_),
    .S(_00816_),
    .X(_01920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12904_ (.A0(_01918_),
    .A1(_01762_),
    .S(_00825_),
    .X(_01919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12905_ (.A0(_01917_),
    .A1(_01849_),
    .S(_00833_),
    .X(_01918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12906_ (.A0(_00775_),
    .A1(_01389_),
    .S(_00840_),
    .X(_01917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12907_ (.A0(_01903_),
    .A1(_00872_),
    .S(_00538_),
    .X(_01904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12908_ (.A0(_01904_),
    .A1(_00784_),
    .S(_00864_),
    .X(_01905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12909_ (.A0(_01425_),
    .A1(_01428_),
    .S(_00535_),
    .X(_01906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12910_ (.A0(_01906_),
    .A1(_01428_),
    .S(_00534_),
    .X(_01907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12911_ (.A0(_01908_),
    .A1(_00525_),
    .S(_01434_),
    .X(_01909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12912_ (.A0(_01909_),
    .A1(_01890_),
    .S(_00590_),
    .X(_01910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12913_ (.A0(_01910_),
    .A1(_01911_),
    .S(_01437_),
    .X(_01912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12914_ (.A0(_01898_),
    .A1(_00381_),
    .S(_00816_),
    .X(_01900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12915_ (.A0(_01898_),
    .A1(_01402_),
    .S(_00816_),
    .X(_01899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12916_ (.A0(_01723_),
    .A1(_01725_),
    .S(_00825_),
    .X(_01898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12917_ (.A0(_01716_),
    .A1(_01718_),
    .S(_00825_),
    .X(_01895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12918_ (.A0(_01895_),
    .A1(_01896_),
    .S(_00816_),
    .X(_01897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12919_ (.A0(_01719_),
    .A1(_01722_),
    .S(_00825_),
    .X(_01896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12920_ (.A0(_01864_),
    .A1(_01846_),
    .S(_00538_),
    .X(_01865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12921_ (.A0(_01865_),
    .A1(_00793_),
    .S(_00864_),
    .X(_01866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12922_ (.A0(_01869_),
    .A1(_01881_),
    .S(_00545_),
    .X(_01882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12923_ (.A0(_01882_),
    .A1(_01873_),
    .S(_00907_),
    .X(_01883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12924_ (.A0(_01883_),
    .A1(_01878_),
    .S(_00551_),
    .X(_01884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12925_ (.A0(_01873_),
    .A1(_01869_),
    .S(_00535_),
    .X(_01874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12926_ (.A0(_01874_),
    .A1(_01869_),
    .S(_00534_),
    .X(_01875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12927_ (.A0(_01885_),
    .A1(_00531_),
    .S(_01434_),
    .X(_01886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12928_ (.A0(_01886_),
    .A1(_01844_),
    .S(_00590_),
    .X(_01887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12929_ (.A0(_01887_),
    .A1(_01888_),
    .S(_01437_),
    .X(_01889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12930_ (.A0(_01879_),
    .A1(_01880_),
    .S(\design_top.XADDR[31] ),
    .X(_01881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12931_ (.A0(_01876_),
    .A1(_01877_),
    .S(\design_top.XADDR[31] ),
    .X(_01878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12932_ (.A0(_01571_),
    .A1(_01871_),
    .S(\design_top.XADDR[3] ),
    .X(_01872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12933_ (.A0(_01870_),
    .A1(_01872_),
    .S(\design_top.XADDR[31] ),
    .X(_01873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12934_ (.A0(_01867_),
    .A1(_01868_),
    .S(\design_top.XADDR[31] ),
    .X(_01869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12935_ (.A0(_01857_),
    .A1(_01860_),
    .S(_00816_),
    .X(_01861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12936_ (.A0(_01678_),
    .A1(_00381_),
    .S(_00825_),
    .X(_01860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12937_ (.A0(_01857_),
    .A1(_01858_),
    .S(_00816_),
    .X(_01859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12938_ (.A0(_01672_),
    .A1(_01674_),
    .S(_00825_),
    .X(_01857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12939_ (.A0(_01665_),
    .A1(_01667_),
    .S(_00825_),
    .X(_01854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12940_ (.A0(_01854_),
    .A1(_01855_),
    .S(_00816_),
    .X(_01856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12941_ (.A0(_01668_),
    .A1(_01671_),
    .S(_00825_),
    .X(_01855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12942_ (.A0(_01850_),
    .A1(_01660_),
    .S(_00825_),
    .X(_01851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12943_ (.A0(_01849_),
    .A1(_01761_),
    .S(_00833_),
    .X(_01850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12944_ (.A0(_00786_),
    .A1(_01391_),
    .S(_00840_),
    .X(_01849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12945_ (.A0(_01818_),
    .A1(_00871_),
    .S(_00538_),
    .X(_01819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12946_ (.A0(_01819_),
    .A1(_00800_),
    .S(_00864_),
    .X(_01820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12947_ (.A0(_01823_),
    .A1(_01835_),
    .S(_00545_),
    .X(_01836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12948_ (.A0(_01836_),
    .A1(_01827_),
    .S(_00907_),
    .X(_01837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12949_ (.A0(_01837_),
    .A1(_01832_),
    .S(_00551_),
    .X(_01838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12950_ (.A0(_01827_),
    .A1(_01823_),
    .S(_00535_),
    .X(_01828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12951_ (.A0(_01828_),
    .A1(_01823_),
    .S(_00534_),
    .X(_01829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12952_ (.A0(_01839_),
    .A1(_00354_),
    .S(_01434_),
    .X(_01840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12953_ (.A0(_01840_),
    .A1(_01801_),
    .S(_00590_),
    .X(_01841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12954_ (.A0(_01841_),
    .A1(_01842_),
    .S(_01437_),
    .X(_01843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12955_ (.A0(_01833_),
    .A1(_01834_),
    .S(\design_top.XADDR[31] ),
    .X(_01835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12956_ (.A0(_01830_),
    .A1(_01831_),
    .S(\design_top.XADDR[31] ),
    .X(_01832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12957_ (.A0(_01571_),
    .A1(_01825_),
    .S(\design_top.XADDR[3] ),
    .X(_01826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12958_ (.A0(_01824_),
    .A1(_01826_),
    .S(\design_top.XADDR[31] ),
    .X(_01827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12959_ (.A0(_01821_),
    .A1(_01822_),
    .S(\design_top.XADDR[31] ),
    .X(_01823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12960_ (.A0(_01811_),
    .A1(_01814_),
    .S(_00816_),
    .X(_01815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12961_ (.A0(_01623_),
    .A1(_00381_),
    .S(_00825_),
    .X(_01814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12962_ (.A0(_01811_),
    .A1(_01812_),
    .S(_00816_),
    .X(_01813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12963_ (.A0(_01614_),
    .A1(_01618_),
    .S(_00825_),
    .X(_01811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12964_ (.A0(_01599_),
    .A1(_01603_),
    .S(_00825_),
    .X(_01808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12965_ (.A0(_01808_),
    .A1(_01809_),
    .S(_00816_),
    .X(_01810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12966_ (.A0(_01606_),
    .A1(_01611_),
    .S(_00825_),
    .X(_01809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12967_ (.A0(_01804_),
    .A1(_01590_),
    .S(_00825_),
    .X(_01805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12968_ (.A0(_01392_),
    .A1(_01394_),
    .S(_00833_),
    .X(_01804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12969_ (.A0(_01776_),
    .A1(_00870_),
    .S(_00538_),
    .X(_01777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12970_ (.A0(_01777_),
    .A1(_00809_),
    .S(_00864_),
    .X(_01778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12971_ (.A0(_01781_),
    .A1(_01792_),
    .S(_00545_),
    .X(_01793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12972_ (.A0(_01793_),
    .A1(_01784_),
    .S(_00907_),
    .X(_01794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12973_ (.A0(_01794_),
    .A1(_01789_),
    .S(_00551_),
    .X(_01795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12974_ (.A0(_01784_),
    .A1(_01781_),
    .S(_00535_),
    .X(_01785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12975_ (.A0(_01785_),
    .A1(_01781_),
    .S(_00534_),
    .X(_01786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12976_ (.A0(_01796_),
    .A1(_00347_),
    .S(_01434_),
    .X(_01797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12977_ (.A0(_01797_),
    .A1(_01757_),
    .S(_00590_),
    .X(_01798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12978_ (.A0(_01798_),
    .A1(_01799_),
    .S(_01437_),
    .X(_01800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12979_ (.A0(_01790_),
    .A1(_01791_),
    .S(\design_top.XADDR[31] ),
    .X(_01792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12980_ (.A0(_01787_),
    .A1(_01788_),
    .S(\design_top.XADDR[31] ),
    .X(_01789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12981_ (.A0(_01782_),
    .A1(_01783_),
    .S(\design_top.XADDR[31] ),
    .X(_01784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12982_ (.A0(_01779_),
    .A1(_01780_),
    .S(\design_top.XADDR[31] ),
    .X(_01781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12983_ (.A0(_01769_),
    .A1(_01772_),
    .S(_00816_),
    .X(_01773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12984_ (.A0(_01550_),
    .A1(_00381_),
    .S(_00825_),
    .X(_01772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12985_ (.A0(_01769_),
    .A1(_01770_),
    .S(_00816_),
    .X(_01771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12986_ (.A0(_01543_),
    .A1(_01547_),
    .S(_00825_),
    .X(_01769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12987_ (.A0(_01528_),
    .A1(_01532_),
    .S(_00825_),
    .X(_01766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12988_ (.A0(_01766_),
    .A1(_01767_),
    .S(_00816_),
    .X(_01768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12989_ (.A0(_01535_),
    .A1(_01540_),
    .S(_00825_),
    .X(_01767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12990_ (.A0(_01762_),
    .A1(_01519_),
    .S(_00825_),
    .X(_01763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12991_ (.A0(_01761_),
    .A1(_01659_),
    .S(_00833_),
    .X(_01762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12992_ (.A0(_00802_),
    .A1(_00810_),
    .S(_00840_),
    .X(_01761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12993_ (.A0(_01732_),
    .A1(_00869_),
    .S(_00538_),
    .X(_01733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12994_ (.A0(_01733_),
    .A1(_00817_),
    .S(_00864_),
    .X(_01734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12995_ (.A0(_01737_),
    .A1(_01748_),
    .S(_00545_),
    .X(_01749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12996_ (.A0(_01749_),
    .A1(_01740_),
    .S(_00907_),
    .X(_01750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12997_ (.A0(_01750_),
    .A1(_01745_),
    .S(_00551_),
    .X(_01751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12998_ (.A0(_01740_),
    .A1(_01737_),
    .S(_00535_),
    .X(_01741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _12999_ (.A0(_01741_),
    .A1(_01737_),
    .S(_00534_),
    .X(_01742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13000_ (.A0(_01752_),
    .A1(_00335_),
    .S(_01434_),
    .X(_01753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13001_ (.A0(_01753_),
    .A1(_01709_),
    .S(_00590_),
    .X(_01754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13002_ (.A0(_01754_),
    .A1(_01755_),
    .S(_01437_),
    .X(_01756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13003_ (.A0(_01746_),
    .A1(_01747_),
    .S(\design_top.XADDR[31] ),
    .X(_01748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13004_ (.A0(_01743_),
    .A1(_01744_),
    .S(\design_top.XADDR[31] ),
    .X(_01745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13005_ (.A0(_01738_),
    .A1(_01739_),
    .S(\design_top.XADDR[31] ),
    .X(_01740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13006_ (.A0(_01735_),
    .A1(_01736_),
    .S(\design_top.XADDR[31] ),
    .X(_01737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13007_ (.A0(_01724_),
    .A1(_01728_),
    .S(_00816_),
    .X(_01729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13008_ (.A0(_01725_),
    .A1(_00381_),
    .S(_00825_),
    .X(_01728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13009_ (.A0(_01724_),
    .A1(_01726_),
    .S(_00816_),
    .X(_01727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13010_ (.A0(_01725_),
    .A1(_01401_),
    .S(_00825_),
    .X(_01726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13011_ (.A0(_01617_),
    .A1(_01619_),
    .S(_00833_),
    .X(_01725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13012_ (.A0(_01722_),
    .A1(_01723_),
    .S(_00825_),
    .X(_01724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13013_ (.A0(_01613_),
    .A1(_01616_),
    .S(_00833_),
    .X(_01723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13014_ (.A0(_01610_),
    .A1(_01612_),
    .S(_00833_),
    .X(_01722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13015_ (.A0(_01595_),
    .A1(_01597_),
    .S(_00833_),
    .X(_01715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13016_ (.A0(_01715_),
    .A1(_01716_),
    .S(_00825_),
    .X(_01717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13017_ (.A0(_01717_),
    .A1(_01720_),
    .S(_00816_),
    .X(_01721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13018_ (.A0(_01718_),
    .A1(_01719_),
    .S(_00825_),
    .X(_01720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13019_ (.A0(_01605_),
    .A1(_01609_),
    .S(_00833_),
    .X(_01719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13020_ (.A0(_01602_),
    .A1(_01604_),
    .S(_00833_),
    .X(_01718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13021_ (.A0(_01598_),
    .A1(_01601_),
    .S(_00833_),
    .X(_01716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13022_ (.A0(_01683_),
    .A1(_01656_),
    .S(_00538_),
    .X(_01684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13023_ (.A0(_01684_),
    .A1(_00826_),
    .S(_00864_),
    .X(_01685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13024_ (.A0(_01688_),
    .A1(_01700_),
    .S(_00545_),
    .X(_01701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13025_ (.A0(_01701_),
    .A1(_01692_),
    .S(_00907_),
    .X(_01702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13026_ (.A0(_01702_),
    .A1(_01697_),
    .S(_00551_),
    .X(_01703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13027_ (.A0(_01692_),
    .A1(_01688_),
    .S(_00535_),
    .X(_01693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13028_ (.A0(_01693_),
    .A1(_01688_),
    .S(_00534_),
    .X(_01694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13029_ (.A0(_01704_),
    .A1(_00310_),
    .S(_01434_),
    .X(_01705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13030_ (.A0(_01705_),
    .A1(_01654_),
    .S(_00590_),
    .X(_01706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13031_ (.A0(_01706_),
    .A1(_01707_),
    .S(_01437_),
    .X(_01708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13032_ (.A0(_01698_),
    .A1(_01699_),
    .S(\design_top.XADDR[31] ),
    .X(_01700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13033_ (.A0(_01695_),
    .A1(_01696_),
    .S(\design_top.XADDR[31] ),
    .X(_01697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13034_ (.A0(_01571_),
    .A1(_01690_),
    .S(\design_top.XADDR[3] ),
    .X(_01691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13035_ (.A0(_01689_),
    .A1(_01691_),
    .S(\design_top.XADDR[31] ),
    .X(_01692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13036_ (.A0(_01686_),
    .A1(_01687_),
    .S(\design_top.XADDR[31] ),
    .X(_01688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13037_ (.A0(_01673_),
    .A1(_01679_),
    .S(_00816_),
    .X(_01680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13038_ (.A0(_01674_),
    .A1(_01678_),
    .S(_00825_),
    .X(_01679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13039_ (.A0(_01549_),
    .A1(_00381_),
    .S(_00833_),
    .X(_01678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13040_ (.A0(_01673_),
    .A1(_01676_),
    .S(_00816_),
    .X(_01677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13041_ (.A0(_01674_),
    .A1(_01675_),
    .S(_00825_),
    .X(_01676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13042_ (.A0(_01546_),
    .A1(_01548_),
    .S(_00833_),
    .X(_01674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13043_ (.A0(_01671_),
    .A1(_01672_),
    .S(_00825_),
    .X(_01673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13044_ (.A0(_01542_),
    .A1(_01545_),
    .S(_00833_),
    .X(_01672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13045_ (.A0(_01539_),
    .A1(_01541_),
    .S(_00833_),
    .X(_01671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13046_ (.A0(_01524_),
    .A1(_01526_),
    .S(_00833_),
    .X(_01664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13047_ (.A0(_01664_),
    .A1(_01665_),
    .S(_00825_),
    .X(_01666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13048_ (.A0(_01666_),
    .A1(_01669_),
    .S(_00816_),
    .X(_01670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13049_ (.A0(_01667_),
    .A1(_01668_),
    .S(_00825_),
    .X(_01669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13050_ (.A0(_01534_),
    .A1(_01538_),
    .S(_00833_),
    .X(_01668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13051_ (.A0(_01531_),
    .A1(_01533_),
    .S(_00833_),
    .X(_01667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13052_ (.A0(_01527_),
    .A1(_01530_),
    .S(_00833_),
    .X(_01665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13053_ (.A0(_01659_),
    .A1(_01518_),
    .S(_00833_),
    .X(_01660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13054_ (.A0(_00819_),
    .A1(_00827_),
    .S(_00840_),
    .X(_01659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13055_ (.A0(_01628_),
    .A1(_00834_),
    .S(_00538_),
    .X(_01629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13056_ (.A0(_01629_),
    .A1(_01587_),
    .S(_00864_),
    .X(_01630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13057_ (.A0(_01633_),
    .A1(_01645_),
    .S(_00545_),
    .X(_01646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13058_ (.A0(_01646_),
    .A1(_01636_),
    .S(_00907_),
    .X(_01647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13059_ (.A0(_01647_),
    .A1(_01642_),
    .S(_00551_),
    .X(_01648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13060_ (.A0(_01636_),
    .A1(_01633_),
    .S(_00535_),
    .X(_01637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13061_ (.A0(_01637_),
    .A1(_01633_),
    .S(_00534_),
    .X(_01638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13062_ (.A0(_01649_),
    .A1(_00325_),
    .S(_01434_),
    .X(_01650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13063_ (.A0(_01650_),
    .A1(_01586_),
    .S(_00590_),
    .X(_01651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13064_ (.A0(_01651_),
    .A1(_01652_),
    .S(_01437_),
    .X(_01653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13065_ (.A0(_01643_),
    .A1(_01644_),
    .S(\design_top.XADDR[31] ),
    .X(_01645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13066_ (.A0(_01571_),
    .A1(_01640_),
    .S(\design_top.XADDR[3] ),
    .X(_01641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13067_ (.A0(_01639_),
    .A1(_01641_),
    .S(\design_top.XADDR[31] ),
    .X(_01642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13068_ (.A0(_01634_),
    .A1(_01635_),
    .S(\design_top.XADDR[31] ),
    .X(_01636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13069_ (.A0(_01631_),
    .A1(_01632_),
    .S(\design_top.XADDR[31] ),
    .X(_01633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13070_ (.A0(_01615_),
    .A1(_01624_),
    .S(_00816_),
    .X(_01625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13071_ (.A0(_01618_),
    .A1(_01623_),
    .S(_00825_),
    .X(_01624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13072_ (.A0(_01619_),
    .A1(_00381_),
    .S(_00833_),
    .X(_01623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13073_ (.A0(_01615_),
    .A1(_01621_),
    .S(_00816_),
    .X(_01622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13074_ (.A0(_01618_),
    .A1(_01620_),
    .S(_00825_),
    .X(_01621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13075_ (.A0(_01619_),
    .A1(_01400_),
    .S(_00833_),
    .X(_01620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13076_ (.A0(_00603_),
    .A1(_00594_),
    .S(_00840_),
    .X(_01619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13077_ (.A0(_01616_),
    .A1(_01617_),
    .S(_00833_),
    .X(_01618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13078_ (.A0(_00620_),
    .A1(_00612_),
    .S(_00840_),
    .X(_01617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13079_ (.A0(_00637_),
    .A1(_00629_),
    .S(_00840_),
    .X(_01616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13080_ (.A0(_01611_),
    .A1(_01614_),
    .S(_00825_),
    .X(_01615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13081_ (.A0(_01612_),
    .A1(_01613_),
    .S(_00833_),
    .X(_01614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13082_ (.A0(_00654_),
    .A1(_00646_),
    .S(_00840_),
    .X(_01613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13083_ (.A0(_00671_),
    .A1(_00663_),
    .S(_00840_),
    .X(_01612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13084_ (.A0(_01609_),
    .A1(_01610_),
    .S(_00833_),
    .X(_01611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13085_ (.A0(_00688_),
    .A1(_00680_),
    .S(_00840_),
    .X(_01610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13086_ (.A0(_00705_),
    .A1(_00697_),
    .S(_00840_),
    .X(_01609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13087_ (.A0(_00827_),
    .A1(_00819_),
    .S(_00840_),
    .X(_01594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13088_ (.A0(_01594_),
    .A1(_01595_),
    .S(_00833_),
    .X(_01596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13089_ (.A0(_01596_),
    .A1(_01599_),
    .S(_00825_),
    .X(_01600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13090_ (.A0(_01600_),
    .A1(_01607_),
    .S(_00816_),
    .X(_01608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13091_ (.A0(_01603_),
    .A1(_01606_),
    .S(_00825_),
    .X(_01607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13092_ (.A0(_01604_),
    .A1(_01605_),
    .S(_00833_),
    .X(_01606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13093_ (.A0(_00722_),
    .A1(_00714_),
    .S(_00840_),
    .X(_01605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13094_ (.A0(_00734_),
    .A1(_00726_),
    .S(_00840_),
    .X(_01604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13095_ (.A0(_01601_),
    .A1(_01602_),
    .S(_00833_),
    .X(_01603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13096_ (.A0(_01383_),
    .A1(_00743_),
    .S(_00840_),
    .X(_01602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13097_ (.A0(_01385_),
    .A1(_00759_),
    .S(_00840_),
    .X(_01601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13098_ (.A0(_01597_),
    .A1(_01598_),
    .S(_00833_),
    .X(_01599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13099_ (.A0(_01389_),
    .A1(_00775_),
    .S(_00840_),
    .X(_01598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13100_ (.A0(_01391_),
    .A1(_00786_),
    .S(_00840_),
    .X(_01597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13101_ (.A0(_00810_),
    .A1(_00802_),
    .S(_00840_),
    .X(_01595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13102_ (.A0(_01554_),
    .A1(_01522_),
    .S(_00532_),
    .X(_01555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13103_ (.A0(_01555_),
    .A1(_00868_),
    .S(_00537_),
    .X(_01556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13104_ (.A0(_01556_),
    .A1(_00841_),
    .S(_01407_),
    .X(_01557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13105_ (.A0(_01557_),
    .A1(_00863_),
    .S(_01408_),
    .X(_01558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13106_ (.A0(_01558_),
    .A1(_00868_),
    .S(_00538_),
    .X(_01559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13107_ (.A0(_01559_),
    .A1(_01517_),
    .S(_00864_),
    .X(_01560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13108_ (.A0(_01564_),
    .A1(_01577_),
    .S(_00545_),
    .X(_01578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13109_ (.A0(_01578_),
    .A1(_01567_),
    .S(_00907_),
    .X(_01579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13110_ (.A0(_01579_),
    .A1(_01574_),
    .S(_00551_),
    .X(_01580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13111_ (.A0(_01567_),
    .A1(_01564_),
    .S(_00535_),
    .X(_01568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13112_ (.A0(_01568_),
    .A1(_01564_),
    .S(_00534_),
    .X(_01569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13113_ (.A0(_01581_),
    .A1(_00326_),
    .S(_01434_),
    .X(_01582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13114_ (.A0(_01582_),
    .A1(_01515_),
    .S(_00590_),
    .X(_01583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13115_ (.A0(_01583_),
    .A1(_01584_),
    .S(_01437_),
    .X(_01585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13116_ (.A0(_01575_),
    .A1(_01576_),
    .S(\design_top.XADDR[31] ),
    .X(_01577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13117_ (.A0(_01571_),
    .A1(_01572_),
    .S(\design_top.XADDR[3] ),
    .X(_01573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13118_ (.A0(_01570_),
    .A1(_01573_),
    .S(\design_top.XADDR[31] ),
    .X(_01574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13119_ (.A0(_01565_),
    .A1(_01566_),
    .S(\design_top.XADDR[31] ),
    .X(_01567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13120_ (.A0(_01561_),
    .A1(_01563_),
    .S(\design_top.XADDR[31] ),
    .X(_01564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13121_ (.A0(_00867_),
    .A1(_00827_),
    .S(_00840_),
    .X(_01523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13122_ (.A0(_01523_),
    .A1(_01524_),
    .S(_00833_),
    .X(_01525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13123_ (.A0(_01525_),
    .A1(_01528_),
    .S(_00825_),
    .X(_01529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13124_ (.A0(_01529_),
    .A1(_01536_),
    .S(_00816_),
    .X(_01537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13125_ (.A0(_01537_),
    .A1(_01552_),
    .S(_00808_),
    .X(_01553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13126_ (.A0(_01544_),
    .A1(_01551_),
    .S(_00816_),
    .X(_01552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13127_ (.A0(_01547_),
    .A1(_01550_),
    .S(_00825_),
    .X(_01551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13128_ (.A0(_01548_),
    .A1(_01549_),
    .S(_00833_),
    .X(_01550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13129_ (.A0(_00594_),
    .A1(_00381_),
    .S(_00840_),
    .X(_01549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13130_ (.A0(_00612_),
    .A1(_00603_),
    .S(_00840_),
    .X(_01548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13131_ (.A0(_01545_),
    .A1(_01546_),
    .S(_00833_),
    .X(_01547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13132_ (.A0(_00629_),
    .A1(_00620_),
    .S(_00840_),
    .X(_01546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13133_ (.A0(_00646_),
    .A1(_00637_),
    .S(_00840_),
    .X(_01545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13134_ (.A0(_01540_),
    .A1(_01543_),
    .S(_00825_),
    .X(_01544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13135_ (.A0(_01541_),
    .A1(_01542_),
    .S(_00833_),
    .X(_01543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13136_ (.A0(_00663_),
    .A1(_00654_),
    .S(_00840_),
    .X(_01542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13137_ (.A0(_00680_),
    .A1(_00671_),
    .S(_00840_),
    .X(_01541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13138_ (.A0(_01538_),
    .A1(_01539_),
    .S(_00833_),
    .X(_01540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13139_ (.A0(_00697_),
    .A1(_00688_),
    .S(_00840_),
    .X(_01539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13140_ (.A0(_00714_),
    .A1(_00705_),
    .S(_00840_),
    .X(_01538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13141_ (.A0(_01532_),
    .A1(_01535_),
    .S(_00825_),
    .X(_01536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13142_ (.A0(_01533_),
    .A1(_01534_),
    .S(_00833_),
    .X(_01535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13143_ (.A0(_00726_),
    .A1(_00722_),
    .S(_00840_),
    .X(_01534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13144_ (.A0(_00743_),
    .A1(_00734_),
    .S(_00840_),
    .X(_01533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13145_ (.A0(_01530_),
    .A1(_01531_),
    .S(_00833_),
    .X(_01532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13146_ (.A0(_00759_),
    .A1(_01383_),
    .S(_00840_),
    .X(_01531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13147_ (.A0(_00775_),
    .A1(_01385_),
    .S(_00840_),
    .X(_01530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13148_ (.A0(_01526_),
    .A1(_01527_),
    .S(_00833_),
    .X(_01528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13149_ (.A0(_00786_),
    .A1(_01389_),
    .S(_00840_),
    .X(_01527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13150_ (.A0(_00802_),
    .A1(_01391_),
    .S(_00840_),
    .X(_01526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13151_ (.A0(_00819_),
    .A1(_00810_),
    .S(_00840_),
    .X(_01524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13152_ (.A0(\design_top.core0.XIDATA[10] ),
    .A1(\design_top.core0.RESMODE[3] ),
    .S(\design_top.core0.XRES ),
    .X(_01442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13153_ (.A0(\design_top.core0.XIDATA[9] ),
    .A1(\design_top.core0.RESMODE[2] ),
    .S(\design_top.core0.XRES ),
    .X(_01441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13154_ (.A0(\design_top.core0.XIDATA[8] ),
    .A1(\design_top.core0.RESMODE[1] ),
    .S(\design_top.core0.XRES ),
    .X(_01440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13155_ (.A0(\design_top.core0.XIDATA[7] ),
    .A1(\design_top.core0.RESMODE[0] ),
    .S(\design_top.core0.XRES ),
    .X(_01439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13156_ (.A0(_01409_),
    .A1(_00894_),
    .S(_00538_),
    .X(_01410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13157_ (.A0(_01410_),
    .A1(_00592_),
    .S(_00864_),
    .X(_01411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13158_ (.A0(_01421_),
    .A1(_01416_),
    .S(_00534_),
    .X(_01422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13159_ (.A0(_01433_),
    .A1(_01360_),
    .S(_01434_),
    .X(_01435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13160_ (.A0(_01435_),
    .A1(_01359_),
    .S(_00590_),
    .X(_01436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13161_ (.A0(_01436_),
    .A1(_00919_),
    .S(_01437_),
    .X(_01438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13162_ (.A0(_01428_),
    .A1(_01419_),
    .S(_00545_),
    .X(_01429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13163_ (.A0(_01429_),
    .A1(_01425_),
    .S(_00907_),
    .X(_01430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13164_ (.A0(_01430_),
    .A1(_01416_),
    .S(_00551_),
    .X(_01431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13165_ (.A0(_01426_),
    .A1(_01427_),
    .S(\design_top.XADDR[31] ),
    .X(_01428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13166_ (.A0(_01423_),
    .A1(_01424_),
    .S(\design_top.XADDR[31] ),
    .X(_01425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13167_ (.A0(_01416_),
    .A1(_01419_),
    .S(_00535_),
    .X(_01420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13168_ (.A0(_01417_),
    .A1(_01418_),
    .S(\design_top.XADDR[31] ),
    .X(_01419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13169_ (.A0(_01414_),
    .A1(_00346_),
    .S(_01413_),
    .X(_01415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13170_ (.A0(_01412_),
    .A1(_01415_),
    .S(\design_top.XADDR[31] ),
    .X(_01416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13171_ (.A0(_01404_),
    .A1(_00381_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_01405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13172_ (.A0(_00381_),
    .A1(_00594_),
    .S(_00840_),
    .X(_01365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13173_ (.A0(_01365_),
    .A1(_01366_),
    .S(_00833_),
    .X(_01367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13174_ (.A0(_01367_),
    .A1(_01370_),
    .S(_00825_),
    .X(_01371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13175_ (.A0(_01371_),
    .A1(_01378_),
    .S(_00816_),
    .X(_01379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13176_ (.A0(_01379_),
    .A1(_01398_),
    .S(_00808_),
    .X(_01399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13177_ (.A0(_01388_),
    .A1(_01397_),
    .S(_00816_),
    .X(_01398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13178_ (.A0(_01393_),
    .A1(_01396_),
    .S(_00825_),
    .X(_01397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13179_ (.A0(_01394_),
    .A1(_01395_),
    .S(_00833_),
    .X(_01396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13180_ (.A0(_00827_),
    .A1(_00867_),
    .S(_00840_),
    .X(_01395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13181_ (.A0(_00810_),
    .A1(_00819_),
    .S(_00840_),
    .X(_01394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13182_ (.A0(_01390_),
    .A1(_01392_),
    .S(_00833_),
    .X(_01393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13183_ (.A0(_01391_),
    .A1(_00802_),
    .S(_00840_),
    .X(_01392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13184_ (.A0(_01389_),
    .A1(_00786_),
    .S(_00840_),
    .X(_01390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13185_ (.A0(_01382_),
    .A1(_01387_),
    .S(_00825_),
    .X(_01388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13186_ (.A0(_01384_),
    .A1(_01386_),
    .S(_00833_),
    .X(_01387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13187_ (.A0(_01385_),
    .A1(_00775_),
    .S(_00840_),
    .X(_01386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13188_ (.A0(_01383_),
    .A1(_00759_),
    .S(_00840_),
    .X(_01384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13189_ (.A0(_01380_),
    .A1(_01381_),
    .S(_00833_),
    .X(_01382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13190_ (.A0(_00734_),
    .A1(_00743_),
    .S(_00840_),
    .X(_01381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13191_ (.A0(_00722_),
    .A1(_00726_),
    .S(_00840_),
    .X(_01380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13192_ (.A0(_01374_),
    .A1(_01377_),
    .S(_00825_),
    .X(_01378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13193_ (.A0(_01375_),
    .A1(_01376_),
    .S(_00833_),
    .X(_01377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13194_ (.A0(_00705_),
    .A1(_00714_),
    .S(_00840_),
    .X(_01376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13195_ (.A0(_00688_),
    .A1(_00697_),
    .S(_00840_),
    .X(_01375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13196_ (.A0(_01372_),
    .A1(_01373_),
    .S(_00833_),
    .X(_01374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13197_ (.A0(_00671_),
    .A1(_00680_),
    .S(_00840_),
    .X(_01373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13198_ (.A0(_00654_),
    .A1(_00663_),
    .S(_00840_),
    .X(_01372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13199_ (.A0(_01368_),
    .A1(_01369_),
    .S(_00833_),
    .X(_01370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13200_ (.A0(_00637_),
    .A1(_00646_),
    .S(_00840_),
    .X(_01369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13201_ (.A0(_00620_),
    .A1(_00629_),
    .S(_00840_),
    .X(_01368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13202_ (.A0(_00603_),
    .A1(_00612_),
    .S(_00840_),
    .X(_01366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13203_ (.A0(_01357_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_01358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13204_ (.A0(_01355_),
    .A1(_01262_),
    .S(_00008_),
    .X(_01356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13205_ (.A0(_01353_),
    .A1(\design_top.IDATA[18] ),
    .S(_00008_),
    .X(_01354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13206_ (.A0(_01351_),
    .A1(\design_top.IDATA[17] ),
    .S(_00008_),
    .X(_01352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13207_ (.A0(_01349_),
    .A1(\design_top.IDATA[16] ),
    .S(_00008_),
    .X(_01350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13208_ (.A0(_01347_),
    .A1(\design_top.IDATA[15] ),
    .S(_00008_),
    .X(_01348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13209_ (.A0(_01345_),
    .A1(\design_top.IDATA[14] ),
    .S(_00008_),
    .X(_01346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13210_ (.A0(_01343_),
    .A1(\design_top.IDATA[13] ),
    .S(_00008_),
    .X(_01344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13211_ (.A0(_01340_),
    .A1(\design_top.IDATA[12] ),
    .S(_00008_),
    .X(_01341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13212_ (.A0(_01341_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_01342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13213_ (.A0(\design_top.ROMFF[11] ),
    .A1(\design_top.ROMFF2[11] ),
    .S(\design_top.HLT2 ),
    .X(_01315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13214_ (.A0(\design_top.ROMFF[29] ),
    .A1(\design_top.ROMFF2[29] ),
    .S(\design_top.HLT2 ),
    .X(_01298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13215_ (.A0(\design_top.ROMFF[28] ),
    .A1(\design_top.ROMFF2[28] ),
    .S(\design_top.HLT2 ),
    .X(_01294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13216_ (.A0(\design_top.ROMFF[27] ),
    .A1(\design_top.ROMFF2[27] ),
    .S(\design_top.HLT2 ),
    .X(_01290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13217_ (.A0(\design_top.ROMFF[26] ),
    .A1(\design_top.ROMFF2[26] ),
    .S(\design_top.HLT2 ),
    .X(_01286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13218_ (.A0(\design_top.ROMFF[25] ),
    .A1(\design_top.ROMFF2[25] ),
    .S(\design_top.HLT2 ),
    .X(_01282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13219_ (.A0(\design_top.ROMFF[24] ),
    .A1(\design_top.ROMFF2[24] ),
    .S(\design_top.HLT2 ),
    .X(_01278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13220_ (.A0(\design_top.ROMFF[19] ),
    .A1(\design_top.ROMFF2[19] ),
    .S(\design_top.HLT2 ),
    .X(_01262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13221_ (.A0(\design_top.ROMFF[6] ),
    .A1(\design_top.ROMFF2[6] ),
    .S(\design_top.HLT2 ),
    .X(_00906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13222_ (.A0(\design_top.ROMFF[5] ),
    .A1(\design_top.ROMFF2[5] ),
    .S(\design_top.HLT2 ),
    .X(_00905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13223_ (.A0(\design_top.ROMFF[4] ),
    .A1(\design_top.ROMFF2[4] ),
    .S(\design_top.HLT2 ),
    .X(_00904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13224_ (.A0(_00868_),
    .A1(_00895_),
    .S(_00537_),
    .X(_00896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13225_ (.A0(_00896_),
    .A1(_00865_),
    .S(_00866_),
    .X(_00897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13226_ (.A0(_00897_),
    .A1(_00863_),
    .S(_00864_),
    .X(_00898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13227_ (.A0(_00898_),
    .A1(_00842_),
    .S(_00533_),
    .X(_00899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13228_ (.A0(_00899_),
    .A1(_00841_),
    .S(_00538_),
    .X(_00900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13229_ (.A0(_00748_),
    .A1(\design_top.core0.UIMM[12] ),
    .S(\design_top.core0.XMCC ),
    .X(_00862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13230_ (.A0(_00739_),
    .A1(\design_top.core0.UIMM[13] ),
    .S(\design_top.core0.XMCC ),
    .X(_00861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13231_ (.A0(_00731_),
    .A1(\design_top.core0.UIMM[14] ),
    .S(\design_top.core0.XMCC ),
    .X(_00860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13232_ (.A0(_00576_),
    .A1(\design_top.core0.UIMM[15] ),
    .S(\design_top.core0.XMCC ),
    .X(_00859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13233_ (.A0(_00719_),
    .A1(\design_top.core0.UIMM[16] ),
    .S(\design_top.core0.XMCC ),
    .X(_00858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13234_ (.A0(_00710_),
    .A1(\design_top.core0.UIMM[17] ),
    .S(\design_top.core0.XMCC ),
    .X(_00857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13235_ (.A0(_00702_),
    .A1(\design_top.core0.UIMM[18] ),
    .S(\design_top.core0.XMCC ),
    .X(_00856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13236_ (.A0(_00693_),
    .A1(\design_top.core0.UIMM[19] ),
    .S(\design_top.core0.XMCC ),
    .X(_00855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13237_ (.A0(_00685_),
    .A1(\design_top.core0.UIMM[20] ),
    .S(\design_top.core0.XMCC ),
    .X(_00854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13238_ (.A0(_00676_),
    .A1(\design_top.core0.UIMM[21] ),
    .S(\design_top.core0.XMCC ),
    .X(_00853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13239_ (.A0(_00668_),
    .A1(\design_top.core0.UIMM[22] ),
    .S(\design_top.core0.XMCC ),
    .X(_00852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13240_ (.A0(_00659_),
    .A1(\design_top.core0.UIMM[23] ),
    .S(\design_top.core0.XMCC ),
    .X(_00851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13241_ (.A0(_00651_),
    .A1(\design_top.core0.UIMM[24] ),
    .S(\design_top.core0.XMCC ),
    .X(_00850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13242_ (.A0(_00642_),
    .A1(\design_top.core0.UIMM[25] ),
    .S(\design_top.core0.XMCC ),
    .X(_00849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13243_ (.A0(_00634_),
    .A1(\design_top.core0.UIMM[26] ),
    .S(\design_top.core0.XMCC ),
    .X(_00848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13244_ (.A0(_00625_),
    .A1(\design_top.core0.UIMM[27] ),
    .S(\design_top.core0.XMCC ),
    .X(_00847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13245_ (.A0(_00617_),
    .A1(\design_top.core0.UIMM[28] ),
    .S(\design_top.core0.XMCC ),
    .X(_00846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13246_ (.A0(_00608_),
    .A1(\design_top.core0.UIMM[29] ),
    .S(\design_top.core0.XMCC ),
    .X(_00845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13247_ (.A0(_00599_),
    .A1(\design_top.core0.UIMM[30] ),
    .S(\design_top.core0.XMCC ),
    .X(_00844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13248_ (.A0(_00582_),
    .A1(\design_top.core0.UIMM[31] ),
    .S(\design_top.core0.XMCC ),
    .X(_00843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13249_ (.A0(_00839_),
    .A1(\design_top.core0.SIMM[0] ),
    .S(\design_top.core0.XMCC ),
    .X(_00840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13250_ (.A0(_00832_),
    .A1(\design_top.core0.SIMM[1] ),
    .S(\design_top.core0.XMCC ),
    .X(_00833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13251_ (.A0(_00824_),
    .A1(\design_top.core0.SIMM[2] ),
    .S(\design_top.core0.XMCC ),
    .X(_00825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13252_ (.A0(_00815_),
    .A1(\design_top.core0.SIMM[3] ),
    .S(\design_top.core0.XMCC ),
    .X(_00816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13253_ (.A0(_00807_),
    .A1(\design_top.core0.SIMM[4] ),
    .S(\design_top.core0.XMCC ),
    .X(_00808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13254_ (.A0(_00798_),
    .A1(\design_top.core0.SIMM[5] ),
    .S(\design_top.core0.XMCC ),
    .X(_00799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13255_ (.A0(_00791_),
    .A1(\design_top.core0.SIMM[6] ),
    .S(\design_top.core0.XMCC ),
    .X(_00792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13256_ (.A0(_00570_),
    .A1(\design_top.core0.SIMM[7] ),
    .S(\design_top.core0.XMCC ),
    .X(_00783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13257_ (.A0(_00780_),
    .A1(\design_top.core0.SIMM[8] ),
    .S(\design_top.core0.XMCC ),
    .X(_00781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13258_ (.A0(_00771_),
    .A1(\design_top.core0.SIMM[9] ),
    .S(\design_top.core0.XMCC ),
    .X(_00772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13259_ (.A0(_00764_),
    .A1(\design_top.core0.SIMM[10] ),
    .S(\design_top.core0.XMCC ),
    .X(_00765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13260_ (.A0(_00755_),
    .A1(\design_top.core0.SIMM[11] ),
    .S(\design_top.core0.XMCC ),
    .X(_00756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13261_ (.A0(_00748_),
    .A1(\design_top.core0.SIMM[12] ),
    .S(\design_top.core0.XMCC ),
    .X(_00749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13262_ (.A0(_00739_),
    .A1(\design_top.core0.SIMM[13] ),
    .S(\design_top.core0.XMCC ),
    .X(_00740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13263_ (.A0(_00731_),
    .A1(\design_top.core0.SIMM[14] ),
    .S(\design_top.core0.XMCC ),
    .X(_00732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13264_ (.A0(_00576_),
    .A1(\design_top.core0.SIMM[15] ),
    .S(\design_top.core0.XMCC ),
    .X(_00723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13265_ (.A0(_00719_),
    .A1(\design_top.core0.SIMM[16] ),
    .S(\design_top.core0.XMCC ),
    .X(_00720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13266_ (.A0(_00710_),
    .A1(\design_top.core0.SIMM[17] ),
    .S(\design_top.core0.XMCC ),
    .X(_00711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13267_ (.A0(_00702_),
    .A1(\design_top.core0.SIMM[18] ),
    .S(\design_top.core0.XMCC ),
    .X(_00703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13268_ (.A0(_00693_),
    .A1(\design_top.core0.SIMM[19] ),
    .S(\design_top.core0.XMCC ),
    .X(_00694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13269_ (.A0(_00685_),
    .A1(\design_top.core0.SIMM[20] ),
    .S(\design_top.core0.XMCC ),
    .X(_00686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13270_ (.A0(_00676_),
    .A1(\design_top.core0.SIMM[21] ),
    .S(\design_top.core0.XMCC ),
    .X(_00677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13271_ (.A0(_00668_),
    .A1(\design_top.core0.SIMM[22] ),
    .S(\design_top.core0.XMCC ),
    .X(_00669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13272_ (.A0(_00659_),
    .A1(\design_top.core0.SIMM[23] ),
    .S(\design_top.core0.XMCC ),
    .X(_00660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13273_ (.A0(_00651_),
    .A1(\design_top.core0.SIMM[24] ),
    .S(\design_top.core0.XMCC ),
    .X(_00652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13274_ (.A0(_00642_),
    .A1(\design_top.core0.SIMM[25] ),
    .S(\design_top.core0.XMCC ),
    .X(_00643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13275_ (.A0(_00634_),
    .A1(\design_top.core0.SIMM[26] ),
    .S(\design_top.core0.XMCC ),
    .X(_00635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13276_ (.A0(_00625_),
    .A1(\design_top.core0.SIMM[27] ),
    .S(\design_top.core0.XMCC ),
    .X(_00626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13277_ (.A0(_00617_),
    .A1(\design_top.core0.SIMM[28] ),
    .S(\design_top.core0.XMCC ),
    .X(_00618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13278_ (.A0(_00608_),
    .A1(\design_top.core0.SIMM[29] ),
    .S(\design_top.core0.XMCC ),
    .X(_00609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13279_ (.A0(_00599_),
    .A1(\design_top.core0.SIMM[30] ),
    .S(\design_top.core0.XMCC ),
    .X(_00600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13280_ (.A0(_00582_),
    .A1(\design_top.core0.SIMM[31] ),
    .S(\design_top.core0.XMCC ),
    .X(_00591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13281_ (.A0(_00552_),
    .A1(_00536_),
    .S(_00539_),
    .X(_00553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13282_ (.A0(_00548_),
    .A1(_00544_),
    .S(_00539_),
    .X(_00549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13283_ (.A0(_00546_),
    .A1(_00544_),
    .S(_00539_),
    .X(_00547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13284_ (.A0(_00541_),
    .A1(_00536_),
    .S(_00539_),
    .X(_00542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13285_ (.A0(_00338_),
    .A1(_00341_),
    .S(_00304_),
    .X(_00342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13286_ (.A0(_00339_),
    .A1(_00340_),
    .S(_00303_),
    .X(_00341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13287_ (.A0(_00336_),
    .A1(_00337_),
    .S(_00303_),
    .X(_00338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13288_ (.A0(_00329_),
    .A1(_00332_),
    .S(_00304_),
    .X(_00333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13289_ (.A0(_00330_),
    .A1(_00331_),
    .S(_00303_),
    .X(_00332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13290_ (.A0(_00327_),
    .A1(_00328_),
    .S(_00303_),
    .X(_00329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13291_ (.A0(_00320_),
    .A1(_00323_),
    .S(_00304_),
    .X(_00324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13292_ (.A0(_00321_),
    .A1(_00322_),
    .S(_00303_),
    .X(_00323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13293_ (.A0(_00318_),
    .A1(_00319_),
    .S(_00303_),
    .X(_00320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13294_ (.A0(_00313_),
    .A1(_00316_),
    .S(_00304_),
    .X(_00317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13295_ (.A0(_00314_),
    .A1(_00315_),
    .S(_00303_),
    .X(_00316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13296_ (.A0(_00311_),
    .A1(_00312_),
    .S(_00303_),
    .X(_00313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13297_ (.A0(_02507_),
    .A1(_02508_),
    .S(_00589_),
    .X(_02509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13298_ (.A0(_02509_),
    .A1(_02506_),
    .S(_00901_),
    .X(_00097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13299_ (.A0(_02503_),
    .A1(_02504_),
    .S(_00589_),
    .X(_02505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13300_ (.A0(_02505_),
    .A1(_02502_),
    .S(_00901_),
    .X(_00096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13301_ (.A0(_02499_),
    .A1(_02500_),
    .S(_00589_),
    .X(_02501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13302_ (.A0(_02501_),
    .A1(_02498_),
    .S(_00901_),
    .X(_00095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13303_ (.A0(_02495_),
    .A1(_02496_),
    .S(_00589_),
    .X(_02497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13304_ (.A0(_02497_),
    .A1(_02494_),
    .S(_00901_),
    .X(_00094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13305_ (.A0(_02491_),
    .A1(_02492_),
    .S(_00589_),
    .X(_02493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13306_ (.A0(_02493_),
    .A1(_02490_),
    .S(_00901_),
    .X(_00093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13307_ (.A0(_02487_),
    .A1(_02488_),
    .S(_00589_),
    .X(_02489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13308_ (.A0(_02489_),
    .A1(_02486_),
    .S(_00901_),
    .X(_00092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13309_ (.A0(_02483_),
    .A1(_02484_),
    .S(_00589_),
    .X(_02485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13310_ (.A0(_02485_),
    .A1(_02482_),
    .S(_00901_),
    .X(_00091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13311_ (.A0(_02479_),
    .A1(_02480_),
    .S(_00589_),
    .X(_02481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13312_ (.A0(_02481_),
    .A1(_02478_),
    .S(_00901_),
    .X(_00090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13313_ (.A0(_02475_),
    .A1(_02476_),
    .S(_00589_),
    .X(_02477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13314_ (.A0(_02477_),
    .A1(_02474_),
    .S(_00901_),
    .X(_00089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13315_ (.A0(_02471_),
    .A1(_02472_),
    .S(_00589_),
    .X(_02473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13316_ (.A0(_02473_),
    .A1(_02470_),
    .S(_00901_),
    .X(_00088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13317_ (.A0(_02467_),
    .A1(_02468_),
    .S(_00589_),
    .X(_02469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13318_ (.A0(_02469_),
    .A1(_02466_),
    .S(_00901_),
    .X(_00087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13319_ (.A0(_02463_),
    .A1(_02464_),
    .S(_00589_),
    .X(_02465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13320_ (.A0(_02465_),
    .A1(_02462_),
    .S(_00901_),
    .X(_00086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13321_ (.A0(_02459_),
    .A1(_02460_),
    .S(_00589_),
    .X(_02461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13322_ (.A0(_02461_),
    .A1(_02458_),
    .S(_00901_),
    .X(_00085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13323_ (.A0(_02455_),
    .A1(_02456_),
    .S(_00589_),
    .X(_02457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13324_ (.A0(_02457_),
    .A1(_02454_),
    .S(_00901_),
    .X(_00084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13325_ (.A0(_02451_),
    .A1(_02452_),
    .S(_00589_),
    .X(_02453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13326_ (.A0(_02453_),
    .A1(_02450_),
    .S(_00901_),
    .X(_00083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13327_ (.A0(_02447_),
    .A1(_02448_),
    .S(_00589_),
    .X(_02449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13328_ (.A0(_02449_),
    .A1(_02446_),
    .S(_00901_),
    .X(_00082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13329_ (.A0(_02443_),
    .A1(_02444_),
    .S(_00589_),
    .X(_02445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13330_ (.A0(_02445_),
    .A1(_02442_),
    .S(_00901_),
    .X(_00081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13331_ (.A0(_02439_),
    .A1(_02440_),
    .S(_00589_),
    .X(_02441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13332_ (.A0(_02441_),
    .A1(_02438_),
    .S(_00901_),
    .X(_00080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13333_ (.A0(_02435_),
    .A1(_02436_),
    .S(_00589_),
    .X(_02437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13334_ (.A0(_02437_),
    .A1(_02434_),
    .S(_00901_),
    .X(_00079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13335_ (.A0(_02431_),
    .A1(_02432_),
    .S(_00589_),
    .X(_02433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13336_ (.A0(_02433_),
    .A1(_02430_),
    .S(_00901_),
    .X(_00108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13337_ (.A0(_02427_),
    .A1(_02428_),
    .S(_00589_),
    .X(_02429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13338_ (.A0(_02429_),
    .A1(_02426_),
    .S(_00901_),
    .X(_00107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13339_ (.A0(_02423_),
    .A1(_02424_),
    .S(_00589_),
    .X(_02425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13340_ (.A0(_02425_),
    .A1(_02422_),
    .S(_00901_),
    .X(_00106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13341_ (.A0(_02419_),
    .A1(_02420_),
    .S(_00589_),
    .X(_02421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13342_ (.A0(_02421_),
    .A1(_02418_),
    .S(_00901_),
    .X(_00105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13343_ (.A0(_02416_),
    .A1(_02415_),
    .S(_00589_),
    .X(_02417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13344_ (.A0(_02417_),
    .A1(_02414_),
    .S(_00901_),
    .X(_00104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13345_ (.A0(_02412_),
    .A1(_00543_),
    .S(_00589_),
    .X(_02413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13346_ (.A0(_02413_),
    .A1(_02411_),
    .S(_00901_),
    .X(_00103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13347_ (.A0(_02409_),
    .A1(\design_top.DADDR[3] ),
    .S(_00589_),
    .X(_02410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13348_ (.A0(_02410_),
    .A1(_02408_),
    .S(_00901_),
    .X(_00102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13349_ (.A0(_02406_),
    .A1(\design_top.DADDR[2] ),
    .S(_00589_),
    .X(_02407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13350_ (.A0(_02407_),
    .A1(_02405_),
    .S(_00901_),
    .X(_00099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13351_ (.A0(_02050_),
    .A1(_02051_),
    .S(\design_top.core0.XRES ),
    .X(_00045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13352_ (.A0(_01514_),
    .A1(_01513_),
    .S(_00309_),
    .X(_00011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13353_ (.A0(_01512_),
    .A1(_00903_),
    .S(_00902_),
    .X(_00078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13354_ (.A0(\design_top.IDATA[15] ),
    .A1(\design_top.core0.S1PTR[0] ),
    .S(\design_top.HLT ),
    .X(_00000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13355_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_00565_),
    .X(_00196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13356_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_00565_),
    .X(_00195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13357_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_00565_),
    .X(_00194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13358_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_00565_),
    .X(_00193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13359_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_00565_),
    .X(_00192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13360_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_00565_),
    .X(_00191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13361_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_00565_),
    .X(_00190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13362_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_00565_),
    .X(_00189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13363_ (.A0(_01337_),
    .A1(\design_top.IDATA[20] ),
    .S(_00008_),
    .X(_01338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13364_ (.A0(_01338_),
    .A1(\design_top.IDATA[7] ),
    .S(_00009_),
    .X(_01339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13365_ (.A0(_01339_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13366_ (.A0(_01334_),
    .A1(\design_top.IDATA[30] ),
    .S(_00008_),
    .X(_01335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13367_ (.A0(_01335_),
    .A1(\design_top.IDATA[30] ),
    .S(_00009_),
    .X(_01336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13368_ (.A0(_01336_),
    .A1(\design_top.IDATA[30] ),
    .S(_00010_),
    .X(_00048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13369_ (.A0(_01331_),
    .A1(_01298_),
    .S(_00008_),
    .X(_01332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13370_ (.A0(_01332_),
    .A1(_01298_),
    .S(_00009_),
    .X(_01333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13371_ (.A0(_01333_),
    .A1(_01298_),
    .S(_00010_),
    .X(_00077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13372_ (.A0(_01328_),
    .A1(_01294_),
    .S(_00008_),
    .X(_01329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13373_ (.A0(_01329_),
    .A1(_01294_),
    .S(_00009_),
    .X(_01330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13374_ (.A0(_01330_),
    .A1(_01294_),
    .S(_00010_),
    .X(_00076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13375_ (.A0(_01325_),
    .A1(_01290_),
    .S(_00008_),
    .X(_01326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13376_ (.A0(_01326_),
    .A1(_01290_),
    .S(_00009_),
    .X(_01327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13377_ (.A0(_01327_),
    .A1(_01290_),
    .S(_00010_),
    .X(_00075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13378_ (.A0(_01322_),
    .A1(_01286_),
    .S(_00008_),
    .X(_01323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13379_ (.A0(_01323_),
    .A1(_01286_),
    .S(_00009_),
    .X(_01324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13380_ (.A0(_01324_),
    .A1(_01286_),
    .S(_00010_),
    .X(_00074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13381_ (.A0(_01319_),
    .A1(_01282_),
    .S(_00008_),
    .X(_01320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13382_ (.A0(_01320_),
    .A1(_01282_),
    .S(_00009_),
    .X(_01321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13383_ (.A0(_01321_),
    .A1(_01282_),
    .S(_00010_),
    .X(_00073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13384_ (.A0(_01316_),
    .A1(_01278_),
    .S(_00008_),
    .X(_01317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13385_ (.A0(_01317_),
    .A1(_01315_),
    .S(_00009_),
    .X(_01318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13386_ (.A0(_01318_),
    .A1(_01315_),
    .S(_00010_),
    .X(_00072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13387_ (.A0(_01312_),
    .A1(\design_top.IDATA[23] ),
    .S(_00008_),
    .X(_01313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13388_ (.A0(_01313_),
    .A1(\design_top.IDATA[10] ),
    .S(_00009_),
    .X(_01314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13389_ (.A0(_01314_),
    .A1(\design_top.IDATA[10] ),
    .S(_00010_),
    .X(_00071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13390_ (.A0(_01309_),
    .A1(\design_top.IDATA[22] ),
    .S(_00008_),
    .X(_01310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13391_ (.A0(_01310_),
    .A1(\design_top.IDATA[9] ),
    .S(_00009_),
    .X(_01311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13392_ (.A0(_01311_),
    .A1(\design_top.IDATA[9] ),
    .S(_00010_),
    .X(_00069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13393_ (.A0(_01306_),
    .A1(\design_top.IDATA[21] ),
    .S(_00008_),
    .X(_01307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13394_ (.A0(_01307_),
    .A1(\design_top.IDATA[8] ),
    .S(_00009_),
    .X(_01308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13395_ (.A0(_01308_),
    .A1(\design_top.IDATA[8] ),
    .S(_00010_),
    .X(_00058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13396_ (.A0(_01305_),
    .A1(\design_top.IDATA[7] ),
    .S(_00010_),
    .X(_00047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13397_ (.A0(\design_top.IDATA[16] ),
    .A1(\design_top.core0.S1PTR[1] ),
    .S(\design_top.HLT ),
    .X(_00001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13398_ (.A0(\design_top.IDATA[30] ),
    .A1(\design_top.IDATA[31] ),
    .S(_01240_),
    .X(_01302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13399_ (.A0(_01302_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_01303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13400_ (.A0(_01303_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_01304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13401_ (.A0(_01304_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13402_ (.A0(_01298_),
    .A1(\design_top.IDATA[31] ),
    .S(_01240_),
    .X(_01299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13403_ (.A0(_01299_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_01300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13404_ (.A0(_01300_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_01301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13405_ (.A0(_01301_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13406_ (.A0(_01294_),
    .A1(\design_top.IDATA[31] ),
    .S(_01240_),
    .X(_01295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13407_ (.A0(_01295_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_01296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13408_ (.A0(_01296_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_01297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13409_ (.A0(_01297_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13410_ (.A0(_01290_),
    .A1(\design_top.IDATA[31] ),
    .S(_01240_),
    .X(_01291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13411_ (.A0(_01291_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_01292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13412_ (.A0(_01292_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_01293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13413_ (.A0(_01293_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13414_ (.A0(_01286_),
    .A1(\design_top.IDATA[31] ),
    .S(_01240_),
    .X(_01287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13415_ (.A0(_01287_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_01288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13416_ (.A0(_01288_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_01289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13417_ (.A0(_01289_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13418_ (.A0(_01282_),
    .A1(\design_top.IDATA[31] ),
    .S(_01240_),
    .X(_01283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13419_ (.A0(_01283_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_01284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13420_ (.A0(_01284_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_01285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13421_ (.A0(_01285_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13422_ (.A0(_01278_),
    .A1(\design_top.IDATA[31] ),
    .S(_01240_),
    .X(_01279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13423_ (.A0(_01279_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_01280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13424_ (.A0(_01280_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_01281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13425_ (.A0(_01281_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13426_ (.A0(\design_top.IDATA[23] ),
    .A1(\design_top.IDATA[31] ),
    .S(_01240_),
    .X(_01275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13427_ (.A0(_01275_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_01276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13428_ (.A0(_01276_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_01277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13429_ (.A0(_01277_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13430_ (.A0(\design_top.IDATA[22] ),
    .A1(\design_top.IDATA[31] ),
    .S(_01240_),
    .X(_01272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13431_ (.A0(_01272_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_01273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13432_ (.A0(_01273_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_01274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13433_ (.A0(_01274_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13434_ (.A0(\design_top.IDATA[21] ),
    .A1(\design_top.IDATA[31] ),
    .S(_01240_),
    .X(_01269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13435_ (.A0(_01269_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_01270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13436_ (.A0(_01270_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_01271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13437_ (.A0(_01271_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13438_ (.A0(\design_top.IDATA[20] ),
    .A1(\design_top.IDATA[31] ),
    .S(_01240_),
    .X(_01266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13439_ (.A0(_01266_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_01267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13440_ (.A0(_01267_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_01268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13441_ (.A0(_01268_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13442_ (.A0(_01262_),
    .A1(\design_top.IDATA[31] ),
    .S(_01240_),
    .X(_01263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13443_ (.A0(_01263_),
    .A1(_01262_),
    .S(_00008_),
    .X(_01264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13444_ (.A0(_01264_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_01265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13445_ (.A0(_01265_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13446_ (.A0(\design_top.IDATA[18] ),
    .A1(\design_top.IDATA[31] ),
    .S(_01240_),
    .X(_01259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13447_ (.A0(_01259_),
    .A1(\design_top.IDATA[18] ),
    .S(_00008_),
    .X(_01260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13448_ (.A0(_01260_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_01261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13449_ (.A0(_01261_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13450_ (.A0(\design_top.IDATA[17] ),
    .A1(\design_top.IDATA[31] ),
    .S(_01240_),
    .X(_01256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13451_ (.A0(_01256_),
    .A1(\design_top.IDATA[17] ),
    .S(_00008_),
    .X(_01257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13452_ (.A0(_01257_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_01258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13453_ (.A0(_01258_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13454_ (.A0(\design_top.IDATA[16] ),
    .A1(\design_top.IDATA[31] ),
    .S(_01240_),
    .X(_01253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13455_ (.A0(_01253_),
    .A1(\design_top.IDATA[16] ),
    .S(_00008_),
    .X(_01254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13456_ (.A0(_01254_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_01255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13457_ (.A0(_01255_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13458_ (.A0(\design_top.IDATA[15] ),
    .A1(\design_top.IDATA[31] ),
    .S(_01240_),
    .X(_01250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13459_ (.A0(_01250_),
    .A1(\design_top.IDATA[15] ),
    .S(_00008_),
    .X(_01251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13460_ (.A0(_01251_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_01252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13461_ (.A0(_01252_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13462_ (.A0(\design_top.IDATA[14] ),
    .A1(\design_top.IDATA[31] ),
    .S(_01240_),
    .X(_01247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13463_ (.A0(_01247_),
    .A1(\design_top.IDATA[14] ),
    .S(_00008_),
    .X(_01248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13464_ (.A0(_01248_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_01249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13465_ (.A0(_01249_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13466_ (.A0(\design_top.IDATA[13] ),
    .A1(\design_top.IDATA[31] ),
    .S(_01240_),
    .X(_01244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13467_ (.A0(_01244_),
    .A1(\design_top.IDATA[13] ),
    .S(_00008_),
    .X(_01245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13468_ (.A0(_01245_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_01246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13469_ (.A0(_01246_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13470_ (.A0(\design_top.IDATA[12] ),
    .A1(\design_top.IDATA[31] ),
    .S(_01240_),
    .X(_01241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13471_ (.A0(_01241_),
    .A1(\design_top.IDATA[12] ),
    .S(_00008_),
    .X(_01242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13472_ (.A0(_01242_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_01243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13473_ (.A0(_01243_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13474_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_00585_),
    .X(_00180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13475_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_00585_),
    .X(_00179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13476_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_00585_),
    .X(_00178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13477_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_00585_),
    .X(_00177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13478_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_00585_),
    .X(_00176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13479_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_00585_),
    .X(_00175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13480_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_00585_),
    .X(_00174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13481_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_00585_),
    .X(_00173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13482_ (.A0(\design_top.IDATA[22] ),
    .A1(\design_top.core0.S2PTR[2] ),
    .S(\design_top.HLT ),
    .X(_00006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13483_ (.A0(\design_top.IDATA[23] ),
    .A1(\design_top.core0.S2PTR[3] ),
    .S(\design_top.HLT ),
    .X(_00007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13484_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_00558_),
    .X(_00260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13485_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_00558_),
    .X(_00259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13486_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_00558_),
    .X(_00258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13487_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_00558_),
    .X(_00257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13488_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_00558_),
    .X(_00256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13489_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_00558_),
    .X(_00255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13490_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_00558_),
    .X(_00254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13491_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_00558_),
    .X(_00253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13492_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_00557_),
    .X(_00268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13493_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_00557_),
    .X(_00267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13494_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_00557_),
    .X(_00266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13495_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_00557_),
    .X(_00265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13496_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_00557_),
    .X(_00264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13497_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_00557_),
    .X(_00263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13498_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_00557_),
    .X(_00262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13499_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_00557_),
    .X(_00261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13500_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_00556_),
    .X(_00276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13501_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_00556_),
    .X(_00275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13502_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_00556_),
    .X(_00274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13503_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_00556_),
    .X(_00273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13504_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_00556_),
    .X(_00272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13505_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_00556_),
    .X(_00271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13506_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_00556_),
    .X(_00270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13507_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_00556_),
    .X(_00269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13508_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_00555_),
    .X(_00284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13509_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_00555_),
    .X(_00283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13510_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_00555_),
    .X(_00282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13511_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_00555_),
    .X(_00281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13512_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_00555_),
    .X(_00280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13513_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_00555_),
    .X(_00279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13514_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_00555_),
    .X(_00278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13515_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_00555_),
    .X(_00277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13516_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_00554_),
    .X(_00292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13517_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_00554_),
    .X(_00291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13518_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_00554_),
    .X(_00290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13519_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_00554_),
    .X(_00289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13520_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_00554_),
    .X(_00288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13521_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_00554_),
    .X(_00287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13522_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_00554_),
    .X(_00286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13523_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_00554_),
    .X(_00285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13524_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_00550_),
    .X(_00300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13525_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_00550_),
    .X(_00299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13526_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_00550_),
    .X(_00298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13527_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_00550_),
    .X(_00297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13528_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_00550_),
    .X(_00296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13529_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_00550_),
    .X(_00295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13530_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_00550_),
    .X(_00294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13531_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_00550_),
    .X(_00293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13532_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_00561_),
    .X(_00236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13533_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_00561_),
    .X(_00235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13534_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_00561_),
    .X(_00234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13535_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_00561_),
    .X(_00233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13536_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_00561_),
    .X(_00232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13537_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_00561_),
    .X(_00231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13538_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_00561_),
    .X(_00230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13539_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_00561_),
    .X(_00229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13540_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_00564_),
    .X(_00204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13541_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_00564_),
    .X(_00203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13542_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_00564_),
    .X(_00202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13543_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_00564_),
    .X(_00201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13544_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_00564_),
    .X(_00200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13545_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_00564_),
    .X(_00199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13546_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_00564_),
    .X(_00198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13547_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_00564_),
    .X(_00197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13548_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_00563_),
    .X(_00212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13549_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_00563_),
    .X(_00211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13550_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_00563_),
    .X(_00210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13551_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_00563_),
    .X(_00209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13552_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_00563_),
    .X(_00208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13553_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_00563_),
    .X(_00207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13554_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_00563_),
    .X(_00206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13555_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_00563_),
    .X(_00205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13556_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_00587_),
    .X(_00220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13557_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_00587_),
    .X(_00219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13558_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_00587_),
    .X(_00218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13559_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_00587_),
    .X(_00217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13560_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_00587_),
    .X(_00216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13561_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_00587_),
    .X(_00215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13562_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_00587_),
    .X(_00214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13563_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_00587_),
    .X(_00213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13564_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_00562_),
    .X(_00228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13565_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_00562_),
    .X(_00227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13566_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_00562_),
    .X(_00226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13567_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_00562_),
    .X(_00225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13568_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_00562_),
    .X(_00224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13569_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_00562_),
    .X(_00223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13570_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_00562_),
    .X(_00222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13571_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_00562_),
    .X(_00221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13572_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_00560_),
    .X(_00244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13573_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_00560_),
    .X(_00243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13574_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_00560_),
    .X(_00242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13575_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_00560_),
    .X(_00241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13576_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_00560_),
    .X(_00240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13577_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_00560_),
    .X(_00239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13578_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_00560_),
    .X(_00238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13579_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_00560_),
    .X(_00237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13580_ (.A0(_01111_),
    .A1(io_out[12]),
    .S(_00588_),
    .X(_00012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13581_ (.A0(\design_top.IDATA[18] ),
    .A1(\design_top.core0.S1PTR[3] ),
    .S(\design_top.HLT ),
    .X(_00003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13582_ (.A0(\design_top.IDATA[21] ),
    .A1(\design_top.core0.S2PTR[1] ),
    .S(\design_top.HLT ),
    .X(_00005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13583_ (.A0(_01110_),
    .A1(\design_top.IOMUX[3][31] ),
    .S(_00345_),
    .X(_00037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13584_ (.A0(_01109_),
    .A1(\design_top.IOMUX[3][30] ),
    .S(_00345_),
    .X(_00036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13585_ (.A0(_01108_),
    .A1(\design_top.IOMUX[3][29] ),
    .S(_00345_),
    .X(_00034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13586_ (.A0(_01107_),
    .A1(\design_top.IOMUX[3][28] ),
    .S(_00345_),
    .X(_00033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13587_ (.A0(_01106_),
    .A1(\design_top.IOMUX[3][27] ),
    .S(_00345_),
    .X(_00032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13588_ (.A0(_01105_),
    .A1(\design_top.IOMUX[3][26] ),
    .S(_00345_),
    .X(_00031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13589_ (.A0(_01104_),
    .A1(\design_top.IOMUX[3][25] ),
    .S(_00345_),
    .X(_00030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13590_ (.A0(_01103_),
    .A1(\design_top.IOMUX[3][24] ),
    .S(_00345_),
    .X(_00029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13591_ (.A0(_01102_),
    .A1(\design_top.IOMUX[3][23] ),
    .S(_00345_),
    .X(_00028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13592_ (.A0(_01101_),
    .A1(\design_top.IOMUX[3][22] ),
    .S(_00345_),
    .X(_00027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13593_ (.A0(_01100_),
    .A1(\design_top.IOMUX[3][21] ),
    .S(_00345_),
    .X(_00026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13594_ (.A0(_01099_),
    .A1(\design_top.IOMUX[3][20] ),
    .S(_00345_),
    .X(_00025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13595_ (.A0(_01098_),
    .A1(\design_top.IOMUX[3][19] ),
    .S(_00345_),
    .X(_00023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13596_ (.A0(_01097_),
    .A1(\design_top.IOMUX[3][18] ),
    .S(_00345_),
    .X(_00022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13597_ (.A0(_01096_),
    .A1(\design_top.IOMUX[3][17] ),
    .S(_00345_),
    .X(_00021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13598_ (.A0(_01095_),
    .A1(\design_top.IOMUX[3][16] ),
    .S(_00345_),
    .X(_00020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13599_ (.A0(_01094_),
    .A1(\design_top.IOMUX[3][15] ),
    .S(_00345_),
    .X(_00019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13600_ (.A0(_01093_),
    .A1(\design_top.IOMUX[3][14] ),
    .S(_00345_),
    .X(_00018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13601_ (.A0(_01092_),
    .A1(\design_top.IOMUX[3][13] ),
    .S(_00345_),
    .X(_00017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13602_ (.A0(_01091_),
    .A1(\design_top.IOMUX[3][12] ),
    .S(_00345_),
    .X(_00016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13603_ (.A0(_01090_),
    .A1(\design_top.IOMUX[3][11] ),
    .S(_00345_),
    .X(_00015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13604_ (.A0(_01089_),
    .A1(\design_top.IOMUX[3][10] ),
    .S(_00345_),
    .X(_00014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13605_ (.A0(_01088_),
    .A1(\design_top.IOMUX[3][9] ),
    .S(_00345_),
    .X(_00044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13606_ (.A0(_01087_),
    .A1(\design_top.IOMUX[3][8] ),
    .S(_00345_),
    .X(_00043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13607_ (.A0(_01086_),
    .A1(\design_top.IOMUX[3][7] ),
    .S(_00345_),
    .X(_00042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13608_ (.A0(_01085_),
    .A1(\design_top.IOMUX[3][6] ),
    .S(_00345_),
    .X(_00041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13609_ (.A0(_01084_),
    .A1(\design_top.IOMUX[3][5] ),
    .S(_00345_),
    .X(_00040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13610_ (.A0(_01083_),
    .A1(\design_top.IOMUX[3][4] ),
    .S(_00345_),
    .X(_00039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13611_ (.A0(_01082_),
    .A1(\design_top.IOMUX[3][3] ),
    .S(_00345_),
    .X(_00038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13612_ (.A0(_01081_),
    .A1(\design_top.IOMUX[3][2] ),
    .S(_00345_),
    .X(_00035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13613_ (.A0(_01080_),
    .A1(\design_top.IOMUX[3][1] ),
    .S(_00345_),
    .X(_00024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13614_ (.A0(_01079_),
    .A1(\design_top.IOMUX[3][0] ),
    .S(_00345_),
    .X(_00013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13615_ (.A0(\design_top.IDATA[17] ),
    .A1(\design_top.core0.S1PTR[2] ),
    .S(\design_top.HLT ),
    .X(_00002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13616_ (.A0(\design_top.IDATA[20] ),
    .A1(\design_top.core0.S2PTR[0] ),
    .S(\design_top.HLT ),
    .X(_00004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13617_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_00559_),
    .X(_00252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13618_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_00559_),
    .X(_00251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13619_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_00559_),
    .X(_00250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13620_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_00559_),
    .X(_00249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13621_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_00559_),
    .X(_00248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13622_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_00559_),
    .X(_00247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13623_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_00559_),
    .X(_00246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13624_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_00559_),
    .X(_00245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13625_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_00584_),
    .X(_00188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13626_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_00584_),
    .X(_00187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13627_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_00584_),
    .X(_00186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13628_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_00584_),
    .X(_00185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13629_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_00584_),
    .X(_00184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13630_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_00584_),
    .X(_00183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13631_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_00584_),
    .X(_00182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13632_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_00584_),
    .X(_00181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13633_ (.A0(_00920_),
    .A1(\design_top.DADDR[31] ),
    .S(_00589_),
    .X(_00921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13634_ (.A0(_00921_),
    .A1(_00918_),
    .S(_00901_),
    .X(_00101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13635_ (.A0(_00915_),
    .A1(_00916_),
    .S(_00589_),
    .X(_00917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13636_ (.A0(_00917_),
    .A1(_00913_),
    .S(_00901_),
    .X(_00100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13637_ (.A0(_00910_),
    .A1(_00911_),
    .S(_00589_),
    .X(_00912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _13638_ (.A0(_00912_),
    .A1(_00908_),
    .S(_00901_),
    .X(_00098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13639_ (.A0(\design_top.uart0.UART_XFIFO[0] ),
    .A1(\design_top.uart0.UART_XFIFO[1] ),
    .A2(\design_top.uart0.UART_XFIFO[2] ),
    .A3(\design_top.uart0.UART_XFIFO[3] ),
    .S0(\design_top.uart0.UART_XSTATE[0] ),
    .S1(\design_top.uart0.UART_XSTATE[1] ),
    .X(_00923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13640_ (.A0(\design_top.uart0.UART_XFIFO[4] ),
    .A1(\design_top.uart0.UART_XFIFO[5] ),
    .A2(\design_top.uart0.UART_XFIFO[6] ),
    .A3(\design_top.uart0.UART_XFIFO[7] ),
    .S0(\design_top.uart0.UART_XSTATE[0] ),
    .S1(\design_top.uart0.UART_XSTATE[1] ),
    .X(_00924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13641_ (.A0(_02397_),
    .A1(_00602_),
    .A2(_01432_),
    .A3(_02398_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_02399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13642_ (.A0(_02393_),
    .A1(_02390_),
    .A2(_02384_),
    .A3(_02385_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_02394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13643_ (.A0(_02377_),
    .A1(_00611_),
    .A2(_01432_),
    .A3(_02378_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_02379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13644_ (.A0(_02373_),
    .A1(_02370_),
    .A2(_02365_),
    .A3(_02366_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_02374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13645_ (.A0(_02357_),
    .A1(_02343_),
    .A2(_01432_),
    .A3(_02358_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_02359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13646_ (.A0(_02353_),
    .A1(_02350_),
    .A2(_02344_),
    .A3(_02345_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_02354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13647_ (.A0(_02335_),
    .A1(_00628_),
    .A2(_01432_),
    .A3(_02336_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_02337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13648_ (.A0(_02331_),
    .A1(_02328_),
    .A2(_02324_),
    .A3(_02325_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_02332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13649_ (.A0(_02316_),
    .A1(_02302_),
    .A2(_01432_),
    .A3(_02317_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_02318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13650_ (.A0(_02312_),
    .A1(_02309_),
    .A2(_02303_),
    .A3(_02304_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_02313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13651_ (.A0(_02294_),
    .A1(_00645_),
    .A2(_01432_),
    .A3(_02295_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_02296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13652_ (.A0(_02290_),
    .A1(_02287_),
    .A2(_02282_),
    .A3(_02283_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_02291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13653_ (.A0(_02274_),
    .A1(_02260_),
    .A2(_01432_),
    .A3(_02275_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_02276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13654_ (.A0(_02270_),
    .A1(_02267_),
    .A2(_02261_),
    .A3(_02262_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_02271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13655_ (.A0(_02252_),
    .A1(_00662_),
    .A2(_01432_),
    .A3(_02253_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_02254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13656_ (.A0(_02248_),
    .A1(_02245_),
    .A2(_02242_),
    .A3(_02243_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_02249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13657_ (.A0(_02234_),
    .A1(_02220_),
    .A2(_01432_),
    .A3(_02235_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_02236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13658_ (.A0(_02230_),
    .A1(_02227_),
    .A2(_02221_),
    .A3(_02222_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_02231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13659_ (.A0(_02212_),
    .A1(_00679_),
    .A2(_01432_),
    .A3(_02213_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_02214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13660_ (.A0(_02208_),
    .A1(_02205_),
    .A2(_02200_),
    .A3(_02201_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_02209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13661_ (.A0(_02192_),
    .A1(_02178_),
    .A2(_01432_),
    .A3(_02193_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_02194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13662_ (.A0(_02188_),
    .A1(_02185_),
    .A2(_02179_),
    .A3(_02180_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_02189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13663_ (.A0(_02170_),
    .A1(_00696_),
    .A2(_01432_),
    .A3(_02171_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_02172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13664_ (.A0(_02166_),
    .A1(_02163_),
    .A2(_02159_),
    .A3(_02160_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_02167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13665_ (.A0(_02151_),
    .A1(_02136_),
    .A2(_01432_),
    .A3(_02152_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_02153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13666_ (.A0(_02147_),
    .A1(_02144_),
    .A2(_02138_),
    .A3(_02139_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_02148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13667_ (.A0(_02128_),
    .A1(_00713_),
    .A2(_01432_),
    .A3(_02129_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_02130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13668_ (.A0(_02124_),
    .A1(_02121_),
    .A2(_02116_),
    .A3(_02117_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_02125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13669_ (.A0(_02108_),
    .A1(_02094_),
    .A2(_01432_),
    .A3(_02109_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_02110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13670_ (.A0(_02104_),
    .A1(_02101_),
    .A2(_02095_),
    .A3(_02096_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_02105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13671_ (.A0(_02086_),
    .A1(_00725_),
    .A2(_01432_),
    .A3(_02087_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_02088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13672_ (.A0(_02081_),
    .A1(_01403_),
    .A2(_02081_),
    .A3(_00381_),
    .S0(_00808_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_02082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13673_ (.A0(_02082_),
    .A1(_02080_),
    .A2(_02078_),
    .A3(_02079_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_02083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13674_ (.A0(_02069_),
    .A1(_02053_),
    .A2(_01432_),
    .A3(_02071_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_02072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13675_ (.A0(_02062_),
    .A1(_02063_),
    .A2(_02062_),
    .A3(_02064_),
    .S0(_00808_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_02065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13676_ (.A0(_02065_),
    .A1(_02061_),
    .A2(_02055_),
    .A3(_02056_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_02066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13677_ (.A0(_02042_),
    .A1(_00742_),
    .A2(_01432_),
    .A3(_02044_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_02045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13678_ (.A0(_02035_),
    .A1(_02036_),
    .A2(_02035_),
    .A3(_02037_),
    .S0(_00808_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_02038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13679_ (.A0(_02038_),
    .A1(_02034_),
    .A2(_02029_),
    .A3(_02030_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_02039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13680_ (.A0(_02020_),
    .A1(_02005_),
    .A2(_01432_),
    .A3(_02022_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_02023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13681_ (.A0(_02013_),
    .A1(_02014_),
    .A2(_02013_),
    .A3(_02015_),
    .S0(_00808_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_02016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13682_ (.A0(_02016_),
    .A1(_02012_),
    .A2(_02006_),
    .A3(_02007_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_02017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13683_ (.A0(_01996_),
    .A1(_00758_),
    .A2(_01432_),
    .A3(_01998_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_01999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13684_ (.A0(_01989_),
    .A1(_01990_),
    .A2(_01989_),
    .A3(_01991_),
    .S0(_00808_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13685_ (.A0(_01992_),
    .A1(_01988_),
    .A2(_01984_),
    .A3(_01985_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_01993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13686_ (.A0(_01975_),
    .A1(_01960_),
    .A2(_01432_),
    .A3(_01977_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_01978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13687_ (.A0(_01968_),
    .A1(_01969_),
    .A2(_01968_),
    .A3(_01970_),
    .S0(_00808_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13688_ (.A0(_01971_),
    .A1(_01967_),
    .A2(_01961_),
    .A3(_01962_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_01972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13689_ (.A0(_01951_),
    .A1(_00774_),
    .A2(_01432_),
    .A3(_01953_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_01954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13690_ (.A0(_01944_),
    .A1(_01945_),
    .A2(_01944_),
    .A3(_01946_),
    .S0(_00808_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13691_ (.A0(_01947_),
    .A1(_01943_),
    .A2(_01938_),
    .A3(_01939_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_01948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13692_ (.A0(_01929_),
    .A1(_01914_),
    .A2(_01432_),
    .A3(_01931_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_01932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13693_ (.A0(_01922_),
    .A1(_01923_),
    .A2(_01922_),
    .A3(_01924_),
    .S0(_00808_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13694_ (.A0(_01925_),
    .A1(_01921_),
    .A2(_01915_),
    .A3(_01916_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_01926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13695_ (.A0(_01905_),
    .A1(_00785_),
    .A2(_01431_),
    .A3(_01907_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_01908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13696_ (.A0(_01897_),
    .A1(_01899_),
    .A2(_01897_),
    .A3(_01900_),
    .S0(_00808_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13697_ (.A0(_01901_),
    .A1(_01894_),
    .A2(_01891_),
    .A3(_01892_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_01902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13698_ (.A0(_01866_),
    .A1(_01845_),
    .A2(_01884_),
    .A3(_01875_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_01885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13699_ (.A0(_01856_),
    .A1(_01859_),
    .A2(_01856_),
    .A3(_01861_),
    .S0(_00808_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13700_ (.A0(_01862_),
    .A1(_01853_),
    .A2(_01847_),
    .A3(_01848_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_01863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13701_ (.A0(_01820_),
    .A1(_00801_),
    .A2(_01838_),
    .A3(_01829_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_01839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13702_ (.A0(_01810_),
    .A1(_01813_),
    .A2(_01810_),
    .A3(_01815_),
    .S0(_00808_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13703_ (.A0(_01816_),
    .A1(_01807_),
    .A2(_01802_),
    .A3(_01803_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_01817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13704_ (.A0(_01778_),
    .A1(_01758_),
    .A2(_01795_),
    .A3(_01786_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_01796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13705_ (.A0(_01768_),
    .A1(_01771_),
    .A2(_01768_),
    .A3(_01773_),
    .S0(_00808_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13706_ (.A0(_01774_),
    .A1(_01765_),
    .A2(_01759_),
    .A3(_01760_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_01775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13707_ (.A0(_01734_),
    .A1(_00818_),
    .A2(_01751_),
    .A3(_01742_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_01752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13708_ (.A0(_01721_),
    .A1(_01727_),
    .A2(_01721_),
    .A3(_01729_),
    .S0(_00808_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13709_ (.A0(_01730_),
    .A1(_01714_),
    .A2(_01710_),
    .A3(_01711_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_01731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13710_ (.A0(_01685_),
    .A1(_01655_),
    .A2(_01703_),
    .A3(_01694_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_01704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13711_ (.A0(_01670_),
    .A1(_01677_),
    .A2(_01670_),
    .A3(_01680_),
    .S0(_00808_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13712_ (.A0(_01681_),
    .A1(_01663_),
    .A2(_01657_),
    .A3(_01658_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_01682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13713_ (.A0(_01630_),
    .A1(_01361_),
    .A2(_01648_),
    .A3(_01638_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_01649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13714_ (.A0(_01608_),
    .A1(_01622_),
    .A2(_01608_),
    .A3(_01625_),
    .S0(_00808_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13715_ (.A0(_01626_),
    .A1(_01593_),
    .A2(_01588_),
    .A3(_01589_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_01627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13716_ (.A0(_01560_),
    .A1(_01516_),
    .A2(_01580_),
    .A3(_01569_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_01581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13717_ (.A0(_01411_),
    .A1(_00593_),
    .A2(_01432_),
    .A3(_01422_),
    .S0(_07035_),
    .S1(io_out[12]),
    .X(_01433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13718_ (.A0(_01405_),
    .A1(_01399_),
    .A2(_01362_),
    .A3(_01364_),
    .S0(_07036_),
    .S1(_00537_),
    .X(_01406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13719_ (.A0(\design_top.core0.REG2[0][0] ),
    .A1(\design_top.core0.REG2[1][0] ),
    .A2(\design_top.core0.REG2[2][0] ),
    .A3(\design_top.core0.REG2[3][0] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13720_ (.A0(\design_top.core0.REG2[4][0] ),
    .A1(\design_top.core0.REG2[5][0] ),
    .A2(\design_top.core0.REG2[6][0] ),
    .A3(\design_top.core0.REG2[7][0] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13721_ (.A0(\design_top.core0.REG2[8][0] ),
    .A1(\design_top.core0.REG2[9][0] ),
    .A2(\design_top.core0.REG2[10][0] ),
    .A3(\design_top.core0.REG2[11][0] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13722_ (.A0(\design_top.core0.REG2[12][0] ),
    .A1(\design_top.core0.REG2[13][0] ),
    .A2(\design_top.core0.REG2[14][0] ),
    .A3(\design_top.core0.REG2[15][0] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13723_ (.A0(_00835_),
    .A1(_00836_),
    .A2(_00837_),
    .A3(_00838_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13724_ (.A0(\design_top.core0.REG2[0][1] ),
    .A1(\design_top.core0.REG2[1][1] ),
    .A2(\design_top.core0.REG2[2][1] ),
    .A3(\design_top.core0.REG2[3][1] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13725_ (.A0(\design_top.core0.REG2[4][1] ),
    .A1(\design_top.core0.REG2[5][1] ),
    .A2(\design_top.core0.REG2[6][1] ),
    .A3(\design_top.core0.REG2[7][1] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13726_ (.A0(\design_top.core0.REG2[8][1] ),
    .A1(\design_top.core0.REG2[9][1] ),
    .A2(\design_top.core0.REG2[10][1] ),
    .A3(\design_top.core0.REG2[11][1] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13727_ (.A0(\design_top.core0.REG2[12][1] ),
    .A1(\design_top.core0.REG2[13][1] ),
    .A2(\design_top.core0.REG2[14][1] ),
    .A3(\design_top.core0.REG2[15][1] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13728_ (.A0(_00828_),
    .A1(_00829_),
    .A2(_00830_),
    .A3(_00831_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13729_ (.A0(\design_top.core0.REG2[0][2] ),
    .A1(\design_top.core0.REG2[1][2] ),
    .A2(\design_top.core0.REG2[2][2] ),
    .A3(\design_top.core0.REG2[3][2] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13730_ (.A0(\design_top.core0.REG2[4][2] ),
    .A1(\design_top.core0.REG2[5][2] ),
    .A2(\design_top.core0.REG2[6][2] ),
    .A3(\design_top.core0.REG2[7][2] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13731_ (.A0(\design_top.core0.REG2[8][2] ),
    .A1(\design_top.core0.REG2[9][2] ),
    .A2(\design_top.core0.REG2[10][2] ),
    .A3(\design_top.core0.REG2[11][2] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13732_ (.A0(\design_top.core0.REG2[12][2] ),
    .A1(\design_top.core0.REG2[13][2] ),
    .A2(\design_top.core0.REG2[14][2] ),
    .A3(\design_top.core0.REG2[15][2] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13733_ (.A0(_00820_),
    .A1(_00821_),
    .A2(_00822_),
    .A3(_00823_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13734_ (.A0(\design_top.core0.REG2[0][3] ),
    .A1(\design_top.core0.REG2[1][3] ),
    .A2(\design_top.core0.REG2[2][3] ),
    .A3(\design_top.core0.REG2[3][3] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13735_ (.A0(\design_top.core0.REG2[4][3] ),
    .A1(\design_top.core0.REG2[5][3] ),
    .A2(\design_top.core0.REG2[6][3] ),
    .A3(\design_top.core0.REG2[7][3] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13736_ (.A0(\design_top.core0.REG2[8][3] ),
    .A1(\design_top.core0.REG2[9][3] ),
    .A2(\design_top.core0.REG2[10][3] ),
    .A3(\design_top.core0.REG2[11][3] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13737_ (.A0(\design_top.core0.REG2[12][3] ),
    .A1(\design_top.core0.REG2[13][3] ),
    .A2(\design_top.core0.REG2[14][3] ),
    .A3(\design_top.core0.REG2[15][3] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13738_ (.A0(_00811_),
    .A1(_00812_),
    .A2(_00813_),
    .A3(_00814_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13739_ (.A0(\design_top.core0.REG2[0][4] ),
    .A1(\design_top.core0.REG2[1][4] ),
    .A2(\design_top.core0.REG2[2][4] ),
    .A3(\design_top.core0.REG2[3][4] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13740_ (.A0(\design_top.core0.REG2[4][4] ),
    .A1(\design_top.core0.REG2[5][4] ),
    .A2(\design_top.core0.REG2[6][4] ),
    .A3(\design_top.core0.REG2[7][4] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13741_ (.A0(\design_top.core0.REG2[8][4] ),
    .A1(\design_top.core0.REG2[9][4] ),
    .A2(\design_top.core0.REG2[10][4] ),
    .A3(\design_top.core0.REG2[11][4] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13742_ (.A0(\design_top.core0.REG2[12][4] ),
    .A1(\design_top.core0.REG2[13][4] ),
    .A2(\design_top.core0.REG2[14][4] ),
    .A3(\design_top.core0.REG2[15][4] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13743_ (.A0(_00803_),
    .A1(_00804_),
    .A2(_00805_),
    .A3(_00806_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13744_ (.A0(\design_top.core0.REG2[0][5] ),
    .A1(\design_top.core0.REG2[1][5] ),
    .A2(\design_top.core0.REG2[2][5] ),
    .A3(\design_top.core0.REG2[3][5] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13745_ (.A0(\design_top.core0.REG2[4][5] ),
    .A1(\design_top.core0.REG2[5][5] ),
    .A2(\design_top.core0.REG2[6][5] ),
    .A3(\design_top.core0.REG2[7][5] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13746_ (.A0(\design_top.core0.REG2[8][5] ),
    .A1(\design_top.core0.REG2[9][5] ),
    .A2(\design_top.core0.REG2[10][5] ),
    .A3(\design_top.core0.REG2[11][5] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13747_ (.A0(\design_top.core0.REG2[12][5] ),
    .A1(\design_top.core0.REG2[13][5] ),
    .A2(\design_top.core0.REG2[14][5] ),
    .A3(\design_top.core0.REG2[15][5] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13748_ (.A0(_00794_),
    .A1(_00795_),
    .A2(_00796_),
    .A3(_00797_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13749_ (.A0(\design_top.core0.REG2[0][6] ),
    .A1(\design_top.core0.REG2[1][6] ),
    .A2(\design_top.core0.REG2[2][6] ),
    .A3(\design_top.core0.REG2[3][6] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13750_ (.A0(\design_top.core0.REG2[4][6] ),
    .A1(\design_top.core0.REG2[5][6] ),
    .A2(\design_top.core0.REG2[6][6] ),
    .A3(\design_top.core0.REG2[7][6] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13751_ (.A0(\design_top.core0.REG2[8][6] ),
    .A1(\design_top.core0.REG2[9][6] ),
    .A2(\design_top.core0.REG2[10][6] ),
    .A3(\design_top.core0.REG2[11][6] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13752_ (.A0(\design_top.core0.REG2[12][6] ),
    .A1(\design_top.core0.REG2[13][6] ),
    .A2(\design_top.core0.REG2[14][6] ),
    .A3(\design_top.core0.REG2[15][6] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13753_ (.A0(_00787_),
    .A1(_00788_),
    .A2(_00789_),
    .A3(_00790_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13754_ (.A0(\design_top.core0.REG2[0][8] ),
    .A1(\design_top.core0.REG2[1][8] ),
    .A2(\design_top.core0.REG2[2][8] ),
    .A3(\design_top.core0.REG2[3][8] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13755_ (.A0(\design_top.core0.REG2[4][8] ),
    .A1(\design_top.core0.REG2[5][8] ),
    .A2(\design_top.core0.REG2[6][8] ),
    .A3(\design_top.core0.REG2[7][8] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13756_ (.A0(\design_top.core0.REG2[8][8] ),
    .A1(\design_top.core0.REG2[9][8] ),
    .A2(\design_top.core0.REG2[10][8] ),
    .A3(\design_top.core0.REG2[11][8] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13757_ (.A0(\design_top.core0.REG2[12][8] ),
    .A1(\design_top.core0.REG2[13][8] ),
    .A2(\design_top.core0.REG2[14][8] ),
    .A3(\design_top.core0.REG2[15][8] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13758_ (.A0(_00776_),
    .A1(_00777_),
    .A2(_00778_),
    .A3(_00779_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13759_ (.A0(\design_top.core0.REG2[0][9] ),
    .A1(\design_top.core0.REG2[1][9] ),
    .A2(\design_top.core0.REG2[2][9] ),
    .A3(\design_top.core0.REG2[3][9] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13760_ (.A0(\design_top.core0.REG2[4][9] ),
    .A1(\design_top.core0.REG2[5][9] ),
    .A2(\design_top.core0.REG2[6][9] ),
    .A3(\design_top.core0.REG2[7][9] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13761_ (.A0(\design_top.core0.REG2[8][9] ),
    .A1(\design_top.core0.REG2[9][9] ),
    .A2(\design_top.core0.REG2[10][9] ),
    .A3(\design_top.core0.REG2[11][9] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13762_ (.A0(\design_top.core0.REG2[12][9] ),
    .A1(\design_top.core0.REG2[13][9] ),
    .A2(\design_top.core0.REG2[14][9] ),
    .A3(\design_top.core0.REG2[15][9] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13763_ (.A0(_00767_),
    .A1(_00768_),
    .A2(_00769_),
    .A3(_00770_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13764_ (.A0(\design_top.core0.REG2[0][10] ),
    .A1(\design_top.core0.REG2[1][10] ),
    .A2(\design_top.core0.REG2[2][10] ),
    .A3(\design_top.core0.REG2[3][10] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13765_ (.A0(\design_top.core0.REG2[4][10] ),
    .A1(\design_top.core0.REG2[5][10] ),
    .A2(\design_top.core0.REG2[6][10] ),
    .A3(\design_top.core0.REG2[7][10] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13766_ (.A0(\design_top.core0.REG2[8][10] ),
    .A1(\design_top.core0.REG2[9][10] ),
    .A2(\design_top.core0.REG2[10][10] ),
    .A3(\design_top.core0.REG2[11][10] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13767_ (.A0(\design_top.core0.REG2[12][10] ),
    .A1(\design_top.core0.REG2[13][10] ),
    .A2(\design_top.core0.REG2[14][10] ),
    .A3(\design_top.core0.REG2[15][10] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13768_ (.A0(_00760_),
    .A1(_00761_),
    .A2(_00762_),
    .A3(_00763_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13769_ (.A0(\design_top.core0.REG2[0][11] ),
    .A1(\design_top.core0.REG2[1][11] ),
    .A2(\design_top.core0.REG2[2][11] ),
    .A3(\design_top.core0.REG2[3][11] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13770_ (.A0(\design_top.core0.REG2[4][11] ),
    .A1(\design_top.core0.REG2[5][11] ),
    .A2(\design_top.core0.REG2[6][11] ),
    .A3(\design_top.core0.REG2[7][11] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13771_ (.A0(\design_top.core0.REG2[8][11] ),
    .A1(\design_top.core0.REG2[9][11] ),
    .A2(\design_top.core0.REG2[10][11] ),
    .A3(\design_top.core0.REG2[11][11] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13772_ (.A0(\design_top.core0.REG2[12][11] ),
    .A1(\design_top.core0.REG2[13][11] ),
    .A2(\design_top.core0.REG2[14][11] ),
    .A3(\design_top.core0.REG2[15][11] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13773_ (.A0(_00751_),
    .A1(_00752_),
    .A2(_00753_),
    .A3(_00754_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13774_ (.A0(\design_top.core0.REG2[0][12] ),
    .A1(\design_top.core0.REG2[1][12] ),
    .A2(\design_top.core0.REG2[2][12] ),
    .A3(\design_top.core0.REG2[3][12] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13775_ (.A0(\design_top.core0.REG2[4][12] ),
    .A1(\design_top.core0.REG2[5][12] ),
    .A2(\design_top.core0.REG2[6][12] ),
    .A3(\design_top.core0.REG2[7][12] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13776_ (.A0(\design_top.core0.REG2[8][12] ),
    .A1(\design_top.core0.REG2[9][12] ),
    .A2(\design_top.core0.REG2[10][12] ),
    .A3(\design_top.core0.REG2[11][12] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13777_ (.A0(\design_top.core0.REG2[12][12] ),
    .A1(\design_top.core0.REG2[13][12] ),
    .A2(\design_top.core0.REG2[14][12] ),
    .A3(\design_top.core0.REG2[15][12] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13778_ (.A0(_00744_),
    .A1(_00745_),
    .A2(_00746_),
    .A3(_00747_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13779_ (.A0(\design_top.core0.REG2[0][13] ),
    .A1(\design_top.core0.REG2[1][13] ),
    .A2(\design_top.core0.REG2[2][13] ),
    .A3(\design_top.core0.REG2[3][13] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13780_ (.A0(\design_top.core0.REG2[4][13] ),
    .A1(\design_top.core0.REG2[5][13] ),
    .A2(\design_top.core0.REG2[6][13] ),
    .A3(\design_top.core0.REG2[7][13] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13781_ (.A0(\design_top.core0.REG2[8][13] ),
    .A1(\design_top.core0.REG2[9][13] ),
    .A2(\design_top.core0.REG2[10][13] ),
    .A3(\design_top.core0.REG2[11][13] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13782_ (.A0(\design_top.core0.REG2[12][13] ),
    .A1(\design_top.core0.REG2[13][13] ),
    .A2(\design_top.core0.REG2[14][13] ),
    .A3(\design_top.core0.REG2[15][13] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13783_ (.A0(_00735_),
    .A1(_00736_),
    .A2(_00737_),
    .A3(_00738_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13784_ (.A0(\design_top.core0.REG2[0][14] ),
    .A1(\design_top.core0.REG2[1][14] ),
    .A2(\design_top.core0.REG2[2][14] ),
    .A3(\design_top.core0.REG2[3][14] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13785_ (.A0(\design_top.core0.REG2[4][14] ),
    .A1(\design_top.core0.REG2[5][14] ),
    .A2(\design_top.core0.REG2[6][14] ),
    .A3(\design_top.core0.REG2[7][14] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13786_ (.A0(\design_top.core0.REG2[8][14] ),
    .A1(\design_top.core0.REG2[9][14] ),
    .A2(\design_top.core0.REG2[10][14] ),
    .A3(\design_top.core0.REG2[11][14] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13787_ (.A0(\design_top.core0.REG2[12][14] ),
    .A1(\design_top.core0.REG2[13][14] ),
    .A2(\design_top.core0.REG2[14][14] ),
    .A3(\design_top.core0.REG2[15][14] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13788_ (.A0(_00727_),
    .A1(_00728_),
    .A2(_00729_),
    .A3(_00730_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13789_ (.A0(\design_top.core0.REG2[0][16] ),
    .A1(\design_top.core0.REG2[1][16] ),
    .A2(\design_top.core0.REG2[2][16] ),
    .A3(\design_top.core0.REG2[3][16] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13790_ (.A0(\design_top.core0.REG2[4][16] ),
    .A1(\design_top.core0.REG2[5][16] ),
    .A2(\design_top.core0.REG2[6][16] ),
    .A3(\design_top.core0.REG2[7][16] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13791_ (.A0(\design_top.core0.REG2[8][16] ),
    .A1(\design_top.core0.REG2[9][16] ),
    .A2(\design_top.core0.REG2[10][16] ),
    .A3(\design_top.core0.REG2[11][16] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13792_ (.A0(\design_top.core0.REG2[12][16] ),
    .A1(\design_top.core0.REG2[13][16] ),
    .A2(\design_top.core0.REG2[14][16] ),
    .A3(\design_top.core0.REG2[15][16] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13793_ (.A0(_00715_),
    .A1(_00716_),
    .A2(_00717_),
    .A3(_00718_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13794_ (.A0(\design_top.core0.REG2[0][17] ),
    .A1(\design_top.core0.REG2[1][17] ),
    .A2(\design_top.core0.REG2[2][17] ),
    .A3(\design_top.core0.REG2[3][17] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13795_ (.A0(\design_top.core0.REG2[4][17] ),
    .A1(\design_top.core0.REG2[5][17] ),
    .A2(\design_top.core0.REG2[6][17] ),
    .A3(\design_top.core0.REG2[7][17] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13796_ (.A0(\design_top.core0.REG2[8][17] ),
    .A1(\design_top.core0.REG2[9][17] ),
    .A2(\design_top.core0.REG2[10][17] ),
    .A3(\design_top.core0.REG2[11][17] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13797_ (.A0(\design_top.core0.REG2[12][17] ),
    .A1(\design_top.core0.REG2[13][17] ),
    .A2(\design_top.core0.REG2[14][17] ),
    .A3(\design_top.core0.REG2[15][17] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13798_ (.A0(_00706_),
    .A1(_00707_),
    .A2(_00708_),
    .A3(_00709_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13799_ (.A0(\design_top.core0.REG2[0][18] ),
    .A1(\design_top.core0.REG2[1][18] ),
    .A2(\design_top.core0.REG2[2][18] ),
    .A3(\design_top.core0.REG2[3][18] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13800_ (.A0(\design_top.core0.REG2[4][18] ),
    .A1(\design_top.core0.REG2[5][18] ),
    .A2(\design_top.core0.REG2[6][18] ),
    .A3(\design_top.core0.REG2[7][18] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13801_ (.A0(\design_top.core0.REG2[8][18] ),
    .A1(\design_top.core0.REG2[9][18] ),
    .A2(\design_top.core0.REG2[10][18] ),
    .A3(\design_top.core0.REG2[11][18] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13802_ (.A0(\design_top.core0.REG2[12][18] ),
    .A1(\design_top.core0.REG2[13][18] ),
    .A2(\design_top.core0.REG2[14][18] ),
    .A3(\design_top.core0.REG2[15][18] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13803_ (.A0(_00698_),
    .A1(_00699_),
    .A2(_00700_),
    .A3(_00701_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13804_ (.A0(\design_top.core0.REG2[0][19] ),
    .A1(\design_top.core0.REG2[1][19] ),
    .A2(\design_top.core0.REG2[2][19] ),
    .A3(\design_top.core0.REG2[3][19] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13805_ (.A0(\design_top.core0.REG2[4][19] ),
    .A1(\design_top.core0.REG2[5][19] ),
    .A2(\design_top.core0.REG2[6][19] ),
    .A3(\design_top.core0.REG2[7][19] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13806_ (.A0(\design_top.core0.REG2[8][19] ),
    .A1(\design_top.core0.REG2[9][19] ),
    .A2(\design_top.core0.REG2[10][19] ),
    .A3(\design_top.core0.REG2[11][19] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13807_ (.A0(\design_top.core0.REG2[12][19] ),
    .A1(\design_top.core0.REG2[13][19] ),
    .A2(\design_top.core0.REG2[14][19] ),
    .A3(\design_top.core0.REG2[15][19] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13808_ (.A0(_00689_),
    .A1(_00690_),
    .A2(_00691_),
    .A3(_00692_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13809_ (.A0(\design_top.core0.REG2[0][20] ),
    .A1(\design_top.core0.REG2[1][20] ),
    .A2(\design_top.core0.REG2[2][20] ),
    .A3(\design_top.core0.REG2[3][20] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13810_ (.A0(\design_top.core0.REG2[4][20] ),
    .A1(\design_top.core0.REG2[5][20] ),
    .A2(\design_top.core0.REG2[6][20] ),
    .A3(\design_top.core0.REG2[7][20] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13811_ (.A0(\design_top.core0.REG2[8][20] ),
    .A1(\design_top.core0.REG2[9][20] ),
    .A2(\design_top.core0.REG2[10][20] ),
    .A3(\design_top.core0.REG2[11][20] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13812_ (.A0(\design_top.core0.REG2[12][20] ),
    .A1(\design_top.core0.REG2[13][20] ),
    .A2(\design_top.core0.REG2[14][20] ),
    .A3(\design_top.core0.REG2[15][20] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13813_ (.A0(_00681_),
    .A1(_00682_),
    .A2(_00683_),
    .A3(_00684_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13814_ (.A0(\design_top.core0.REG2[0][21] ),
    .A1(\design_top.core0.REG2[1][21] ),
    .A2(\design_top.core0.REG2[2][21] ),
    .A3(\design_top.core0.REG2[3][21] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13815_ (.A0(\design_top.core0.REG2[4][21] ),
    .A1(\design_top.core0.REG2[5][21] ),
    .A2(\design_top.core0.REG2[6][21] ),
    .A3(\design_top.core0.REG2[7][21] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13816_ (.A0(\design_top.core0.REG2[8][21] ),
    .A1(\design_top.core0.REG2[9][21] ),
    .A2(\design_top.core0.REG2[10][21] ),
    .A3(\design_top.core0.REG2[11][21] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13817_ (.A0(\design_top.core0.REG2[12][21] ),
    .A1(\design_top.core0.REG2[13][21] ),
    .A2(\design_top.core0.REG2[14][21] ),
    .A3(\design_top.core0.REG2[15][21] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13818_ (.A0(_00672_),
    .A1(_00673_),
    .A2(_00674_),
    .A3(_00675_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13819_ (.A0(\design_top.core0.REG2[0][22] ),
    .A1(\design_top.core0.REG2[1][22] ),
    .A2(\design_top.core0.REG2[2][22] ),
    .A3(\design_top.core0.REG2[3][22] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13820_ (.A0(\design_top.core0.REG2[4][22] ),
    .A1(\design_top.core0.REG2[5][22] ),
    .A2(\design_top.core0.REG2[6][22] ),
    .A3(\design_top.core0.REG2[7][22] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13821_ (.A0(\design_top.core0.REG2[8][22] ),
    .A1(\design_top.core0.REG2[9][22] ),
    .A2(\design_top.core0.REG2[10][22] ),
    .A3(\design_top.core0.REG2[11][22] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13822_ (.A0(\design_top.core0.REG2[12][22] ),
    .A1(\design_top.core0.REG2[13][22] ),
    .A2(\design_top.core0.REG2[14][22] ),
    .A3(\design_top.core0.REG2[15][22] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13823_ (.A0(_00664_),
    .A1(_00665_),
    .A2(_00666_),
    .A3(_00667_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13824_ (.A0(\design_top.core0.REG2[0][23] ),
    .A1(\design_top.core0.REG2[1][23] ),
    .A2(\design_top.core0.REG2[2][23] ),
    .A3(\design_top.core0.REG2[3][23] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13825_ (.A0(\design_top.core0.REG2[4][23] ),
    .A1(\design_top.core0.REG2[5][23] ),
    .A2(\design_top.core0.REG2[6][23] ),
    .A3(\design_top.core0.REG2[7][23] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13826_ (.A0(\design_top.core0.REG2[8][23] ),
    .A1(\design_top.core0.REG2[9][23] ),
    .A2(\design_top.core0.REG2[10][23] ),
    .A3(\design_top.core0.REG2[11][23] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13827_ (.A0(\design_top.core0.REG2[12][23] ),
    .A1(\design_top.core0.REG2[13][23] ),
    .A2(\design_top.core0.REG2[14][23] ),
    .A3(\design_top.core0.REG2[15][23] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13828_ (.A0(_00655_),
    .A1(_00656_),
    .A2(_00657_),
    .A3(_00658_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13829_ (.A0(\design_top.core0.REG2[0][24] ),
    .A1(\design_top.core0.REG2[1][24] ),
    .A2(\design_top.core0.REG2[2][24] ),
    .A3(\design_top.core0.REG2[3][24] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13830_ (.A0(\design_top.core0.REG2[4][24] ),
    .A1(\design_top.core0.REG2[5][24] ),
    .A2(\design_top.core0.REG2[6][24] ),
    .A3(\design_top.core0.REG2[7][24] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13831_ (.A0(\design_top.core0.REG2[8][24] ),
    .A1(\design_top.core0.REG2[9][24] ),
    .A2(\design_top.core0.REG2[10][24] ),
    .A3(\design_top.core0.REG2[11][24] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13832_ (.A0(\design_top.core0.REG2[12][24] ),
    .A1(\design_top.core0.REG2[13][24] ),
    .A2(\design_top.core0.REG2[14][24] ),
    .A3(\design_top.core0.REG2[15][24] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13833_ (.A0(_00647_),
    .A1(_00648_),
    .A2(_00649_),
    .A3(_00650_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13834_ (.A0(\design_top.core0.REG2[0][25] ),
    .A1(\design_top.core0.REG2[1][25] ),
    .A2(\design_top.core0.REG2[2][25] ),
    .A3(\design_top.core0.REG2[3][25] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13835_ (.A0(\design_top.core0.REG2[4][25] ),
    .A1(\design_top.core0.REG2[5][25] ),
    .A2(\design_top.core0.REG2[6][25] ),
    .A3(\design_top.core0.REG2[7][25] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13836_ (.A0(\design_top.core0.REG2[8][25] ),
    .A1(\design_top.core0.REG2[9][25] ),
    .A2(\design_top.core0.REG2[10][25] ),
    .A3(\design_top.core0.REG2[11][25] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13837_ (.A0(\design_top.core0.REG2[12][25] ),
    .A1(\design_top.core0.REG2[13][25] ),
    .A2(\design_top.core0.REG2[14][25] ),
    .A3(\design_top.core0.REG2[15][25] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13838_ (.A0(_00638_),
    .A1(_00639_),
    .A2(_00640_),
    .A3(_00641_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13839_ (.A0(\design_top.core0.REG2[0][26] ),
    .A1(\design_top.core0.REG2[1][26] ),
    .A2(\design_top.core0.REG2[2][26] ),
    .A3(\design_top.core0.REG2[3][26] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13840_ (.A0(\design_top.core0.REG2[4][26] ),
    .A1(\design_top.core0.REG2[5][26] ),
    .A2(\design_top.core0.REG2[6][26] ),
    .A3(\design_top.core0.REG2[7][26] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13841_ (.A0(\design_top.core0.REG2[8][26] ),
    .A1(\design_top.core0.REG2[9][26] ),
    .A2(\design_top.core0.REG2[10][26] ),
    .A3(\design_top.core0.REG2[11][26] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13842_ (.A0(\design_top.core0.REG2[12][26] ),
    .A1(\design_top.core0.REG2[13][26] ),
    .A2(\design_top.core0.REG2[14][26] ),
    .A3(\design_top.core0.REG2[15][26] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13843_ (.A0(_00630_),
    .A1(_00631_),
    .A2(_00632_),
    .A3(_00633_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13844_ (.A0(\design_top.core0.REG2[0][27] ),
    .A1(\design_top.core0.REG2[1][27] ),
    .A2(\design_top.core0.REG2[2][27] ),
    .A3(\design_top.core0.REG2[3][27] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13845_ (.A0(\design_top.core0.REG2[4][27] ),
    .A1(\design_top.core0.REG2[5][27] ),
    .A2(\design_top.core0.REG2[6][27] ),
    .A3(\design_top.core0.REG2[7][27] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13846_ (.A0(\design_top.core0.REG2[8][27] ),
    .A1(\design_top.core0.REG2[9][27] ),
    .A2(\design_top.core0.REG2[10][27] ),
    .A3(\design_top.core0.REG2[11][27] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13847_ (.A0(\design_top.core0.REG2[12][27] ),
    .A1(\design_top.core0.REG2[13][27] ),
    .A2(\design_top.core0.REG2[14][27] ),
    .A3(\design_top.core0.REG2[15][27] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13848_ (.A0(_00621_),
    .A1(_00622_),
    .A2(_00623_),
    .A3(_00624_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13849_ (.A0(\design_top.core0.REG2[0][28] ),
    .A1(\design_top.core0.REG2[1][28] ),
    .A2(\design_top.core0.REG2[2][28] ),
    .A3(\design_top.core0.REG2[3][28] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13850_ (.A0(\design_top.core0.REG2[4][28] ),
    .A1(\design_top.core0.REG2[5][28] ),
    .A2(\design_top.core0.REG2[6][28] ),
    .A3(\design_top.core0.REG2[7][28] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13851_ (.A0(\design_top.core0.REG2[8][28] ),
    .A1(\design_top.core0.REG2[9][28] ),
    .A2(\design_top.core0.REG2[10][28] ),
    .A3(\design_top.core0.REG2[11][28] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13852_ (.A0(\design_top.core0.REG2[12][28] ),
    .A1(\design_top.core0.REG2[13][28] ),
    .A2(\design_top.core0.REG2[14][28] ),
    .A3(\design_top.core0.REG2[15][28] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13853_ (.A0(_00613_),
    .A1(_00614_),
    .A2(_00615_),
    .A3(_00616_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13854_ (.A0(\design_top.core0.REG2[0][29] ),
    .A1(\design_top.core0.REG2[1][29] ),
    .A2(\design_top.core0.REG2[2][29] ),
    .A3(\design_top.core0.REG2[3][29] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13855_ (.A0(\design_top.core0.REG2[4][29] ),
    .A1(\design_top.core0.REG2[5][29] ),
    .A2(\design_top.core0.REG2[6][29] ),
    .A3(\design_top.core0.REG2[7][29] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13856_ (.A0(\design_top.core0.REG2[8][29] ),
    .A1(\design_top.core0.REG2[9][29] ),
    .A2(\design_top.core0.REG2[10][29] ),
    .A3(\design_top.core0.REG2[11][29] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13857_ (.A0(\design_top.core0.REG2[12][29] ),
    .A1(\design_top.core0.REG2[13][29] ),
    .A2(\design_top.core0.REG2[14][29] ),
    .A3(\design_top.core0.REG2[15][29] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13858_ (.A0(_00604_),
    .A1(_00605_),
    .A2(_00606_),
    .A3(_00607_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13859_ (.A0(\design_top.core0.REG2[0][30] ),
    .A1(\design_top.core0.REG2[1][30] ),
    .A2(\design_top.core0.REG2[2][30] ),
    .A3(\design_top.core0.REG2[3][30] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13860_ (.A0(\design_top.core0.REG2[4][30] ),
    .A1(\design_top.core0.REG2[5][30] ),
    .A2(\design_top.core0.REG2[6][30] ),
    .A3(\design_top.core0.REG2[7][30] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13861_ (.A0(\design_top.core0.REG2[8][30] ),
    .A1(\design_top.core0.REG2[9][30] ),
    .A2(\design_top.core0.REG2[10][30] ),
    .A3(\design_top.core0.REG2[11][30] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13862_ (.A0(\design_top.core0.REG2[12][30] ),
    .A1(\design_top.core0.REG2[13][30] ),
    .A2(\design_top.core0.REG2[14][30] ),
    .A3(\design_top.core0.REG2[15][30] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13863_ (.A0(_00595_),
    .A1(_00596_),
    .A2(_00597_),
    .A3(_00598_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13864_ (.A0(\design_top.core0.REG2[0][31] ),
    .A1(\design_top.core0.REG2[1][31] ),
    .A2(\design_top.core0.REG2[2][31] ),
    .A3(\design_top.core0.REG2[3][31] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13865_ (.A0(\design_top.core0.REG2[4][31] ),
    .A1(\design_top.core0.REG2[5][31] ),
    .A2(\design_top.core0.REG2[6][31] ),
    .A3(\design_top.core0.REG2[7][31] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13866_ (.A0(\design_top.core0.REG2[8][31] ),
    .A1(\design_top.core0.REG2[9][31] ),
    .A2(\design_top.core0.REG2[10][31] ),
    .A3(\design_top.core0.REG2[11][31] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13867_ (.A0(\design_top.core0.REG2[12][31] ),
    .A1(\design_top.core0.REG2[13][31] ),
    .A2(\design_top.core0.REG2[14][31] ),
    .A3(\design_top.core0.REG2[15][31] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13868_ (.A0(_00578_),
    .A1(_00579_),
    .A2(_00580_),
    .A3(_00581_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13869_ (.A0(\design_top.core0.REG2[0][15] ),
    .A1(\design_top.core0.REG2[1][15] ),
    .A2(\design_top.core0.REG2[2][15] ),
    .A3(\design_top.core0.REG2[3][15] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13870_ (.A0(\design_top.core0.REG2[4][15] ),
    .A1(\design_top.core0.REG2[5][15] ),
    .A2(\design_top.core0.REG2[6][15] ),
    .A3(\design_top.core0.REG2[7][15] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13871_ (.A0(\design_top.core0.REG2[8][15] ),
    .A1(\design_top.core0.REG2[9][15] ),
    .A2(\design_top.core0.REG2[10][15] ),
    .A3(\design_top.core0.REG2[11][15] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13872_ (.A0(\design_top.core0.REG2[12][15] ),
    .A1(\design_top.core0.REG2[13][15] ),
    .A2(\design_top.core0.REG2[14][15] ),
    .A3(\design_top.core0.REG2[15][15] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13873_ (.A0(_00572_),
    .A1(_00573_),
    .A2(_00574_),
    .A3(_00575_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13874_ (.A0(\design_top.core0.REG2[0][7] ),
    .A1(\design_top.core0.REG2[1][7] ),
    .A2(\design_top.core0.REG2[2][7] ),
    .A3(\design_top.core0.REG2[3][7] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13875_ (.A0(\design_top.core0.REG2[4][7] ),
    .A1(\design_top.core0.REG2[5][7] ),
    .A2(\design_top.core0.REG2[6][7] ),
    .A3(\design_top.core0.REG2[7][7] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13876_ (.A0(\design_top.core0.REG2[8][7] ),
    .A1(\design_top.core0.REG2[9][7] ),
    .A2(\design_top.core0.REG2[10][7] ),
    .A3(\design_top.core0.REG2[11][7] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13877_ (.A0(\design_top.core0.REG2[12][7] ),
    .A1(\design_top.core0.REG2[13][7] ),
    .A2(\design_top.core0.REG2[14][7] ),
    .A3(\design_top.core0.REG2[15][7] ),
    .S0(_00305_),
    .S1(_00306_),
    .X(_00569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13878_ (.A0(_00566_),
    .A1(_00567_),
    .A2(_00568_),
    .A3(_00569_),
    .S0(_00307_),
    .S1(_00308_),
    .X(_00570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13879_ (.A0(\design_top.core0.REG1[0][6] ),
    .A1(\design_top.core0.REG1[1][6] ),
    .A2(\design_top.core0.REG1[2][6] ),
    .A3(\design_top.core0.REG1[3][6] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13880_ (.A0(\design_top.core0.REG1[4][6] ),
    .A1(\design_top.core0.REG1[5][6] ),
    .A2(\design_top.core0.REG1[6][6] ),
    .A3(\design_top.core0.REG1[7][6] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13881_ (.A0(\design_top.core0.REG1[8][6] ),
    .A1(\design_top.core0.REG1[9][6] ),
    .A2(\design_top.core0.REG1[10][6] ),
    .A3(\design_top.core0.REG1[11][6] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13882_ (.A0(\design_top.core0.REG1[12][6] ),
    .A1(\design_top.core0.REG1[13][6] ),
    .A2(\design_top.core0.REG1[14][6] ),
    .A3(\design_top.core0.REG1[15][6] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13883_ (.A0(_00526_),
    .A1(_00527_),
    .A2(_00528_),
    .A3(_00529_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13884_ (.A0(\design_top.core0.REG1[0][7] ),
    .A1(\design_top.core0.REG1[1][7] ),
    .A2(\design_top.core0.REG1[2][7] ),
    .A3(\design_top.core0.REG1[3][7] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13885_ (.A0(\design_top.core0.REG1[4][7] ),
    .A1(\design_top.core0.REG1[5][7] ),
    .A2(\design_top.core0.REG1[6][7] ),
    .A3(\design_top.core0.REG1[7][7] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13886_ (.A0(\design_top.core0.REG1[8][7] ),
    .A1(\design_top.core0.REG1[9][7] ),
    .A2(\design_top.core0.REG1[10][7] ),
    .A3(\design_top.core0.REG1[11][7] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13887_ (.A0(\design_top.core0.REG1[12][7] ),
    .A1(\design_top.core0.REG1[13][7] ),
    .A2(\design_top.core0.REG1[14][7] ),
    .A3(\design_top.core0.REG1[15][7] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13888_ (.A0(_00520_),
    .A1(_00521_),
    .A2(_00522_),
    .A3(_00523_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13889_ (.A0(\design_top.core0.REG1[0][8] ),
    .A1(\design_top.core0.REG1[1][8] ),
    .A2(\design_top.core0.REG1[2][8] ),
    .A3(\design_top.core0.REG1[3][8] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13890_ (.A0(\design_top.core0.REG1[4][8] ),
    .A1(\design_top.core0.REG1[5][8] ),
    .A2(\design_top.core0.REG1[6][8] ),
    .A3(\design_top.core0.REG1[7][8] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13891_ (.A0(\design_top.core0.REG1[8][8] ),
    .A1(\design_top.core0.REG1[9][8] ),
    .A2(\design_top.core0.REG1[10][8] ),
    .A3(\design_top.core0.REG1[11][8] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13892_ (.A0(\design_top.core0.REG1[12][8] ),
    .A1(\design_top.core0.REG1[13][8] ),
    .A2(\design_top.core0.REG1[14][8] ),
    .A3(\design_top.core0.REG1[15][8] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13893_ (.A0(_00514_),
    .A1(_00515_),
    .A2(_00516_),
    .A3(_00517_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13894_ (.A0(\design_top.core0.REG1[0][9] ),
    .A1(\design_top.core0.REG1[1][9] ),
    .A2(\design_top.core0.REG1[2][9] ),
    .A3(\design_top.core0.REG1[3][9] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13895_ (.A0(\design_top.core0.REG1[4][9] ),
    .A1(\design_top.core0.REG1[5][9] ),
    .A2(\design_top.core0.REG1[6][9] ),
    .A3(\design_top.core0.REG1[7][9] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13896_ (.A0(\design_top.core0.REG1[8][9] ),
    .A1(\design_top.core0.REG1[9][9] ),
    .A2(\design_top.core0.REG1[10][9] ),
    .A3(\design_top.core0.REG1[11][9] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13897_ (.A0(\design_top.core0.REG1[12][9] ),
    .A1(\design_top.core0.REG1[13][9] ),
    .A2(\design_top.core0.REG1[14][9] ),
    .A3(\design_top.core0.REG1[15][9] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13898_ (.A0(_00508_),
    .A1(_00509_),
    .A2(_00510_),
    .A3(_00511_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13899_ (.A0(\design_top.core0.REG1[0][10] ),
    .A1(\design_top.core0.REG1[1][10] ),
    .A2(\design_top.core0.REG1[2][10] ),
    .A3(\design_top.core0.REG1[3][10] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13900_ (.A0(\design_top.core0.REG1[4][10] ),
    .A1(\design_top.core0.REG1[5][10] ),
    .A2(\design_top.core0.REG1[6][10] ),
    .A3(\design_top.core0.REG1[7][10] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13901_ (.A0(\design_top.core0.REG1[8][10] ),
    .A1(\design_top.core0.REG1[9][10] ),
    .A2(\design_top.core0.REG1[10][10] ),
    .A3(\design_top.core0.REG1[11][10] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13902_ (.A0(\design_top.core0.REG1[12][10] ),
    .A1(\design_top.core0.REG1[13][10] ),
    .A2(\design_top.core0.REG1[14][10] ),
    .A3(\design_top.core0.REG1[15][10] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13903_ (.A0(_00502_),
    .A1(_00503_),
    .A2(_00504_),
    .A3(_00505_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13904_ (.A0(\design_top.core0.REG1[0][11] ),
    .A1(\design_top.core0.REG1[1][11] ),
    .A2(\design_top.core0.REG1[2][11] ),
    .A3(\design_top.core0.REG1[3][11] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13905_ (.A0(\design_top.core0.REG1[4][11] ),
    .A1(\design_top.core0.REG1[5][11] ),
    .A2(\design_top.core0.REG1[6][11] ),
    .A3(\design_top.core0.REG1[7][11] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13906_ (.A0(\design_top.core0.REG1[8][11] ),
    .A1(\design_top.core0.REG1[9][11] ),
    .A2(\design_top.core0.REG1[10][11] ),
    .A3(\design_top.core0.REG1[11][11] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13907_ (.A0(\design_top.core0.REG1[12][11] ),
    .A1(\design_top.core0.REG1[13][11] ),
    .A2(\design_top.core0.REG1[14][11] ),
    .A3(\design_top.core0.REG1[15][11] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13908_ (.A0(_00496_),
    .A1(_00497_),
    .A2(_00498_),
    .A3(_00499_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13909_ (.A0(\design_top.core0.REG1[0][12] ),
    .A1(\design_top.core0.REG1[1][12] ),
    .A2(\design_top.core0.REG1[2][12] ),
    .A3(\design_top.core0.REG1[3][12] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13910_ (.A0(\design_top.core0.REG1[4][12] ),
    .A1(\design_top.core0.REG1[5][12] ),
    .A2(\design_top.core0.REG1[6][12] ),
    .A3(\design_top.core0.REG1[7][12] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13911_ (.A0(\design_top.core0.REG1[8][12] ),
    .A1(\design_top.core0.REG1[9][12] ),
    .A2(\design_top.core0.REG1[10][12] ),
    .A3(\design_top.core0.REG1[11][12] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13912_ (.A0(\design_top.core0.REG1[12][12] ),
    .A1(\design_top.core0.REG1[13][12] ),
    .A2(\design_top.core0.REG1[14][12] ),
    .A3(\design_top.core0.REG1[15][12] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13913_ (.A0(_00490_),
    .A1(_00491_),
    .A2(_00492_),
    .A3(_00493_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13914_ (.A0(\design_top.core0.REG1[0][13] ),
    .A1(\design_top.core0.REG1[1][13] ),
    .A2(\design_top.core0.REG1[2][13] ),
    .A3(\design_top.core0.REG1[3][13] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13915_ (.A0(\design_top.core0.REG1[4][13] ),
    .A1(\design_top.core0.REG1[5][13] ),
    .A2(\design_top.core0.REG1[6][13] ),
    .A3(\design_top.core0.REG1[7][13] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13916_ (.A0(\design_top.core0.REG1[8][13] ),
    .A1(\design_top.core0.REG1[9][13] ),
    .A2(\design_top.core0.REG1[10][13] ),
    .A3(\design_top.core0.REG1[11][13] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13917_ (.A0(\design_top.core0.REG1[12][13] ),
    .A1(\design_top.core0.REG1[13][13] ),
    .A2(\design_top.core0.REG1[14][13] ),
    .A3(\design_top.core0.REG1[15][13] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13918_ (.A0(_00484_),
    .A1(_00485_),
    .A2(_00486_),
    .A3(_00487_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13919_ (.A0(\design_top.core0.REG1[0][14] ),
    .A1(\design_top.core0.REG1[1][14] ),
    .A2(\design_top.core0.REG1[2][14] ),
    .A3(\design_top.core0.REG1[3][14] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13920_ (.A0(\design_top.core0.REG1[4][14] ),
    .A1(\design_top.core0.REG1[5][14] ),
    .A2(\design_top.core0.REG1[6][14] ),
    .A3(\design_top.core0.REG1[7][14] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13921_ (.A0(\design_top.core0.REG1[8][14] ),
    .A1(\design_top.core0.REG1[9][14] ),
    .A2(\design_top.core0.REG1[10][14] ),
    .A3(\design_top.core0.REG1[11][14] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13922_ (.A0(\design_top.core0.REG1[12][14] ),
    .A1(\design_top.core0.REG1[13][14] ),
    .A2(\design_top.core0.REG1[14][14] ),
    .A3(\design_top.core0.REG1[15][14] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13923_ (.A0(_00478_),
    .A1(_00479_),
    .A2(_00480_),
    .A3(_00481_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13924_ (.A0(\design_top.core0.REG1[0][15] ),
    .A1(\design_top.core0.REG1[1][15] ),
    .A2(\design_top.core0.REG1[2][15] ),
    .A3(\design_top.core0.REG1[3][15] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13925_ (.A0(\design_top.core0.REG1[4][15] ),
    .A1(\design_top.core0.REG1[5][15] ),
    .A2(\design_top.core0.REG1[6][15] ),
    .A3(\design_top.core0.REG1[7][15] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13926_ (.A0(\design_top.core0.REG1[8][15] ),
    .A1(\design_top.core0.REG1[9][15] ),
    .A2(\design_top.core0.REG1[10][15] ),
    .A3(\design_top.core0.REG1[11][15] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13927_ (.A0(\design_top.core0.REG1[12][15] ),
    .A1(\design_top.core0.REG1[13][15] ),
    .A2(\design_top.core0.REG1[14][15] ),
    .A3(\design_top.core0.REG1[15][15] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13928_ (.A0(_00472_),
    .A1(_00473_),
    .A2(_00474_),
    .A3(_00475_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13929_ (.A0(\design_top.core0.REG1[0][16] ),
    .A1(\design_top.core0.REG1[1][16] ),
    .A2(\design_top.core0.REG1[2][16] ),
    .A3(\design_top.core0.REG1[3][16] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13930_ (.A0(\design_top.core0.REG1[4][16] ),
    .A1(\design_top.core0.REG1[5][16] ),
    .A2(\design_top.core0.REG1[6][16] ),
    .A3(\design_top.core0.REG1[7][16] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13931_ (.A0(\design_top.core0.REG1[8][16] ),
    .A1(\design_top.core0.REG1[9][16] ),
    .A2(\design_top.core0.REG1[10][16] ),
    .A3(\design_top.core0.REG1[11][16] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13932_ (.A0(\design_top.core0.REG1[12][16] ),
    .A1(\design_top.core0.REG1[13][16] ),
    .A2(\design_top.core0.REG1[14][16] ),
    .A3(\design_top.core0.REG1[15][16] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13933_ (.A0(_00466_),
    .A1(_00467_),
    .A2(_00468_),
    .A3(_00469_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13934_ (.A0(\design_top.core0.REG1[0][17] ),
    .A1(\design_top.core0.REG1[1][17] ),
    .A2(\design_top.core0.REG1[2][17] ),
    .A3(\design_top.core0.REG1[3][17] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13935_ (.A0(\design_top.core0.REG1[4][17] ),
    .A1(\design_top.core0.REG1[5][17] ),
    .A2(\design_top.core0.REG1[6][17] ),
    .A3(\design_top.core0.REG1[7][17] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13936_ (.A0(\design_top.core0.REG1[8][17] ),
    .A1(\design_top.core0.REG1[9][17] ),
    .A2(\design_top.core0.REG1[10][17] ),
    .A3(\design_top.core0.REG1[11][17] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13937_ (.A0(\design_top.core0.REG1[12][17] ),
    .A1(\design_top.core0.REG1[13][17] ),
    .A2(\design_top.core0.REG1[14][17] ),
    .A3(\design_top.core0.REG1[15][17] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13938_ (.A0(_00460_),
    .A1(_00461_),
    .A2(_00462_),
    .A3(_00463_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13939_ (.A0(\design_top.core0.REG1[0][18] ),
    .A1(\design_top.core0.REG1[1][18] ),
    .A2(\design_top.core0.REG1[2][18] ),
    .A3(\design_top.core0.REG1[3][18] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13940_ (.A0(\design_top.core0.REG1[4][18] ),
    .A1(\design_top.core0.REG1[5][18] ),
    .A2(\design_top.core0.REG1[6][18] ),
    .A3(\design_top.core0.REG1[7][18] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13941_ (.A0(\design_top.core0.REG1[8][18] ),
    .A1(\design_top.core0.REG1[9][18] ),
    .A2(\design_top.core0.REG1[10][18] ),
    .A3(\design_top.core0.REG1[11][18] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13942_ (.A0(\design_top.core0.REG1[12][18] ),
    .A1(\design_top.core0.REG1[13][18] ),
    .A2(\design_top.core0.REG1[14][18] ),
    .A3(\design_top.core0.REG1[15][18] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13943_ (.A0(_00454_),
    .A1(_00455_),
    .A2(_00456_),
    .A3(_00457_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13944_ (.A0(\design_top.core0.REG1[0][19] ),
    .A1(\design_top.core0.REG1[1][19] ),
    .A2(\design_top.core0.REG1[2][19] ),
    .A3(\design_top.core0.REG1[3][19] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13945_ (.A0(\design_top.core0.REG1[4][19] ),
    .A1(\design_top.core0.REG1[5][19] ),
    .A2(\design_top.core0.REG1[6][19] ),
    .A3(\design_top.core0.REG1[7][19] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13946_ (.A0(\design_top.core0.REG1[8][19] ),
    .A1(\design_top.core0.REG1[9][19] ),
    .A2(\design_top.core0.REG1[10][19] ),
    .A3(\design_top.core0.REG1[11][19] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13947_ (.A0(\design_top.core0.REG1[12][19] ),
    .A1(\design_top.core0.REG1[13][19] ),
    .A2(\design_top.core0.REG1[14][19] ),
    .A3(\design_top.core0.REG1[15][19] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13948_ (.A0(_00448_),
    .A1(_00449_),
    .A2(_00450_),
    .A3(_00451_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13949_ (.A0(\design_top.core0.REG1[0][20] ),
    .A1(\design_top.core0.REG1[1][20] ),
    .A2(\design_top.core0.REG1[2][20] ),
    .A3(\design_top.core0.REG1[3][20] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13950_ (.A0(\design_top.core0.REG1[4][20] ),
    .A1(\design_top.core0.REG1[5][20] ),
    .A2(\design_top.core0.REG1[6][20] ),
    .A3(\design_top.core0.REG1[7][20] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13951_ (.A0(\design_top.core0.REG1[8][20] ),
    .A1(\design_top.core0.REG1[9][20] ),
    .A2(\design_top.core0.REG1[10][20] ),
    .A3(\design_top.core0.REG1[11][20] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13952_ (.A0(\design_top.core0.REG1[12][20] ),
    .A1(\design_top.core0.REG1[13][20] ),
    .A2(\design_top.core0.REG1[14][20] ),
    .A3(\design_top.core0.REG1[15][20] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13953_ (.A0(_00442_),
    .A1(_00443_),
    .A2(_00444_),
    .A3(_00445_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13954_ (.A0(\design_top.core0.REG1[0][21] ),
    .A1(\design_top.core0.REG1[1][21] ),
    .A2(\design_top.core0.REG1[2][21] ),
    .A3(\design_top.core0.REG1[3][21] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13955_ (.A0(\design_top.core0.REG1[4][21] ),
    .A1(\design_top.core0.REG1[5][21] ),
    .A2(\design_top.core0.REG1[6][21] ),
    .A3(\design_top.core0.REG1[7][21] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13956_ (.A0(\design_top.core0.REG1[8][21] ),
    .A1(\design_top.core0.REG1[9][21] ),
    .A2(\design_top.core0.REG1[10][21] ),
    .A3(\design_top.core0.REG1[11][21] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13957_ (.A0(\design_top.core0.REG1[12][21] ),
    .A1(\design_top.core0.REG1[13][21] ),
    .A2(\design_top.core0.REG1[14][21] ),
    .A3(\design_top.core0.REG1[15][21] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13958_ (.A0(_00436_),
    .A1(_00437_),
    .A2(_00438_),
    .A3(_00439_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13959_ (.A0(\design_top.core0.REG1[0][22] ),
    .A1(\design_top.core0.REG1[1][22] ),
    .A2(\design_top.core0.REG1[2][22] ),
    .A3(\design_top.core0.REG1[3][22] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13960_ (.A0(\design_top.core0.REG1[4][22] ),
    .A1(\design_top.core0.REG1[5][22] ),
    .A2(\design_top.core0.REG1[6][22] ),
    .A3(\design_top.core0.REG1[7][22] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13961_ (.A0(\design_top.core0.REG1[8][22] ),
    .A1(\design_top.core0.REG1[9][22] ),
    .A2(\design_top.core0.REG1[10][22] ),
    .A3(\design_top.core0.REG1[11][22] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13962_ (.A0(\design_top.core0.REG1[12][22] ),
    .A1(\design_top.core0.REG1[13][22] ),
    .A2(\design_top.core0.REG1[14][22] ),
    .A3(\design_top.core0.REG1[15][22] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13963_ (.A0(_00430_),
    .A1(_00431_),
    .A2(_00432_),
    .A3(_00433_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13964_ (.A0(\design_top.core0.REG1[0][23] ),
    .A1(\design_top.core0.REG1[1][23] ),
    .A2(\design_top.core0.REG1[2][23] ),
    .A3(\design_top.core0.REG1[3][23] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13965_ (.A0(\design_top.core0.REG1[4][23] ),
    .A1(\design_top.core0.REG1[5][23] ),
    .A2(\design_top.core0.REG1[6][23] ),
    .A3(\design_top.core0.REG1[7][23] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13966_ (.A0(\design_top.core0.REG1[8][23] ),
    .A1(\design_top.core0.REG1[9][23] ),
    .A2(\design_top.core0.REG1[10][23] ),
    .A3(\design_top.core0.REG1[11][23] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13967_ (.A0(\design_top.core0.REG1[12][23] ),
    .A1(\design_top.core0.REG1[13][23] ),
    .A2(\design_top.core0.REG1[14][23] ),
    .A3(\design_top.core0.REG1[15][23] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13968_ (.A0(_00424_),
    .A1(_00425_),
    .A2(_00426_),
    .A3(_00427_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13969_ (.A0(\design_top.core0.REG1[0][24] ),
    .A1(\design_top.core0.REG1[1][24] ),
    .A2(\design_top.core0.REG1[2][24] ),
    .A3(\design_top.core0.REG1[3][24] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13970_ (.A0(\design_top.core0.REG1[4][24] ),
    .A1(\design_top.core0.REG1[5][24] ),
    .A2(\design_top.core0.REG1[6][24] ),
    .A3(\design_top.core0.REG1[7][24] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13971_ (.A0(\design_top.core0.REG1[8][24] ),
    .A1(\design_top.core0.REG1[9][24] ),
    .A2(\design_top.core0.REG1[10][24] ),
    .A3(\design_top.core0.REG1[11][24] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13972_ (.A0(\design_top.core0.REG1[12][24] ),
    .A1(\design_top.core0.REG1[13][24] ),
    .A2(\design_top.core0.REG1[14][24] ),
    .A3(\design_top.core0.REG1[15][24] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13973_ (.A0(_00418_),
    .A1(_00419_),
    .A2(_00420_),
    .A3(_00421_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13974_ (.A0(\design_top.core0.REG1[0][25] ),
    .A1(\design_top.core0.REG1[1][25] ),
    .A2(\design_top.core0.REG1[2][25] ),
    .A3(\design_top.core0.REG1[3][25] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13975_ (.A0(\design_top.core0.REG1[4][25] ),
    .A1(\design_top.core0.REG1[5][25] ),
    .A2(\design_top.core0.REG1[6][25] ),
    .A3(\design_top.core0.REG1[7][25] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13976_ (.A0(\design_top.core0.REG1[8][25] ),
    .A1(\design_top.core0.REG1[9][25] ),
    .A2(\design_top.core0.REG1[10][25] ),
    .A3(\design_top.core0.REG1[11][25] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13977_ (.A0(\design_top.core0.REG1[12][25] ),
    .A1(\design_top.core0.REG1[13][25] ),
    .A2(\design_top.core0.REG1[14][25] ),
    .A3(\design_top.core0.REG1[15][25] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13978_ (.A0(_00412_),
    .A1(_00413_),
    .A2(_00414_),
    .A3(_00415_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13979_ (.A0(\design_top.core0.REG1[0][26] ),
    .A1(\design_top.core0.REG1[1][26] ),
    .A2(\design_top.core0.REG1[2][26] ),
    .A3(\design_top.core0.REG1[3][26] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13980_ (.A0(\design_top.core0.REG1[4][26] ),
    .A1(\design_top.core0.REG1[5][26] ),
    .A2(\design_top.core0.REG1[6][26] ),
    .A3(\design_top.core0.REG1[7][26] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13981_ (.A0(\design_top.core0.REG1[8][26] ),
    .A1(\design_top.core0.REG1[9][26] ),
    .A2(\design_top.core0.REG1[10][26] ),
    .A3(\design_top.core0.REG1[11][26] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13982_ (.A0(\design_top.core0.REG1[12][26] ),
    .A1(\design_top.core0.REG1[13][26] ),
    .A2(\design_top.core0.REG1[14][26] ),
    .A3(\design_top.core0.REG1[15][26] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13983_ (.A0(_00406_),
    .A1(_00407_),
    .A2(_00408_),
    .A3(_00409_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13984_ (.A0(\design_top.core0.REG1[0][27] ),
    .A1(\design_top.core0.REG1[1][27] ),
    .A2(\design_top.core0.REG1[2][27] ),
    .A3(\design_top.core0.REG1[3][27] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13985_ (.A0(\design_top.core0.REG1[4][27] ),
    .A1(\design_top.core0.REG1[5][27] ),
    .A2(\design_top.core0.REG1[6][27] ),
    .A3(\design_top.core0.REG1[7][27] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13986_ (.A0(\design_top.core0.REG1[8][27] ),
    .A1(\design_top.core0.REG1[9][27] ),
    .A2(\design_top.core0.REG1[10][27] ),
    .A3(\design_top.core0.REG1[11][27] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13987_ (.A0(\design_top.core0.REG1[12][27] ),
    .A1(\design_top.core0.REG1[13][27] ),
    .A2(\design_top.core0.REG1[14][27] ),
    .A3(\design_top.core0.REG1[15][27] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13988_ (.A0(_00400_),
    .A1(_00401_),
    .A2(_00402_),
    .A3(_00403_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13989_ (.A0(\design_top.core0.REG1[0][28] ),
    .A1(\design_top.core0.REG1[1][28] ),
    .A2(\design_top.core0.REG1[2][28] ),
    .A3(\design_top.core0.REG1[3][28] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13990_ (.A0(\design_top.core0.REG1[4][28] ),
    .A1(\design_top.core0.REG1[5][28] ),
    .A2(\design_top.core0.REG1[6][28] ),
    .A3(\design_top.core0.REG1[7][28] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13991_ (.A0(\design_top.core0.REG1[8][28] ),
    .A1(\design_top.core0.REG1[9][28] ),
    .A2(\design_top.core0.REG1[10][28] ),
    .A3(\design_top.core0.REG1[11][28] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13992_ (.A0(\design_top.core0.REG1[12][28] ),
    .A1(\design_top.core0.REG1[13][28] ),
    .A2(\design_top.core0.REG1[14][28] ),
    .A3(\design_top.core0.REG1[15][28] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13993_ (.A0(_00394_),
    .A1(_00395_),
    .A2(_00396_),
    .A3(_00397_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13994_ (.A0(\design_top.core0.REG1[0][29] ),
    .A1(\design_top.core0.REG1[1][29] ),
    .A2(\design_top.core0.REG1[2][29] ),
    .A3(\design_top.core0.REG1[3][29] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13995_ (.A0(\design_top.core0.REG1[4][29] ),
    .A1(\design_top.core0.REG1[5][29] ),
    .A2(\design_top.core0.REG1[6][29] ),
    .A3(\design_top.core0.REG1[7][29] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13996_ (.A0(\design_top.core0.REG1[8][29] ),
    .A1(\design_top.core0.REG1[9][29] ),
    .A2(\design_top.core0.REG1[10][29] ),
    .A3(\design_top.core0.REG1[11][29] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13997_ (.A0(\design_top.core0.REG1[12][29] ),
    .A1(\design_top.core0.REG1[13][29] ),
    .A2(\design_top.core0.REG1[14][29] ),
    .A3(\design_top.core0.REG1[15][29] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13998_ (.A0(_00388_),
    .A1(_00389_),
    .A2(_00390_),
    .A3(_00391_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _13999_ (.A0(\design_top.core0.REG1[0][30] ),
    .A1(\design_top.core0.REG1[1][30] ),
    .A2(\design_top.core0.REG1[2][30] ),
    .A3(\design_top.core0.REG1[3][30] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14000_ (.A0(\design_top.core0.REG1[4][30] ),
    .A1(\design_top.core0.REG1[5][30] ),
    .A2(\design_top.core0.REG1[6][30] ),
    .A3(\design_top.core0.REG1[7][30] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14001_ (.A0(\design_top.core0.REG1[8][30] ),
    .A1(\design_top.core0.REG1[9][30] ),
    .A2(\design_top.core0.REG1[10][30] ),
    .A3(\design_top.core0.REG1[11][30] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14002_ (.A0(\design_top.core0.REG1[12][30] ),
    .A1(\design_top.core0.REG1[13][30] ),
    .A2(\design_top.core0.REG1[14][30] ),
    .A3(\design_top.core0.REG1[15][30] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14003_ (.A0(_00382_),
    .A1(_00383_),
    .A2(_00384_),
    .A3(_00385_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14004_ (.A0(_00361_),
    .A1(_00362_),
    .A2(_00363_),
    .A3(_00364_),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14005_ (.A0(_00366_),
    .A1(_00367_),
    .A2(_00368_),
    .A3(_00369_),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14006_ (.A0(_00371_),
    .A1(_00372_),
    .A2(_00373_),
    .A3(_00374_),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14007_ (.A0(_00376_),
    .A1(_00377_),
    .A2(_00378_),
    .A3(_00379_),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14008_ (.A0(_00365_),
    .A1(_00370_),
    .A2(_00375_),
    .A3(_00380_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14009_ (.A0(\design_top.core0.REG1[0][5] ),
    .A1(\design_top.core0.REG1[1][5] ),
    .A2(\design_top.core0.REG1[2][5] ),
    .A3(\design_top.core0.REG1[3][5] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14010_ (.A0(\design_top.core0.REG1[4][5] ),
    .A1(\design_top.core0.REG1[5][5] ),
    .A2(\design_top.core0.REG1[6][5] ),
    .A3(\design_top.core0.REG1[7][5] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14011_ (.A0(\design_top.core0.REG1[8][5] ),
    .A1(\design_top.core0.REG1[9][5] ),
    .A2(\design_top.core0.REG1[10][5] ),
    .A3(\design_top.core0.REG1[11][5] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14012_ (.A0(\design_top.core0.REG1[12][5] ),
    .A1(\design_top.core0.REG1[13][5] ),
    .A2(\design_top.core0.REG1[14][5] ),
    .A3(\design_top.core0.REG1[15][5] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14013_ (.A0(_00355_),
    .A1(_00356_),
    .A2(_00357_),
    .A3(_00358_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14014_ (.A0(\design_top.core0.REG1[0][4] ),
    .A1(\design_top.core0.REG1[1][4] ),
    .A2(\design_top.core0.REG1[2][4] ),
    .A3(\design_top.core0.REG1[3][4] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14015_ (.A0(\design_top.core0.REG1[4][4] ),
    .A1(\design_top.core0.REG1[5][4] ),
    .A2(\design_top.core0.REG1[6][4] ),
    .A3(\design_top.core0.REG1[7][4] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14016_ (.A0(\design_top.core0.REG1[8][4] ),
    .A1(\design_top.core0.REG1[9][4] ),
    .A2(\design_top.core0.REG1[10][4] ),
    .A3(\design_top.core0.REG1[11][4] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14017_ (.A0(\design_top.core0.REG1[12][4] ),
    .A1(\design_top.core0.REG1[13][4] ),
    .A2(\design_top.core0.REG1[14][4] ),
    .A3(\design_top.core0.REG1[15][4] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14018_ (.A0(_00348_),
    .A1(_00349_),
    .A2(_00350_),
    .A3(_00351_),
    .S0(_00303_),
    .S1(_00304_),
    .X(_00352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14019_ (.A0(\design_top.core0.REG1[8][3] ),
    .A1(\design_top.core0.REG1[9][3] ),
    .A2(\design_top.core0.REG1[10][3] ),
    .A3(\design_top.core0.REG1[11][3] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14020_ (.A0(\design_top.core0.REG1[12][3] ),
    .A1(\design_top.core0.REG1[13][3] ),
    .A2(\design_top.core0.REG1[14][3] ),
    .A3(\design_top.core0.REG1[15][3] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14021_ (.A0(\design_top.core0.REG1[0][3] ),
    .A1(\design_top.core0.REG1[1][3] ),
    .A2(\design_top.core0.REG1[2][3] ),
    .A3(\design_top.core0.REG1[3][3] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14022_ (.A0(\design_top.core0.REG1[4][3] ),
    .A1(\design_top.core0.REG1[5][3] ),
    .A2(\design_top.core0.REG1[6][3] ),
    .A3(\design_top.core0.REG1[7][3] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14023_ (.A0(\design_top.core0.REG1[8][0] ),
    .A1(\design_top.core0.REG1[9][0] ),
    .A2(\design_top.core0.REG1[10][0] ),
    .A3(\design_top.core0.REG1[11][0] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14024_ (.A0(\design_top.core0.REG1[12][0] ),
    .A1(\design_top.core0.REG1[13][0] ),
    .A2(\design_top.core0.REG1[14][0] ),
    .A3(\design_top.core0.REG1[15][0] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14025_ (.A0(\design_top.core0.REG1[0][0] ),
    .A1(\design_top.core0.REG1[1][0] ),
    .A2(\design_top.core0.REG1[2][0] ),
    .A3(\design_top.core0.REG1[3][0] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14026_ (.A0(\design_top.core0.REG1[4][0] ),
    .A1(\design_top.core0.REG1[5][0] ),
    .A2(\design_top.core0.REG1[6][0] ),
    .A3(\design_top.core0.REG1[7][0] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14027_ (.A0(\design_top.core0.REG1[8][1] ),
    .A1(\design_top.core0.REG1[9][1] ),
    .A2(\design_top.core0.REG1[10][1] ),
    .A3(\design_top.core0.REG1[11][1] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14028_ (.A0(\design_top.core0.REG1[12][1] ),
    .A1(\design_top.core0.REG1[13][1] ),
    .A2(\design_top.core0.REG1[14][1] ),
    .A3(\design_top.core0.REG1[15][1] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14029_ (.A0(\design_top.core0.REG1[0][1] ),
    .A1(\design_top.core0.REG1[1][1] ),
    .A2(\design_top.core0.REG1[2][1] ),
    .A3(\design_top.core0.REG1[3][1] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14030_ (.A0(\design_top.core0.REG1[4][1] ),
    .A1(\design_top.core0.REG1[5][1] ),
    .A2(\design_top.core0.REG1[6][1] ),
    .A3(\design_top.core0.REG1[7][1] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14031_ (.A0(\design_top.core0.REG1[8][2] ),
    .A1(\design_top.core0.REG1[9][2] ),
    .A2(\design_top.core0.REG1[10][2] ),
    .A3(\design_top.core0.REG1[11][2] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14032_ (.A0(\design_top.core0.REG1[12][2] ),
    .A1(\design_top.core0.REG1[13][2] ),
    .A2(\design_top.core0.REG1[14][2] ),
    .A3(\design_top.core0.REG1[15][2] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14033_ (.A0(\design_top.core0.REG1[0][2] ),
    .A1(\design_top.core0.REG1[1][2] ),
    .A2(\design_top.core0.REG1[2][2] ),
    .A3(\design_top.core0.REG1[3][2] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14034_ (.A0(\design_top.core0.REG1[4][2] ),
    .A1(\design_top.core0.REG1[5][2] ),
    .A2(\design_top.core0.REG1[6][2] ),
    .A3(\design_top.core0.REG1[7][2] ),
    .S0(_00301_),
    .S1(_00302_),
    .X(_00312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14035_ (.A0(\design_top.MEM[15][31] ),
    .A1(\design_top.MEM[14][31] ),
    .A2(\design_top.MEM[13][31] ),
    .A3(\design_top.MEM[12][31] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14036_ (.A0(\design_top.MEM[11][31] ),
    .A1(\design_top.MEM[10][31] ),
    .A2(\design_top.MEM[9][31] ),
    .A3(\design_top.MEM[8][31] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14037_ (.A0(\design_top.MEM[7][31] ),
    .A1(\design_top.MEM[6][31] ),
    .A2(\design_top.MEM[5][31] ),
    .A3(\design_top.MEM[4][31] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14038_ (.A0(\design_top.MEM[3][31] ),
    .A1(\design_top.MEM[2][31] ),
    .A2(\design_top.MEM[1][31] ),
    .A3(\design_top.MEM[0][31] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14039_ (.A0(_01239_),
    .A1(_01238_),
    .A2(_01237_),
    .A3(_01236_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14040_ (.A0(\design_top.MEM[15][30] ),
    .A1(\design_top.MEM[14][30] ),
    .A2(\design_top.MEM[13][30] ),
    .A3(\design_top.MEM[12][30] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14041_ (.A0(\design_top.MEM[11][30] ),
    .A1(\design_top.MEM[10][30] ),
    .A2(\design_top.MEM[9][30] ),
    .A3(\design_top.MEM[8][30] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14042_ (.A0(\design_top.MEM[7][30] ),
    .A1(\design_top.MEM[6][30] ),
    .A2(\design_top.MEM[5][30] ),
    .A3(\design_top.MEM[4][30] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14043_ (.A0(\design_top.MEM[3][30] ),
    .A1(\design_top.MEM[2][30] ),
    .A2(\design_top.MEM[1][30] ),
    .A3(\design_top.MEM[0][30] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14044_ (.A0(_01235_),
    .A1(_01234_),
    .A2(_01233_),
    .A3(_01232_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14045_ (.A0(\design_top.MEM[15][29] ),
    .A1(\design_top.MEM[14][29] ),
    .A2(\design_top.MEM[13][29] ),
    .A3(\design_top.MEM[12][29] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14046_ (.A0(\design_top.MEM[11][29] ),
    .A1(\design_top.MEM[10][29] ),
    .A2(\design_top.MEM[9][29] ),
    .A3(\design_top.MEM[8][29] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14047_ (.A0(\design_top.MEM[7][29] ),
    .A1(\design_top.MEM[6][29] ),
    .A2(\design_top.MEM[5][29] ),
    .A3(\design_top.MEM[4][29] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14048_ (.A0(\design_top.MEM[3][29] ),
    .A1(\design_top.MEM[2][29] ),
    .A2(\design_top.MEM[1][29] ),
    .A3(\design_top.MEM[0][29] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14049_ (.A0(_01231_),
    .A1(_01230_),
    .A2(_01229_),
    .A3(_01228_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14050_ (.A0(\design_top.MEM[15][28] ),
    .A1(\design_top.MEM[14][28] ),
    .A2(\design_top.MEM[13][28] ),
    .A3(\design_top.MEM[12][28] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14051_ (.A0(\design_top.MEM[11][28] ),
    .A1(\design_top.MEM[10][28] ),
    .A2(\design_top.MEM[9][28] ),
    .A3(\design_top.MEM[8][28] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14052_ (.A0(\design_top.MEM[7][28] ),
    .A1(\design_top.MEM[6][28] ),
    .A2(\design_top.MEM[5][28] ),
    .A3(\design_top.MEM[4][28] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14053_ (.A0(\design_top.MEM[3][28] ),
    .A1(\design_top.MEM[2][28] ),
    .A2(\design_top.MEM[1][28] ),
    .A3(\design_top.MEM[0][28] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14054_ (.A0(_01227_),
    .A1(_01226_),
    .A2(_01225_),
    .A3(_01224_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14055_ (.A0(\design_top.MEM[15][27] ),
    .A1(\design_top.MEM[14][27] ),
    .A2(\design_top.MEM[13][27] ),
    .A3(\design_top.MEM[12][27] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14056_ (.A0(\design_top.MEM[11][27] ),
    .A1(\design_top.MEM[10][27] ),
    .A2(\design_top.MEM[9][27] ),
    .A3(\design_top.MEM[8][27] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14057_ (.A0(\design_top.MEM[7][27] ),
    .A1(\design_top.MEM[6][27] ),
    .A2(\design_top.MEM[5][27] ),
    .A3(\design_top.MEM[4][27] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14058_ (.A0(\design_top.MEM[3][27] ),
    .A1(\design_top.MEM[2][27] ),
    .A2(\design_top.MEM[1][27] ),
    .A3(\design_top.MEM[0][27] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14059_ (.A0(_01223_),
    .A1(_01222_),
    .A2(_01221_),
    .A3(_01220_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14060_ (.A0(\design_top.MEM[15][26] ),
    .A1(\design_top.MEM[14][26] ),
    .A2(\design_top.MEM[13][26] ),
    .A3(\design_top.MEM[12][26] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14061_ (.A0(\design_top.MEM[11][26] ),
    .A1(\design_top.MEM[10][26] ),
    .A2(\design_top.MEM[9][26] ),
    .A3(\design_top.MEM[8][26] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14062_ (.A0(\design_top.MEM[7][26] ),
    .A1(\design_top.MEM[6][26] ),
    .A2(\design_top.MEM[5][26] ),
    .A3(\design_top.MEM[4][26] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14063_ (.A0(\design_top.MEM[3][26] ),
    .A1(\design_top.MEM[2][26] ),
    .A2(\design_top.MEM[1][26] ),
    .A3(\design_top.MEM[0][26] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14064_ (.A0(_01219_),
    .A1(_01218_),
    .A2(_01217_),
    .A3(_01216_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14065_ (.A0(\design_top.MEM[15][25] ),
    .A1(\design_top.MEM[14][25] ),
    .A2(\design_top.MEM[13][25] ),
    .A3(\design_top.MEM[12][25] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14066_ (.A0(\design_top.MEM[11][25] ),
    .A1(\design_top.MEM[10][25] ),
    .A2(\design_top.MEM[9][25] ),
    .A3(\design_top.MEM[8][25] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14067_ (.A0(\design_top.MEM[7][25] ),
    .A1(\design_top.MEM[6][25] ),
    .A2(\design_top.MEM[5][25] ),
    .A3(\design_top.MEM[4][25] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14068_ (.A0(\design_top.MEM[3][25] ),
    .A1(\design_top.MEM[2][25] ),
    .A2(\design_top.MEM[1][25] ),
    .A3(\design_top.MEM[0][25] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14069_ (.A0(_01215_),
    .A1(_01214_),
    .A2(_01213_),
    .A3(_01212_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14070_ (.A0(\design_top.MEM[15][24] ),
    .A1(\design_top.MEM[14][24] ),
    .A2(\design_top.MEM[13][24] ),
    .A3(\design_top.MEM[12][24] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14071_ (.A0(\design_top.MEM[11][24] ),
    .A1(\design_top.MEM[10][24] ),
    .A2(\design_top.MEM[9][24] ),
    .A3(\design_top.MEM[8][24] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14072_ (.A0(\design_top.MEM[7][24] ),
    .A1(\design_top.MEM[6][24] ),
    .A2(\design_top.MEM[5][24] ),
    .A3(\design_top.MEM[4][24] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14073_ (.A0(\design_top.MEM[3][24] ),
    .A1(\design_top.MEM[2][24] ),
    .A2(\design_top.MEM[1][24] ),
    .A3(\design_top.MEM[0][24] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14074_ (.A0(_01211_),
    .A1(_01210_),
    .A2(_01209_),
    .A3(_01208_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14075_ (.A0(\design_top.MEM[15][23] ),
    .A1(\design_top.MEM[14][23] ),
    .A2(\design_top.MEM[13][23] ),
    .A3(\design_top.MEM[12][23] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14076_ (.A0(\design_top.MEM[11][23] ),
    .A1(\design_top.MEM[10][23] ),
    .A2(\design_top.MEM[9][23] ),
    .A3(\design_top.MEM[8][23] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14077_ (.A0(\design_top.MEM[7][23] ),
    .A1(\design_top.MEM[6][23] ),
    .A2(\design_top.MEM[5][23] ),
    .A3(\design_top.MEM[4][23] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14078_ (.A0(\design_top.MEM[3][23] ),
    .A1(\design_top.MEM[2][23] ),
    .A2(\design_top.MEM[1][23] ),
    .A3(\design_top.MEM[0][23] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14079_ (.A0(_01207_),
    .A1(_01206_),
    .A2(_01205_),
    .A3(_01204_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14080_ (.A0(\design_top.MEM[15][22] ),
    .A1(\design_top.MEM[14][22] ),
    .A2(\design_top.MEM[13][22] ),
    .A3(\design_top.MEM[12][22] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14081_ (.A0(\design_top.MEM[11][22] ),
    .A1(\design_top.MEM[10][22] ),
    .A2(\design_top.MEM[9][22] ),
    .A3(\design_top.MEM[8][22] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14082_ (.A0(\design_top.MEM[7][22] ),
    .A1(\design_top.MEM[6][22] ),
    .A2(\design_top.MEM[5][22] ),
    .A3(\design_top.MEM[4][22] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14083_ (.A0(\design_top.MEM[3][22] ),
    .A1(\design_top.MEM[2][22] ),
    .A2(\design_top.MEM[1][22] ),
    .A3(\design_top.MEM[0][22] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14084_ (.A0(_01203_),
    .A1(_01202_),
    .A2(_01201_),
    .A3(_01200_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14085_ (.A0(\design_top.MEM[15][21] ),
    .A1(\design_top.MEM[14][21] ),
    .A2(\design_top.MEM[13][21] ),
    .A3(\design_top.MEM[12][21] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14086_ (.A0(\design_top.MEM[11][21] ),
    .A1(\design_top.MEM[10][21] ),
    .A2(\design_top.MEM[9][21] ),
    .A3(\design_top.MEM[8][21] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14087_ (.A0(\design_top.MEM[7][21] ),
    .A1(\design_top.MEM[6][21] ),
    .A2(\design_top.MEM[5][21] ),
    .A3(\design_top.MEM[4][21] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14088_ (.A0(\design_top.MEM[3][21] ),
    .A1(\design_top.MEM[2][21] ),
    .A2(\design_top.MEM[1][21] ),
    .A3(\design_top.MEM[0][21] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14089_ (.A0(_01199_),
    .A1(_01198_),
    .A2(_01197_),
    .A3(_01196_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14090_ (.A0(\design_top.MEM[15][20] ),
    .A1(\design_top.MEM[14][20] ),
    .A2(\design_top.MEM[13][20] ),
    .A3(\design_top.MEM[12][20] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14091_ (.A0(\design_top.MEM[11][20] ),
    .A1(\design_top.MEM[10][20] ),
    .A2(\design_top.MEM[9][20] ),
    .A3(\design_top.MEM[8][20] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14092_ (.A0(\design_top.MEM[7][20] ),
    .A1(\design_top.MEM[6][20] ),
    .A2(\design_top.MEM[5][20] ),
    .A3(\design_top.MEM[4][20] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14093_ (.A0(\design_top.MEM[3][20] ),
    .A1(\design_top.MEM[2][20] ),
    .A2(\design_top.MEM[1][20] ),
    .A3(\design_top.MEM[0][20] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14094_ (.A0(_01195_),
    .A1(_01194_),
    .A2(_01193_),
    .A3(_01192_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14095_ (.A0(\design_top.MEM[15][19] ),
    .A1(\design_top.MEM[14][19] ),
    .A2(\design_top.MEM[13][19] ),
    .A3(\design_top.MEM[12][19] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14096_ (.A0(\design_top.MEM[11][19] ),
    .A1(\design_top.MEM[10][19] ),
    .A2(\design_top.MEM[9][19] ),
    .A3(\design_top.MEM[8][19] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14097_ (.A0(\design_top.MEM[7][19] ),
    .A1(\design_top.MEM[6][19] ),
    .A2(\design_top.MEM[5][19] ),
    .A3(\design_top.MEM[4][19] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14098_ (.A0(\design_top.MEM[3][19] ),
    .A1(\design_top.MEM[2][19] ),
    .A2(\design_top.MEM[1][19] ),
    .A3(\design_top.MEM[0][19] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14099_ (.A0(_01191_),
    .A1(_01190_),
    .A2(_01189_),
    .A3(_01188_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14100_ (.A0(\design_top.MEM[15][18] ),
    .A1(\design_top.MEM[14][18] ),
    .A2(\design_top.MEM[13][18] ),
    .A3(\design_top.MEM[12][18] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14101_ (.A0(\design_top.MEM[11][18] ),
    .A1(\design_top.MEM[10][18] ),
    .A2(\design_top.MEM[9][18] ),
    .A3(\design_top.MEM[8][18] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14102_ (.A0(\design_top.MEM[7][18] ),
    .A1(\design_top.MEM[6][18] ),
    .A2(\design_top.MEM[5][18] ),
    .A3(\design_top.MEM[4][18] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14103_ (.A0(\design_top.MEM[3][18] ),
    .A1(\design_top.MEM[2][18] ),
    .A2(\design_top.MEM[1][18] ),
    .A3(\design_top.MEM[0][18] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14104_ (.A0(_01187_),
    .A1(_01186_),
    .A2(_01185_),
    .A3(_01184_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14105_ (.A0(\design_top.MEM[15][17] ),
    .A1(\design_top.MEM[14][17] ),
    .A2(\design_top.MEM[13][17] ),
    .A3(\design_top.MEM[12][17] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14106_ (.A0(\design_top.MEM[11][17] ),
    .A1(\design_top.MEM[10][17] ),
    .A2(\design_top.MEM[9][17] ),
    .A3(\design_top.MEM[8][17] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14107_ (.A0(\design_top.MEM[7][17] ),
    .A1(\design_top.MEM[6][17] ),
    .A2(\design_top.MEM[5][17] ),
    .A3(\design_top.MEM[4][17] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14108_ (.A0(\design_top.MEM[3][17] ),
    .A1(\design_top.MEM[2][17] ),
    .A2(\design_top.MEM[1][17] ),
    .A3(\design_top.MEM[0][17] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14109_ (.A0(_01183_),
    .A1(_01182_),
    .A2(_01181_),
    .A3(_01180_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14110_ (.A0(\design_top.MEM[15][16] ),
    .A1(\design_top.MEM[14][16] ),
    .A2(\design_top.MEM[13][16] ),
    .A3(\design_top.MEM[12][16] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14111_ (.A0(\design_top.MEM[11][16] ),
    .A1(\design_top.MEM[10][16] ),
    .A2(\design_top.MEM[9][16] ),
    .A3(\design_top.MEM[8][16] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14112_ (.A0(\design_top.MEM[7][16] ),
    .A1(\design_top.MEM[6][16] ),
    .A2(\design_top.MEM[5][16] ),
    .A3(\design_top.MEM[4][16] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14113_ (.A0(\design_top.MEM[3][16] ),
    .A1(\design_top.MEM[2][16] ),
    .A2(\design_top.MEM[1][16] ),
    .A3(\design_top.MEM[0][16] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14114_ (.A0(_01179_),
    .A1(_01178_),
    .A2(_01177_),
    .A3(_01176_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14115_ (.A0(\design_top.MEM[15][15] ),
    .A1(\design_top.MEM[14][15] ),
    .A2(\design_top.MEM[13][15] ),
    .A3(\design_top.MEM[12][15] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14116_ (.A0(\design_top.MEM[11][15] ),
    .A1(\design_top.MEM[10][15] ),
    .A2(\design_top.MEM[9][15] ),
    .A3(\design_top.MEM[8][15] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14117_ (.A0(\design_top.MEM[7][15] ),
    .A1(\design_top.MEM[6][15] ),
    .A2(\design_top.MEM[5][15] ),
    .A3(\design_top.MEM[4][15] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14118_ (.A0(\design_top.MEM[3][15] ),
    .A1(\design_top.MEM[2][15] ),
    .A2(\design_top.MEM[1][15] ),
    .A3(\design_top.MEM[0][15] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14119_ (.A0(_01175_),
    .A1(_01174_),
    .A2(_01173_),
    .A3(_01172_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14120_ (.A0(\design_top.MEM[15][14] ),
    .A1(\design_top.MEM[14][14] ),
    .A2(\design_top.MEM[13][14] ),
    .A3(\design_top.MEM[12][14] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14121_ (.A0(\design_top.MEM[11][14] ),
    .A1(\design_top.MEM[10][14] ),
    .A2(\design_top.MEM[9][14] ),
    .A3(\design_top.MEM[8][14] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14122_ (.A0(\design_top.MEM[7][14] ),
    .A1(\design_top.MEM[6][14] ),
    .A2(\design_top.MEM[5][14] ),
    .A3(\design_top.MEM[4][14] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14123_ (.A0(\design_top.MEM[3][14] ),
    .A1(\design_top.MEM[2][14] ),
    .A2(\design_top.MEM[1][14] ),
    .A3(\design_top.MEM[0][14] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14124_ (.A0(_01171_),
    .A1(_01170_),
    .A2(_01169_),
    .A3(_01168_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14125_ (.A0(\design_top.MEM[15][13] ),
    .A1(\design_top.MEM[14][13] ),
    .A2(\design_top.MEM[13][13] ),
    .A3(\design_top.MEM[12][13] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14126_ (.A0(\design_top.MEM[11][13] ),
    .A1(\design_top.MEM[10][13] ),
    .A2(\design_top.MEM[9][13] ),
    .A3(\design_top.MEM[8][13] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14127_ (.A0(\design_top.MEM[7][13] ),
    .A1(\design_top.MEM[6][13] ),
    .A2(\design_top.MEM[5][13] ),
    .A3(\design_top.MEM[4][13] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14128_ (.A0(\design_top.MEM[3][13] ),
    .A1(\design_top.MEM[2][13] ),
    .A2(\design_top.MEM[1][13] ),
    .A3(\design_top.MEM[0][13] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14129_ (.A0(_01167_),
    .A1(_01166_),
    .A2(_01165_),
    .A3(_01164_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14130_ (.A0(\design_top.MEM[15][12] ),
    .A1(\design_top.MEM[14][12] ),
    .A2(\design_top.MEM[13][12] ),
    .A3(\design_top.MEM[12][12] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14131_ (.A0(\design_top.MEM[11][12] ),
    .A1(\design_top.MEM[10][12] ),
    .A2(\design_top.MEM[9][12] ),
    .A3(\design_top.MEM[8][12] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14132_ (.A0(\design_top.MEM[7][12] ),
    .A1(\design_top.MEM[6][12] ),
    .A2(\design_top.MEM[5][12] ),
    .A3(\design_top.MEM[4][12] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14133_ (.A0(\design_top.MEM[3][12] ),
    .A1(\design_top.MEM[2][12] ),
    .A2(\design_top.MEM[1][12] ),
    .A3(\design_top.MEM[0][12] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14134_ (.A0(_01163_),
    .A1(_01162_),
    .A2(_01161_),
    .A3(_01160_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14135_ (.A0(\design_top.MEM[15][11] ),
    .A1(\design_top.MEM[14][11] ),
    .A2(\design_top.MEM[13][11] ),
    .A3(\design_top.MEM[12][11] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14136_ (.A0(\design_top.MEM[11][11] ),
    .A1(\design_top.MEM[10][11] ),
    .A2(\design_top.MEM[9][11] ),
    .A3(\design_top.MEM[8][11] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14137_ (.A0(\design_top.MEM[7][11] ),
    .A1(\design_top.MEM[6][11] ),
    .A2(\design_top.MEM[5][11] ),
    .A3(\design_top.MEM[4][11] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14138_ (.A0(\design_top.MEM[3][11] ),
    .A1(\design_top.MEM[2][11] ),
    .A2(\design_top.MEM[1][11] ),
    .A3(\design_top.MEM[0][11] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14139_ (.A0(_01159_),
    .A1(_01158_),
    .A2(_01157_),
    .A3(_01156_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14140_ (.A0(\design_top.MEM[15][10] ),
    .A1(\design_top.MEM[14][10] ),
    .A2(\design_top.MEM[13][10] ),
    .A3(\design_top.MEM[12][10] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14141_ (.A0(\design_top.MEM[11][10] ),
    .A1(\design_top.MEM[10][10] ),
    .A2(\design_top.MEM[9][10] ),
    .A3(\design_top.MEM[8][10] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14142_ (.A0(\design_top.MEM[7][10] ),
    .A1(\design_top.MEM[6][10] ),
    .A2(\design_top.MEM[5][10] ),
    .A3(\design_top.MEM[4][10] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14143_ (.A0(\design_top.MEM[3][10] ),
    .A1(\design_top.MEM[2][10] ),
    .A2(\design_top.MEM[1][10] ),
    .A3(\design_top.MEM[0][10] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14144_ (.A0(_01155_),
    .A1(_01154_),
    .A2(_01153_),
    .A3(_01152_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14145_ (.A0(\design_top.MEM[15][9] ),
    .A1(\design_top.MEM[14][9] ),
    .A2(\design_top.MEM[13][9] ),
    .A3(\design_top.MEM[12][9] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14146_ (.A0(\design_top.MEM[11][9] ),
    .A1(\design_top.MEM[10][9] ),
    .A2(\design_top.MEM[9][9] ),
    .A3(\design_top.MEM[8][9] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14147_ (.A0(\design_top.MEM[7][9] ),
    .A1(\design_top.MEM[6][9] ),
    .A2(\design_top.MEM[5][9] ),
    .A3(\design_top.MEM[4][9] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14148_ (.A0(\design_top.MEM[3][9] ),
    .A1(\design_top.MEM[2][9] ),
    .A2(\design_top.MEM[1][9] ),
    .A3(\design_top.MEM[0][9] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14149_ (.A0(_01151_),
    .A1(_01150_),
    .A2(_01149_),
    .A3(_01148_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14150_ (.A0(\design_top.MEM[15][8] ),
    .A1(\design_top.MEM[14][8] ),
    .A2(\design_top.MEM[13][8] ),
    .A3(\design_top.MEM[12][8] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14151_ (.A0(\design_top.MEM[11][8] ),
    .A1(\design_top.MEM[10][8] ),
    .A2(\design_top.MEM[9][8] ),
    .A3(\design_top.MEM[8][8] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14152_ (.A0(\design_top.MEM[7][8] ),
    .A1(\design_top.MEM[6][8] ),
    .A2(\design_top.MEM[5][8] ),
    .A3(\design_top.MEM[4][8] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14153_ (.A0(\design_top.MEM[3][8] ),
    .A1(\design_top.MEM[2][8] ),
    .A2(\design_top.MEM[1][8] ),
    .A3(\design_top.MEM[0][8] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14154_ (.A0(_01147_),
    .A1(_01146_),
    .A2(_01145_),
    .A3(_01144_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14155_ (.A0(\design_top.MEM[15][7] ),
    .A1(\design_top.MEM[14][7] ),
    .A2(\design_top.MEM[13][7] ),
    .A3(\design_top.MEM[12][7] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14156_ (.A0(\design_top.MEM[11][7] ),
    .A1(\design_top.MEM[10][7] ),
    .A2(\design_top.MEM[9][7] ),
    .A3(\design_top.MEM[8][7] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14157_ (.A0(\design_top.MEM[7][7] ),
    .A1(\design_top.MEM[6][7] ),
    .A2(\design_top.MEM[5][7] ),
    .A3(\design_top.MEM[4][7] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14158_ (.A0(\design_top.MEM[3][7] ),
    .A1(\design_top.MEM[2][7] ),
    .A2(\design_top.MEM[1][7] ),
    .A3(\design_top.MEM[0][7] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14159_ (.A0(_01143_),
    .A1(_01142_),
    .A2(_01141_),
    .A3(_01140_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14160_ (.A0(\design_top.MEM[15][6] ),
    .A1(\design_top.MEM[14][6] ),
    .A2(\design_top.MEM[13][6] ),
    .A3(\design_top.MEM[12][6] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14161_ (.A0(\design_top.MEM[11][6] ),
    .A1(\design_top.MEM[10][6] ),
    .A2(\design_top.MEM[9][6] ),
    .A3(\design_top.MEM[8][6] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14162_ (.A0(\design_top.MEM[7][6] ),
    .A1(\design_top.MEM[6][6] ),
    .A2(\design_top.MEM[5][6] ),
    .A3(\design_top.MEM[4][6] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14163_ (.A0(\design_top.MEM[3][6] ),
    .A1(\design_top.MEM[2][6] ),
    .A2(\design_top.MEM[1][6] ),
    .A3(\design_top.MEM[0][6] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14164_ (.A0(_01139_),
    .A1(_01138_),
    .A2(_01137_),
    .A3(_01136_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14165_ (.A0(\design_top.MEM[15][5] ),
    .A1(\design_top.MEM[14][5] ),
    .A2(\design_top.MEM[13][5] ),
    .A3(\design_top.MEM[12][5] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14166_ (.A0(\design_top.MEM[11][5] ),
    .A1(\design_top.MEM[10][5] ),
    .A2(\design_top.MEM[9][5] ),
    .A3(\design_top.MEM[8][5] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14167_ (.A0(\design_top.MEM[7][5] ),
    .A1(\design_top.MEM[6][5] ),
    .A2(\design_top.MEM[5][5] ),
    .A3(\design_top.MEM[4][5] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14168_ (.A0(\design_top.MEM[3][5] ),
    .A1(\design_top.MEM[2][5] ),
    .A2(\design_top.MEM[1][5] ),
    .A3(\design_top.MEM[0][5] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14169_ (.A0(_01135_),
    .A1(_01134_),
    .A2(_01133_),
    .A3(_01132_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14170_ (.A0(\design_top.MEM[15][4] ),
    .A1(\design_top.MEM[14][4] ),
    .A2(\design_top.MEM[13][4] ),
    .A3(\design_top.MEM[12][4] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14171_ (.A0(\design_top.MEM[11][4] ),
    .A1(\design_top.MEM[10][4] ),
    .A2(\design_top.MEM[9][4] ),
    .A3(\design_top.MEM[8][4] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14172_ (.A0(\design_top.MEM[7][4] ),
    .A1(\design_top.MEM[6][4] ),
    .A2(\design_top.MEM[5][4] ),
    .A3(\design_top.MEM[4][4] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14173_ (.A0(\design_top.MEM[3][4] ),
    .A1(\design_top.MEM[2][4] ),
    .A2(\design_top.MEM[1][4] ),
    .A3(\design_top.MEM[0][4] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14174_ (.A0(_01131_),
    .A1(_01130_),
    .A2(_01129_),
    .A3(_01128_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14175_ (.A0(\design_top.MEM[15][3] ),
    .A1(\design_top.MEM[14][3] ),
    .A2(\design_top.MEM[13][3] ),
    .A3(\design_top.MEM[12][3] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14176_ (.A0(\design_top.MEM[11][3] ),
    .A1(\design_top.MEM[10][3] ),
    .A2(\design_top.MEM[9][3] ),
    .A3(\design_top.MEM[8][3] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14177_ (.A0(\design_top.MEM[7][3] ),
    .A1(\design_top.MEM[6][3] ),
    .A2(\design_top.MEM[5][3] ),
    .A3(\design_top.MEM[4][3] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14178_ (.A0(\design_top.MEM[3][3] ),
    .A1(\design_top.MEM[2][3] ),
    .A2(\design_top.MEM[1][3] ),
    .A3(\design_top.MEM[0][3] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14179_ (.A0(_01127_),
    .A1(_01126_),
    .A2(_01125_),
    .A3(_01124_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14180_ (.A0(\design_top.MEM[15][2] ),
    .A1(\design_top.MEM[14][2] ),
    .A2(\design_top.MEM[13][2] ),
    .A3(\design_top.MEM[12][2] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14181_ (.A0(\design_top.MEM[11][2] ),
    .A1(\design_top.MEM[10][2] ),
    .A2(\design_top.MEM[9][2] ),
    .A3(\design_top.MEM[8][2] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14182_ (.A0(\design_top.MEM[7][2] ),
    .A1(\design_top.MEM[6][2] ),
    .A2(\design_top.MEM[5][2] ),
    .A3(\design_top.MEM[4][2] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14183_ (.A0(\design_top.MEM[3][2] ),
    .A1(\design_top.MEM[2][2] ),
    .A2(\design_top.MEM[1][2] ),
    .A3(\design_top.MEM[0][2] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14184_ (.A0(_01123_),
    .A1(_01122_),
    .A2(_01121_),
    .A3(_01120_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14185_ (.A0(\design_top.MEM[15][1] ),
    .A1(\design_top.MEM[14][1] ),
    .A2(\design_top.MEM[13][1] ),
    .A3(\design_top.MEM[12][1] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14186_ (.A0(\design_top.MEM[11][1] ),
    .A1(\design_top.MEM[10][1] ),
    .A2(\design_top.MEM[9][1] ),
    .A3(\design_top.MEM[8][1] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14187_ (.A0(\design_top.MEM[7][1] ),
    .A1(\design_top.MEM[6][1] ),
    .A2(\design_top.MEM[5][1] ),
    .A3(\design_top.MEM[4][1] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14188_ (.A0(\design_top.MEM[3][1] ),
    .A1(\design_top.MEM[2][1] ),
    .A2(\design_top.MEM[1][1] ),
    .A3(\design_top.MEM[0][1] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14189_ (.A0(_01119_),
    .A1(_01118_),
    .A2(_01117_),
    .A3(_01116_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14190_ (.A0(\design_top.MEM[15][0] ),
    .A1(\design_top.MEM[14][0] ),
    .A2(\design_top.MEM[13][0] ),
    .A3(\design_top.MEM[12][0] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14191_ (.A0(\design_top.MEM[11][0] ),
    .A1(\design_top.MEM[10][0] ),
    .A2(\design_top.MEM[9][0] ),
    .A3(\design_top.MEM[8][0] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14192_ (.A0(\design_top.MEM[7][0] ),
    .A1(\design_top.MEM[6][0] ),
    .A2(\design_top.MEM[5][0] ),
    .A3(\design_top.MEM[4][0] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14193_ (.A0(\design_top.MEM[3][0] ),
    .A1(\design_top.MEM[2][0] ),
    .A2(\design_top.MEM[1][0] ),
    .A3(\design_top.MEM[0][0] ),
    .S0(_00334_),
    .S1(_00343_),
    .X(_01112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14194_ (.A0(_01115_),
    .A1(_01114_),
    .A2(_01113_),
    .A3(_01112_),
    .S0(_00353_),
    .S1(_00360_),
    .X(_00109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14195_ (.A0(\design_top.MEM[0][31] ),
    .A1(\design_top.MEM[1][31] ),
    .A2(\design_top.MEM[2][31] ),
    .A3(\design_top.MEM[3][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14196_ (.A0(\design_top.MEM[4][31] ),
    .A1(\design_top.MEM[5][31] ),
    .A2(\design_top.MEM[6][31] ),
    .A3(\design_top.MEM[7][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14197_ (.A0(\design_top.MEM[8][31] ),
    .A1(\design_top.MEM[9][31] ),
    .A2(\design_top.MEM[10][31] ),
    .A3(\design_top.MEM[11][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14198_ (.A0(\design_top.MEM[12][31] ),
    .A1(\design_top.MEM[13][31] ),
    .A2(\design_top.MEM[14][31] ),
    .A3(\design_top.MEM[15][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14199_ (.A0(_01051_),
    .A1(_01052_),
    .A2(_01053_),
    .A3(_01054_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14200_ (.A0(\design_top.MEM[0][30] ),
    .A1(\design_top.MEM[1][30] ),
    .A2(\design_top.MEM[2][30] ),
    .A3(\design_top.MEM[3][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14201_ (.A0(\design_top.MEM[4][30] ),
    .A1(\design_top.MEM[5][30] ),
    .A2(\design_top.MEM[6][30] ),
    .A3(\design_top.MEM[7][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14202_ (.A0(\design_top.MEM[8][30] ),
    .A1(\design_top.MEM[9][30] ),
    .A2(\design_top.MEM[10][30] ),
    .A3(\design_top.MEM[11][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14203_ (.A0(\design_top.MEM[12][30] ),
    .A1(\design_top.MEM[13][30] ),
    .A2(\design_top.MEM[14][30] ),
    .A3(\design_top.MEM[15][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14204_ (.A0(_01047_),
    .A1(_01048_),
    .A2(_01049_),
    .A3(_01050_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14205_ (.A0(\design_top.MEM[0][29] ),
    .A1(\design_top.MEM[1][29] ),
    .A2(\design_top.MEM[2][29] ),
    .A3(\design_top.MEM[3][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14206_ (.A0(\design_top.MEM[4][29] ),
    .A1(\design_top.MEM[5][29] ),
    .A2(\design_top.MEM[6][29] ),
    .A3(\design_top.MEM[7][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14207_ (.A0(\design_top.MEM[8][29] ),
    .A1(\design_top.MEM[9][29] ),
    .A2(\design_top.MEM[10][29] ),
    .A3(\design_top.MEM[11][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14208_ (.A0(\design_top.MEM[12][29] ),
    .A1(\design_top.MEM[13][29] ),
    .A2(\design_top.MEM[14][29] ),
    .A3(\design_top.MEM[15][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14209_ (.A0(_01043_),
    .A1(_01044_),
    .A2(_01045_),
    .A3(_01046_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14210_ (.A0(\design_top.MEM[0][28] ),
    .A1(\design_top.MEM[1][28] ),
    .A2(\design_top.MEM[2][28] ),
    .A3(\design_top.MEM[3][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14211_ (.A0(\design_top.MEM[4][28] ),
    .A1(\design_top.MEM[5][28] ),
    .A2(\design_top.MEM[6][28] ),
    .A3(\design_top.MEM[7][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14212_ (.A0(\design_top.MEM[8][28] ),
    .A1(\design_top.MEM[9][28] ),
    .A2(\design_top.MEM[10][28] ),
    .A3(\design_top.MEM[11][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14213_ (.A0(\design_top.MEM[12][28] ),
    .A1(\design_top.MEM[13][28] ),
    .A2(\design_top.MEM[14][28] ),
    .A3(\design_top.MEM[15][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14214_ (.A0(_01039_),
    .A1(_01040_),
    .A2(_01041_),
    .A3(_01042_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14215_ (.A0(\design_top.MEM[0][27] ),
    .A1(\design_top.MEM[1][27] ),
    .A2(\design_top.MEM[2][27] ),
    .A3(\design_top.MEM[3][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14216_ (.A0(\design_top.MEM[4][27] ),
    .A1(\design_top.MEM[5][27] ),
    .A2(\design_top.MEM[6][27] ),
    .A3(\design_top.MEM[7][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14217_ (.A0(\design_top.MEM[8][27] ),
    .A1(\design_top.MEM[9][27] ),
    .A2(\design_top.MEM[10][27] ),
    .A3(\design_top.MEM[11][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14218_ (.A0(\design_top.MEM[12][27] ),
    .A1(\design_top.MEM[13][27] ),
    .A2(\design_top.MEM[14][27] ),
    .A3(\design_top.MEM[15][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14219_ (.A0(_01035_),
    .A1(_01036_),
    .A2(_01037_),
    .A3(_01038_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14220_ (.A0(\design_top.MEM[0][26] ),
    .A1(\design_top.MEM[1][26] ),
    .A2(\design_top.MEM[2][26] ),
    .A3(\design_top.MEM[3][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14221_ (.A0(\design_top.MEM[4][26] ),
    .A1(\design_top.MEM[5][26] ),
    .A2(\design_top.MEM[6][26] ),
    .A3(\design_top.MEM[7][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14222_ (.A0(\design_top.MEM[8][26] ),
    .A1(\design_top.MEM[9][26] ),
    .A2(\design_top.MEM[10][26] ),
    .A3(\design_top.MEM[11][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14223_ (.A0(\design_top.MEM[12][26] ),
    .A1(\design_top.MEM[13][26] ),
    .A2(\design_top.MEM[14][26] ),
    .A3(\design_top.MEM[15][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14224_ (.A0(_01031_),
    .A1(_01032_),
    .A2(_01033_),
    .A3(_01034_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14225_ (.A0(\design_top.MEM[0][25] ),
    .A1(\design_top.MEM[1][25] ),
    .A2(\design_top.MEM[2][25] ),
    .A3(\design_top.MEM[3][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14226_ (.A0(\design_top.MEM[4][25] ),
    .A1(\design_top.MEM[5][25] ),
    .A2(\design_top.MEM[6][25] ),
    .A3(\design_top.MEM[7][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14227_ (.A0(\design_top.MEM[8][25] ),
    .A1(\design_top.MEM[9][25] ),
    .A2(\design_top.MEM[10][25] ),
    .A3(\design_top.MEM[11][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14228_ (.A0(\design_top.MEM[12][25] ),
    .A1(\design_top.MEM[13][25] ),
    .A2(\design_top.MEM[14][25] ),
    .A3(\design_top.MEM[15][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14229_ (.A0(_01027_),
    .A1(_01028_),
    .A2(_01029_),
    .A3(_01030_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14230_ (.A0(\design_top.MEM[0][24] ),
    .A1(\design_top.MEM[1][24] ),
    .A2(\design_top.MEM[2][24] ),
    .A3(\design_top.MEM[3][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14231_ (.A0(\design_top.MEM[4][24] ),
    .A1(\design_top.MEM[5][24] ),
    .A2(\design_top.MEM[6][24] ),
    .A3(\design_top.MEM[7][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14232_ (.A0(\design_top.MEM[8][24] ),
    .A1(\design_top.MEM[9][24] ),
    .A2(\design_top.MEM[10][24] ),
    .A3(\design_top.MEM[11][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14233_ (.A0(\design_top.MEM[12][24] ),
    .A1(\design_top.MEM[13][24] ),
    .A2(\design_top.MEM[14][24] ),
    .A3(\design_top.MEM[15][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14234_ (.A0(_01023_),
    .A1(_01024_),
    .A2(_01025_),
    .A3(_01026_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14235_ (.A0(\design_top.MEM[0][23] ),
    .A1(\design_top.MEM[1][23] ),
    .A2(\design_top.MEM[2][23] ),
    .A3(\design_top.MEM[3][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14236_ (.A0(\design_top.MEM[4][23] ),
    .A1(\design_top.MEM[5][23] ),
    .A2(\design_top.MEM[6][23] ),
    .A3(\design_top.MEM[7][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14237_ (.A0(\design_top.MEM[8][23] ),
    .A1(\design_top.MEM[9][23] ),
    .A2(\design_top.MEM[10][23] ),
    .A3(\design_top.MEM[11][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14238_ (.A0(\design_top.MEM[12][23] ),
    .A1(\design_top.MEM[13][23] ),
    .A2(\design_top.MEM[14][23] ),
    .A3(\design_top.MEM[15][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14239_ (.A0(_01019_),
    .A1(_01020_),
    .A2(_01021_),
    .A3(_01022_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14240_ (.A0(\design_top.MEM[0][22] ),
    .A1(\design_top.MEM[1][22] ),
    .A2(\design_top.MEM[2][22] ),
    .A3(\design_top.MEM[3][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14241_ (.A0(\design_top.MEM[4][22] ),
    .A1(\design_top.MEM[5][22] ),
    .A2(\design_top.MEM[6][22] ),
    .A3(\design_top.MEM[7][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14242_ (.A0(\design_top.MEM[8][22] ),
    .A1(\design_top.MEM[9][22] ),
    .A2(\design_top.MEM[10][22] ),
    .A3(\design_top.MEM[11][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14243_ (.A0(\design_top.MEM[12][22] ),
    .A1(\design_top.MEM[13][22] ),
    .A2(\design_top.MEM[14][22] ),
    .A3(\design_top.MEM[15][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14244_ (.A0(_01015_),
    .A1(_01016_),
    .A2(_01017_),
    .A3(_01018_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14245_ (.A0(\design_top.MEM[0][21] ),
    .A1(\design_top.MEM[1][21] ),
    .A2(\design_top.MEM[2][21] ),
    .A3(\design_top.MEM[3][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14246_ (.A0(\design_top.MEM[4][21] ),
    .A1(\design_top.MEM[5][21] ),
    .A2(\design_top.MEM[6][21] ),
    .A3(\design_top.MEM[7][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14247_ (.A0(\design_top.MEM[8][21] ),
    .A1(\design_top.MEM[9][21] ),
    .A2(\design_top.MEM[10][21] ),
    .A3(\design_top.MEM[11][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14248_ (.A0(\design_top.MEM[12][21] ),
    .A1(\design_top.MEM[13][21] ),
    .A2(\design_top.MEM[14][21] ),
    .A3(\design_top.MEM[15][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14249_ (.A0(_01011_),
    .A1(_01012_),
    .A2(_01013_),
    .A3(_01014_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14250_ (.A0(\design_top.MEM[0][20] ),
    .A1(\design_top.MEM[1][20] ),
    .A2(\design_top.MEM[2][20] ),
    .A3(\design_top.MEM[3][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14251_ (.A0(\design_top.MEM[4][20] ),
    .A1(\design_top.MEM[5][20] ),
    .A2(\design_top.MEM[6][20] ),
    .A3(\design_top.MEM[7][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14252_ (.A0(\design_top.MEM[8][20] ),
    .A1(\design_top.MEM[9][20] ),
    .A2(\design_top.MEM[10][20] ),
    .A3(\design_top.MEM[11][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14253_ (.A0(\design_top.MEM[12][20] ),
    .A1(\design_top.MEM[13][20] ),
    .A2(\design_top.MEM[14][20] ),
    .A3(\design_top.MEM[15][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14254_ (.A0(_01007_),
    .A1(_01008_),
    .A2(_01009_),
    .A3(_01010_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14255_ (.A0(\design_top.MEM[0][19] ),
    .A1(\design_top.MEM[1][19] ),
    .A2(\design_top.MEM[2][19] ),
    .A3(\design_top.MEM[3][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14256_ (.A0(\design_top.MEM[4][19] ),
    .A1(\design_top.MEM[5][19] ),
    .A2(\design_top.MEM[6][19] ),
    .A3(\design_top.MEM[7][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14257_ (.A0(\design_top.MEM[8][19] ),
    .A1(\design_top.MEM[9][19] ),
    .A2(\design_top.MEM[10][19] ),
    .A3(\design_top.MEM[11][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14258_ (.A0(\design_top.MEM[12][19] ),
    .A1(\design_top.MEM[13][19] ),
    .A2(\design_top.MEM[14][19] ),
    .A3(\design_top.MEM[15][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14259_ (.A0(_01003_),
    .A1(_01004_),
    .A2(_01005_),
    .A3(_01006_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14260_ (.A0(\design_top.MEM[0][18] ),
    .A1(\design_top.MEM[1][18] ),
    .A2(\design_top.MEM[2][18] ),
    .A3(\design_top.MEM[3][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14261_ (.A0(\design_top.MEM[4][18] ),
    .A1(\design_top.MEM[5][18] ),
    .A2(\design_top.MEM[6][18] ),
    .A3(\design_top.MEM[7][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14262_ (.A0(\design_top.MEM[8][18] ),
    .A1(\design_top.MEM[9][18] ),
    .A2(\design_top.MEM[10][18] ),
    .A3(\design_top.MEM[11][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14263_ (.A0(\design_top.MEM[12][18] ),
    .A1(\design_top.MEM[13][18] ),
    .A2(\design_top.MEM[14][18] ),
    .A3(\design_top.MEM[15][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_01002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14264_ (.A0(_00999_),
    .A1(_01000_),
    .A2(_01001_),
    .A3(_01002_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14265_ (.A0(\design_top.MEM[0][17] ),
    .A1(\design_top.MEM[1][17] ),
    .A2(\design_top.MEM[2][17] ),
    .A3(\design_top.MEM[3][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14266_ (.A0(\design_top.MEM[4][17] ),
    .A1(\design_top.MEM[5][17] ),
    .A2(\design_top.MEM[6][17] ),
    .A3(\design_top.MEM[7][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14267_ (.A0(\design_top.MEM[8][17] ),
    .A1(\design_top.MEM[9][17] ),
    .A2(\design_top.MEM[10][17] ),
    .A3(\design_top.MEM[11][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14268_ (.A0(\design_top.MEM[12][17] ),
    .A1(\design_top.MEM[13][17] ),
    .A2(\design_top.MEM[14][17] ),
    .A3(\design_top.MEM[15][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14269_ (.A0(_00995_),
    .A1(_00996_),
    .A2(_00997_),
    .A3(_00998_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14270_ (.A0(\design_top.MEM[0][16] ),
    .A1(\design_top.MEM[1][16] ),
    .A2(\design_top.MEM[2][16] ),
    .A3(\design_top.MEM[3][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14271_ (.A0(\design_top.MEM[4][16] ),
    .A1(\design_top.MEM[5][16] ),
    .A2(\design_top.MEM[6][16] ),
    .A3(\design_top.MEM[7][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14272_ (.A0(\design_top.MEM[8][16] ),
    .A1(\design_top.MEM[9][16] ),
    .A2(\design_top.MEM[10][16] ),
    .A3(\design_top.MEM[11][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14273_ (.A0(\design_top.MEM[12][16] ),
    .A1(\design_top.MEM[13][16] ),
    .A2(\design_top.MEM[14][16] ),
    .A3(\design_top.MEM[15][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14274_ (.A0(_00991_),
    .A1(_00992_),
    .A2(_00993_),
    .A3(_00994_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14275_ (.A0(\design_top.MEM[0][15] ),
    .A1(\design_top.MEM[1][15] ),
    .A2(\design_top.MEM[2][15] ),
    .A3(\design_top.MEM[3][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14276_ (.A0(\design_top.MEM[4][15] ),
    .A1(\design_top.MEM[5][15] ),
    .A2(\design_top.MEM[6][15] ),
    .A3(\design_top.MEM[7][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14277_ (.A0(\design_top.MEM[8][15] ),
    .A1(\design_top.MEM[9][15] ),
    .A2(\design_top.MEM[10][15] ),
    .A3(\design_top.MEM[11][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14278_ (.A0(\design_top.MEM[12][15] ),
    .A1(\design_top.MEM[13][15] ),
    .A2(\design_top.MEM[14][15] ),
    .A3(\design_top.MEM[15][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14279_ (.A0(_00987_),
    .A1(_00988_),
    .A2(_00989_),
    .A3(_00990_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14280_ (.A0(\design_top.MEM[0][14] ),
    .A1(\design_top.MEM[1][14] ),
    .A2(\design_top.MEM[2][14] ),
    .A3(\design_top.MEM[3][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14281_ (.A0(\design_top.MEM[4][14] ),
    .A1(\design_top.MEM[5][14] ),
    .A2(\design_top.MEM[6][14] ),
    .A3(\design_top.MEM[7][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14282_ (.A0(\design_top.MEM[8][14] ),
    .A1(\design_top.MEM[9][14] ),
    .A2(\design_top.MEM[10][14] ),
    .A3(\design_top.MEM[11][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14283_ (.A0(\design_top.MEM[12][14] ),
    .A1(\design_top.MEM[13][14] ),
    .A2(\design_top.MEM[14][14] ),
    .A3(\design_top.MEM[15][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14284_ (.A0(_00983_),
    .A1(_00984_),
    .A2(_00985_),
    .A3(_00986_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14285_ (.A0(\design_top.MEM[0][13] ),
    .A1(\design_top.MEM[1][13] ),
    .A2(\design_top.MEM[2][13] ),
    .A3(\design_top.MEM[3][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14286_ (.A0(\design_top.MEM[4][13] ),
    .A1(\design_top.MEM[5][13] ),
    .A2(\design_top.MEM[6][13] ),
    .A3(\design_top.MEM[7][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14287_ (.A0(\design_top.MEM[8][13] ),
    .A1(\design_top.MEM[9][13] ),
    .A2(\design_top.MEM[10][13] ),
    .A3(\design_top.MEM[11][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14288_ (.A0(\design_top.MEM[12][13] ),
    .A1(\design_top.MEM[13][13] ),
    .A2(\design_top.MEM[14][13] ),
    .A3(\design_top.MEM[15][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14289_ (.A0(_00979_),
    .A1(_00980_),
    .A2(_00981_),
    .A3(_00982_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14290_ (.A0(\design_top.MEM[0][12] ),
    .A1(\design_top.MEM[1][12] ),
    .A2(\design_top.MEM[2][12] ),
    .A3(\design_top.MEM[3][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14291_ (.A0(\design_top.MEM[4][12] ),
    .A1(\design_top.MEM[5][12] ),
    .A2(\design_top.MEM[6][12] ),
    .A3(\design_top.MEM[7][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14292_ (.A0(\design_top.MEM[8][12] ),
    .A1(\design_top.MEM[9][12] ),
    .A2(\design_top.MEM[10][12] ),
    .A3(\design_top.MEM[11][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14293_ (.A0(\design_top.MEM[12][12] ),
    .A1(\design_top.MEM[13][12] ),
    .A2(\design_top.MEM[14][12] ),
    .A3(\design_top.MEM[15][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14294_ (.A0(_00975_),
    .A1(_00976_),
    .A2(_00977_),
    .A3(_00978_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14295_ (.A0(\design_top.MEM[0][11] ),
    .A1(\design_top.MEM[1][11] ),
    .A2(\design_top.MEM[2][11] ),
    .A3(\design_top.MEM[3][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14296_ (.A0(\design_top.MEM[4][11] ),
    .A1(\design_top.MEM[5][11] ),
    .A2(\design_top.MEM[6][11] ),
    .A3(\design_top.MEM[7][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14297_ (.A0(\design_top.MEM[8][11] ),
    .A1(\design_top.MEM[9][11] ),
    .A2(\design_top.MEM[10][11] ),
    .A3(\design_top.MEM[11][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14298_ (.A0(\design_top.MEM[12][11] ),
    .A1(\design_top.MEM[13][11] ),
    .A2(\design_top.MEM[14][11] ),
    .A3(\design_top.MEM[15][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14299_ (.A0(_00971_),
    .A1(_00972_),
    .A2(_00973_),
    .A3(_00974_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14300_ (.A0(\design_top.MEM[0][10] ),
    .A1(\design_top.MEM[1][10] ),
    .A2(\design_top.MEM[2][10] ),
    .A3(\design_top.MEM[3][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14301_ (.A0(\design_top.MEM[4][10] ),
    .A1(\design_top.MEM[5][10] ),
    .A2(\design_top.MEM[6][10] ),
    .A3(\design_top.MEM[7][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14302_ (.A0(\design_top.MEM[8][10] ),
    .A1(\design_top.MEM[9][10] ),
    .A2(\design_top.MEM[10][10] ),
    .A3(\design_top.MEM[11][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14303_ (.A0(\design_top.MEM[12][10] ),
    .A1(\design_top.MEM[13][10] ),
    .A2(\design_top.MEM[14][10] ),
    .A3(\design_top.MEM[15][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14304_ (.A0(_00967_),
    .A1(_00968_),
    .A2(_00969_),
    .A3(_00970_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14305_ (.A0(\design_top.MEM[0][9] ),
    .A1(\design_top.MEM[1][9] ),
    .A2(\design_top.MEM[2][9] ),
    .A3(\design_top.MEM[3][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14306_ (.A0(\design_top.MEM[4][9] ),
    .A1(\design_top.MEM[5][9] ),
    .A2(\design_top.MEM[6][9] ),
    .A3(\design_top.MEM[7][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14307_ (.A0(\design_top.MEM[8][9] ),
    .A1(\design_top.MEM[9][9] ),
    .A2(\design_top.MEM[10][9] ),
    .A3(\design_top.MEM[11][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14308_ (.A0(\design_top.MEM[12][9] ),
    .A1(\design_top.MEM[13][9] ),
    .A2(\design_top.MEM[14][9] ),
    .A3(\design_top.MEM[15][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14309_ (.A0(_00963_),
    .A1(_00964_),
    .A2(_00965_),
    .A3(_00966_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14310_ (.A0(\design_top.MEM[0][8] ),
    .A1(\design_top.MEM[1][8] ),
    .A2(\design_top.MEM[2][8] ),
    .A3(\design_top.MEM[3][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14311_ (.A0(\design_top.MEM[4][8] ),
    .A1(\design_top.MEM[5][8] ),
    .A2(\design_top.MEM[6][8] ),
    .A3(\design_top.MEM[7][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14312_ (.A0(\design_top.MEM[8][8] ),
    .A1(\design_top.MEM[9][8] ),
    .A2(\design_top.MEM[10][8] ),
    .A3(\design_top.MEM[11][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14313_ (.A0(\design_top.MEM[12][8] ),
    .A1(\design_top.MEM[13][8] ),
    .A2(\design_top.MEM[14][8] ),
    .A3(\design_top.MEM[15][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14314_ (.A0(_00959_),
    .A1(_00960_),
    .A2(_00961_),
    .A3(_00962_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14315_ (.A0(\design_top.MEM[0][7] ),
    .A1(\design_top.MEM[1][7] ),
    .A2(\design_top.MEM[2][7] ),
    .A3(\design_top.MEM[3][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14316_ (.A0(\design_top.MEM[4][7] ),
    .A1(\design_top.MEM[5][7] ),
    .A2(\design_top.MEM[6][7] ),
    .A3(\design_top.MEM[7][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14317_ (.A0(\design_top.MEM[8][7] ),
    .A1(\design_top.MEM[9][7] ),
    .A2(\design_top.MEM[10][7] ),
    .A3(\design_top.MEM[11][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14318_ (.A0(\design_top.MEM[12][7] ),
    .A1(\design_top.MEM[13][7] ),
    .A2(\design_top.MEM[14][7] ),
    .A3(\design_top.MEM[15][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14319_ (.A0(_00955_),
    .A1(_00956_),
    .A2(_00957_),
    .A3(_00958_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14320_ (.A0(\design_top.MEM[0][6] ),
    .A1(\design_top.MEM[1][6] ),
    .A2(\design_top.MEM[2][6] ),
    .A3(\design_top.MEM[3][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14321_ (.A0(\design_top.MEM[4][6] ),
    .A1(\design_top.MEM[5][6] ),
    .A2(\design_top.MEM[6][6] ),
    .A3(\design_top.MEM[7][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14322_ (.A0(\design_top.MEM[8][6] ),
    .A1(\design_top.MEM[9][6] ),
    .A2(\design_top.MEM[10][6] ),
    .A3(\design_top.MEM[11][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14323_ (.A0(\design_top.MEM[12][6] ),
    .A1(\design_top.MEM[13][6] ),
    .A2(\design_top.MEM[14][6] ),
    .A3(\design_top.MEM[15][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14324_ (.A0(_00951_),
    .A1(_00952_),
    .A2(_00953_),
    .A3(_00954_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14325_ (.A0(\design_top.MEM[0][5] ),
    .A1(\design_top.MEM[1][5] ),
    .A2(\design_top.MEM[2][5] ),
    .A3(\design_top.MEM[3][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14326_ (.A0(\design_top.MEM[4][5] ),
    .A1(\design_top.MEM[5][5] ),
    .A2(\design_top.MEM[6][5] ),
    .A3(\design_top.MEM[7][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14327_ (.A0(\design_top.MEM[8][5] ),
    .A1(\design_top.MEM[9][5] ),
    .A2(\design_top.MEM[10][5] ),
    .A3(\design_top.MEM[11][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14328_ (.A0(\design_top.MEM[12][5] ),
    .A1(\design_top.MEM[13][5] ),
    .A2(\design_top.MEM[14][5] ),
    .A3(\design_top.MEM[15][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14329_ (.A0(_00947_),
    .A1(_00948_),
    .A2(_00949_),
    .A3(_00950_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14330_ (.A0(\design_top.MEM[0][4] ),
    .A1(\design_top.MEM[1][4] ),
    .A2(\design_top.MEM[2][4] ),
    .A3(\design_top.MEM[3][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14331_ (.A0(\design_top.MEM[4][4] ),
    .A1(\design_top.MEM[5][4] ),
    .A2(\design_top.MEM[6][4] ),
    .A3(\design_top.MEM[7][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14332_ (.A0(\design_top.MEM[8][4] ),
    .A1(\design_top.MEM[9][4] ),
    .A2(\design_top.MEM[10][4] ),
    .A3(\design_top.MEM[11][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14333_ (.A0(\design_top.MEM[12][4] ),
    .A1(\design_top.MEM[13][4] ),
    .A2(\design_top.MEM[14][4] ),
    .A3(\design_top.MEM[15][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14334_ (.A0(_00943_),
    .A1(_00944_),
    .A2(_00945_),
    .A3(_00946_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14335_ (.A0(\design_top.MEM[0][3] ),
    .A1(\design_top.MEM[1][3] ),
    .A2(\design_top.MEM[2][3] ),
    .A3(\design_top.MEM[3][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14336_ (.A0(\design_top.MEM[4][3] ),
    .A1(\design_top.MEM[5][3] ),
    .A2(\design_top.MEM[6][3] ),
    .A3(\design_top.MEM[7][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14337_ (.A0(\design_top.MEM[8][3] ),
    .A1(\design_top.MEM[9][3] ),
    .A2(\design_top.MEM[10][3] ),
    .A3(\design_top.MEM[11][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14338_ (.A0(\design_top.MEM[12][3] ),
    .A1(\design_top.MEM[13][3] ),
    .A2(\design_top.MEM[14][3] ),
    .A3(\design_top.MEM[15][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14339_ (.A0(_00939_),
    .A1(_00940_),
    .A2(_00941_),
    .A3(_00942_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14340_ (.A0(\design_top.MEM[0][2] ),
    .A1(\design_top.MEM[1][2] ),
    .A2(\design_top.MEM[2][2] ),
    .A3(\design_top.MEM[3][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14341_ (.A0(\design_top.MEM[4][2] ),
    .A1(\design_top.MEM[5][2] ),
    .A2(\design_top.MEM[6][2] ),
    .A3(\design_top.MEM[7][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14342_ (.A0(\design_top.MEM[8][2] ),
    .A1(\design_top.MEM[9][2] ),
    .A2(\design_top.MEM[10][2] ),
    .A3(\design_top.MEM[11][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14343_ (.A0(\design_top.MEM[12][2] ),
    .A1(\design_top.MEM[13][2] ),
    .A2(\design_top.MEM[14][2] ),
    .A3(\design_top.MEM[15][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14344_ (.A0(_00935_),
    .A1(_00936_),
    .A2(_00937_),
    .A3(_00938_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14345_ (.A0(\design_top.MEM[0][1] ),
    .A1(\design_top.MEM[1][1] ),
    .A2(\design_top.MEM[2][1] ),
    .A3(\design_top.MEM[3][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14346_ (.A0(\design_top.MEM[4][1] ),
    .A1(\design_top.MEM[5][1] ),
    .A2(\design_top.MEM[6][1] ),
    .A3(\design_top.MEM[7][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14347_ (.A0(\design_top.MEM[8][1] ),
    .A1(\design_top.MEM[9][1] ),
    .A2(\design_top.MEM[10][1] ),
    .A3(\design_top.MEM[11][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14348_ (.A0(\design_top.MEM[12][1] ),
    .A1(\design_top.MEM[13][1] ),
    .A2(\design_top.MEM[14][1] ),
    .A3(\design_top.MEM[15][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14349_ (.A0(_00931_),
    .A1(_00932_),
    .A2(_00933_),
    .A3(_00934_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14350_ (.A0(\design_top.MEM[0][0] ),
    .A1(\design_top.MEM[1][0] ),
    .A2(\design_top.MEM[2][0] ),
    .A3(\design_top.MEM[3][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14351_ (.A0(\design_top.MEM[4][0] ),
    .A1(\design_top.MEM[5][0] ),
    .A2(\design_top.MEM[6][0] ),
    .A3(\design_top.MEM[7][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14352_ (.A0(\design_top.MEM[8][0] ),
    .A1(\design_top.MEM[9][0] ),
    .A2(\design_top.MEM[10][0] ),
    .A3(\design_top.MEM[11][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14353_ (.A0(\design_top.MEM[12][0] ),
    .A1(\design_top.MEM[13][0] ),
    .A2(\design_top.MEM[14][0] ),
    .A3(\design_top.MEM[15][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _14354_ (.A0(_00927_),
    .A1(_00928_),
    .A2(_00929_),
    .A3(_00930_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14355_ (.D(_00046_),
    .Q(\design_top.core0.XRES ),
    .CLK(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14356_ (.D(io_in[1]),
    .Q(\design_top.uart0.UART_RXDFF[0] ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14357_ (.D(\design_top.uart0.UART_RXDFF[0] ),
    .Q(\design_top.uart0.UART_RXDFF[1] ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14358_ (.D(\design_top.uart0.UART_RXDFF[1] ),
    .Q(\design_top.uart0.UART_RXDFF[2] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14359_ (.D(\design_top.XRES_reg ),
    .Q(\design_top.XRES ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14360_ (.D(io_in[0]),
    .Q(\design_top.XRES_reg ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14361_ (.D(\design_top.HLT ),
    .Q(\design_top.HLT2 ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14362_ (.D(\design_top.DADDR[2] ),
    .Q(\design_top.XADDR[2] ),
    .CLK(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14363_ (.D(\design_top.DADDR[3] ),
    .Q(\design_top.XADDR[3] ),
    .CLK(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14364_ (.D(\design_top.DADDR[31] ),
    .Q(\design_top.XADDR[31] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14365_ (.D(_00141_),
    .Q(\design_top.ROMFF[0] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14366_ (.D(_00152_),
    .Q(\design_top.ROMFF[1] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14367_ (.D(_00163_),
    .Q(\design_top.ROMFF[2] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14368_ (.D(_00166_),
    .Q(\design_top.ROMFF[3] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14369_ (.D(_00167_),
    .Q(\design_top.ROMFF[4] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14370_ (.D(_00168_),
    .Q(\design_top.ROMFF[5] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14371_ (.D(_00169_),
    .Q(\design_top.ROMFF[6] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14372_ (.D(_00170_),
    .Q(\design_top.ROMFF[7] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14373_ (.D(_00171_),
    .Q(\design_top.ROMFF[8] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14374_ (.D(_00172_),
    .Q(\design_top.ROMFF[9] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14375_ (.D(_00142_),
    .Q(\design_top.ROMFF[10] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14376_ (.D(_00143_),
    .Q(\design_top.ROMFF[11] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14377_ (.D(_00144_),
    .Q(\design_top.ROMFF[12] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14378_ (.D(_00145_),
    .Q(\design_top.ROMFF[13] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14379_ (.D(_00146_),
    .Q(\design_top.ROMFF[14] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14380_ (.D(_00147_),
    .Q(\design_top.ROMFF[15] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14381_ (.D(_00148_),
    .Q(\design_top.ROMFF[16] ),
    .CLK(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14382_ (.D(_00149_),
    .Q(\design_top.ROMFF[17] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14383_ (.D(_00150_),
    .Q(\design_top.ROMFF[18] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14384_ (.D(_00151_),
    .Q(\design_top.ROMFF[19] ),
    .CLK(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14385_ (.D(_00153_),
    .Q(\design_top.ROMFF[20] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14386_ (.D(_00154_),
    .Q(\design_top.ROMFF[21] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14387_ (.D(_00155_),
    .Q(\design_top.ROMFF[22] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14388_ (.D(_00156_),
    .Q(\design_top.ROMFF[23] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14389_ (.D(_00157_),
    .Q(\design_top.ROMFF[24] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14390_ (.D(_00158_),
    .Q(\design_top.ROMFF[25] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14391_ (.D(_00159_),
    .Q(\design_top.ROMFF[26] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14392_ (.D(_00160_),
    .Q(\design_top.ROMFF[27] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14393_ (.D(_00161_),
    .Q(\design_top.ROMFF[28] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14394_ (.D(_00162_),
    .Q(\design_top.ROMFF[29] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14395_ (.D(_00164_),
    .Q(\design_top.ROMFF[30] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14396_ (.D(_00165_),
    .Q(\design_top.ROMFF[31] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14397_ (.D(_00109_),
    .Q(\design_top.RAMFF[0] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14398_ (.D(_00120_),
    .Q(\design_top.RAMFF[1] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14399_ (.D(_00131_),
    .Q(\design_top.RAMFF[2] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14400_ (.D(_00134_),
    .Q(\design_top.RAMFF[3] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14401_ (.D(_00135_),
    .Q(\design_top.RAMFF[4] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14402_ (.D(_00136_),
    .Q(\design_top.RAMFF[5] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14403_ (.D(_00137_),
    .Q(\design_top.RAMFF[6] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14404_ (.D(_00138_),
    .Q(\design_top.RAMFF[7] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14405_ (.D(_00139_),
    .Q(\design_top.RAMFF[8] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14406_ (.D(_00140_),
    .Q(\design_top.RAMFF[9] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14407_ (.D(_00110_),
    .Q(\design_top.RAMFF[10] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14408_ (.D(_00111_),
    .Q(\design_top.RAMFF[11] ),
    .CLK(clknet_leaf_235_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14409_ (.D(_00112_),
    .Q(\design_top.RAMFF[12] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14410_ (.D(_00113_),
    .Q(\design_top.RAMFF[13] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14411_ (.D(_00114_),
    .Q(\design_top.RAMFF[14] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14412_ (.D(_00115_),
    .Q(\design_top.RAMFF[15] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14413_ (.D(_00116_),
    .Q(\design_top.RAMFF[16] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14414_ (.D(_00117_),
    .Q(\design_top.RAMFF[17] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14415_ (.D(_00118_),
    .Q(\design_top.RAMFF[18] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14416_ (.D(_00119_),
    .Q(\design_top.RAMFF[19] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14417_ (.D(_00121_),
    .Q(\design_top.RAMFF[20] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14418_ (.D(_00122_),
    .Q(\design_top.RAMFF[21] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14419_ (.D(_00123_),
    .Q(\design_top.RAMFF[22] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14420_ (.D(_00124_),
    .Q(\design_top.RAMFF[23] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14421_ (.D(_00125_),
    .Q(\design_top.RAMFF[24] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14422_ (.D(_00126_),
    .Q(\design_top.RAMFF[25] ),
    .CLK(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14423_ (.D(_00127_),
    .Q(\design_top.RAMFF[26] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14424_ (.D(_00128_),
    .Q(\design_top.RAMFF[27] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14425_ (.D(_00129_),
    .Q(\design_top.RAMFF[28] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14426_ (.D(_00130_),
    .Q(\design_top.RAMFF[29] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14427_ (.D(_00132_),
    .Q(\design_top.RAMFF[30] ),
    .CLK(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14428_ (.D(_00133_),
    .Q(\design_top.RAMFF[31] ),
    .CLK(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14429_ (.D(_02514_),
    .Q(\design_top.core0.NXPC[0] ),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14430_ (.D(_02515_),
    .Q(\design_top.core0.NXPC[1] ),
    .CLK(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14431_ (.D(_02516_),
    .Q(\design_top.core0.NXPC[2] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14432_ (.D(_02517_),
    .Q(\design_top.core0.NXPC[3] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14433_ (.D(_02518_),
    .Q(\design_top.core0.NXPC[4] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14434_ (.D(_02519_),
    .Q(\design_top.core0.NXPC[5] ),
    .CLK(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14435_ (.D(_02520_),
    .Q(\design_top.core0.NXPC[6] ),
    .CLK(clknet_leaf_29_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14436_ (.D(_02521_),
    .Q(\design_top.core0.NXPC[7] ),
    .CLK(clknet_leaf_29_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14437_ (.D(_02522_),
    .Q(\design_top.core0.NXPC[8] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14438_ (.D(_02523_),
    .Q(\design_top.core0.NXPC[9] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14439_ (.D(_02524_),
    .Q(\design_top.core0.NXPC[10] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14440_ (.D(_02525_),
    .Q(\design_top.core0.NXPC[11] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14441_ (.D(_02526_),
    .Q(\design_top.core0.NXPC[12] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14442_ (.D(_02527_),
    .Q(\design_top.core0.NXPC[13] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14443_ (.D(_02528_),
    .Q(\design_top.core0.NXPC[14] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14444_ (.D(_02529_),
    .Q(\design_top.core0.NXPC[15] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14445_ (.D(_02530_),
    .Q(\design_top.core0.NXPC[16] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14446_ (.D(_02531_),
    .Q(\design_top.core0.NXPC[17] ),
    .CLK(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14447_ (.D(_02532_),
    .Q(\design_top.core0.NXPC[18] ),
    .CLK(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14448_ (.D(_02533_),
    .Q(\design_top.core0.NXPC[19] ),
    .CLK(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14449_ (.D(_02534_),
    .Q(\design_top.core0.NXPC[20] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14450_ (.D(_02535_),
    .Q(\design_top.core0.NXPC[21] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14451_ (.D(_02536_),
    .Q(\design_top.core0.NXPC[22] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14452_ (.D(_02537_),
    .Q(\design_top.core0.NXPC[23] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14453_ (.D(_02538_),
    .Q(\design_top.core0.NXPC[24] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14454_ (.D(_02539_),
    .Q(\design_top.core0.NXPC[25] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14455_ (.D(_02540_),
    .Q(\design_top.core0.NXPC[26] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14456_ (.D(_02541_),
    .Q(\design_top.core0.NXPC[27] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14457_ (.D(_02542_),
    .Q(\design_top.core0.NXPC[28] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14458_ (.D(_02543_),
    .Q(\design_top.core0.NXPC[29] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14459_ (.D(_02544_),
    .Q(\design_top.core0.NXPC[30] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14460_ (.D(_02545_),
    .Q(\design_top.core0.NXPC[31] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14461_ (.D(_02546_),
    .Q(\design_top.core0.PC[0] ),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14462_ (.D(_02547_),
    .Q(\design_top.core0.PC[1] ),
    .CLK(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14463_ (.D(_02548_),
    .Q(\design_top.core0.PC[2] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14464_ (.D(_02549_),
    .Q(\design_top.core0.PC[3] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14465_ (.D(_02550_),
    .Q(\design_top.core0.PC[4] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14466_ (.D(_02551_),
    .Q(\design_top.core0.PC[5] ),
    .CLK(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14467_ (.D(_02552_),
    .Q(\design_top.core0.PC[6] ),
    .CLK(clknet_leaf_29_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14468_ (.D(_02553_),
    .Q(\design_top.core0.PC[7] ),
    .CLK(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14469_ (.D(_02554_),
    .Q(\design_top.core0.PC[8] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14470_ (.D(_02555_),
    .Q(\design_top.core0.PC[9] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14471_ (.D(_02556_),
    .Q(\design_top.core0.PC[10] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14472_ (.D(_02557_),
    .Q(\design_top.core0.PC[11] ),
    .CLK(clknet_leaf_31_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14473_ (.D(_02558_),
    .Q(\design_top.core0.PC[12] ),
    .CLK(clknet_leaf_31_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14474_ (.D(_02559_),
    .Q(\design_top.core0.PC[13] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14475_ (.D(_02560_),
    .Q(\design_top.core0.PC[14] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14476_ (.D(_02561_),
    .Q(\design_top.core0.PC[15] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14477_ (.D(_02562_),
    .Q(\design_top.core0.PC[16] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14478_ (.D(_02563_),
    .Q(\design_top.core0.PC[17] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14479_ (.D(_02564_),
    .Q(\design_top.core0.PC[18] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14480_ (.D(_02565_),
    .Q(\design_top.core0.PC[19] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14481_ (.D(_02566_),
    .Q(\design_top.core0.PC[20] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14482_ (.D(_02567_),
    .Q(\design_top.core0.PC[21] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14483_ (.D(_02568_),
    .Q(\design_top.core0.PC[22] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14484_ (.D(_02569_),
    .Q(\design_top.core0.PC[23] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14485_ (.D(_02570_),
    .Q(\design_top.core0.PC[24] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14486_ (.D(_02571_),
    .Q(\design_top.core0.PC[25] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14487_ (.D(_02572_),
    .Q(\design_top.core0.PC[26] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14488_ (.D(_02573_),
    .Q(\design_top.core0.PC[27] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14489_ (.D(_02574_),
    .Q(\design_top.core0.PC[28] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14490_ (.D(_02575_),
    .Q(\design_top.core0.PC[29] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14491_ (.D(_02576_),
    .Q(\design_top.core0.PC[30] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14492_ (.D(_02577_),
    .Q(\design_top.core0.PC[31] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14493_ (.D(_02578_),
    .Q(\design_top.uart0.UART_RFIFO[0] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14494_ (.D(_02579_),
    .Q(\design_top.uart0.UART_RFIFO[1] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14495_ (.D(_02580_),
    .Q(\design_top.uart0.UART_RFIFO[2] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14496_ (.D(_02581_),
    .Q(\design_top.uart0.UART_RFIFO[3] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14497_ (.D(_02582_),
    .Q(\design_top.uart0.UART_RFIFO[4] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14498_ (.D(_02583_),
    .Q(\design_top.uart0.UART_RFIFO[5] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14499_ (.D(_02584_),
    .Q(\design_top.uart0.UART_RFIFO[6] ),
    .CLK(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14500_ (.D(_02585_),
    .Q(\design_top.uart0.UART_RFIFO[7] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14501_ (.D(_02586_),
    .Q(\design_top.uart0.UART_RREQ ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14502_ (.D(_02587_),
    .Q(\design_top.uart0.UART_XACK ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14503_ (.D(_02588_),
    .Q(\design_top.ROMFF2[0] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14504_ (.D(_02589_),
    .Q(\design_top.ROMFF2[1] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14505_ (.D(_02590_),
    .Q(\design_top.ROMFF2[2] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14506_ (.D(_02591_),
    .Q(\design_top.ROMFF2[3] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14507_ (.D(_02592_),
    .Q(\design_top.ROMFF2[4] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14508_ (.D(_02593_),
    .Q(\design_top.ROMFF2[5] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14509_ (.D(_02594_),
    .Q(\design_top.ROMFF2[6] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14510_ (.D(_02595_),
    .Q(\design_top.ROMFF2[7] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14511_ (.D(_02596_),
    .Q(\design_top.ROMFF2[8] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14512_ (.D(_02597_),
    .Q(\design_top.ROMFF2[9] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14513_ (.D(_02598_),
    .Q(\design_top.ROMFF2[10] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14514_ (.D(_02599_),
    .Q(\design_top.ROMFF2[11] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14515_ (.D(_02600_),
    .Q(\design_top.ROMFF2[12] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14516_ (.D(_02601_),
    .Q(\design_top.ROMFF2[13] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14517_ (.D(_02602_),
    .Q(\design_top.ROMFF2[14] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14518_ (.D(_02603_),
    .Q(\design_top.ROMFF2[15] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14519_ (.D(_02604_),
    .Q(\design_top.ROMFF2[16] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14520_ (.D(_02605_),
    .Q(\design_top.ROMFF2[17] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14521_ (.D(_02606_),
    .Q(\design_top.ROMFF2[18] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14522_ (.D(_02607_),
    .Q(\design_top.ROMFF2[19] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14523_ (.D(_02608_),
    .Q(\design_top.ROMFF2[20] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14524_ (.D(_02609_),
    .Q(\design_top.ROMFF2[21] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14525_ (.D(_02610_),
    .Q(\design_top.ROMFF2[22] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14526_ (.D(_02611_),
    .Q(\design_top.ROMFF2[23] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14527_ (.D(_02612_),
    .Q(\design_top.ROMFF2[24] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14528_ (.D(_02613_),
    .Q(\design_top.ROMFF2[25] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14529_ (.D(_02614_),
    .Q(\design_top.ROMFF2[26] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14530_ (.D(_02615_),
    .Q(\design_top.ROMFF2[27] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14531_ (.D(_02616_),
    .Q(\design_top.ROMFF2[28] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14532_ (.D(_02617_),
    .Q(\design_top.ROMFF2[29] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14533_ (.D(_02618_),
    .Q(\design_top.ROMFF2[30] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14534_ (.D(_02619_),
    .Q(\design_top.ROMFF2[31] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14535_ (.D(_02620_),
    .Q(io_out[8]),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14536_ (.D(_02621_),
    .Q(io_out[9]),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14537_ (.D(_02622_),
    .Q(io_out[10]),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14538_ (.D(_02623_),
    .Q(io_out[11]),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14539_ (.D(_02624_),
    .Q(\design_top.LEDFF[4] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14540_ (.D(_02625_),
    .Q(\design_top.LEDFF[5] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14541_ (.D(_02626_),
    .Q(\design_top.LEDFF[6] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14542_ (.D(_02627_),
    .Q(\design_top.LEDFF[7] ),
    .CLK(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14543_ (.D(_02628_),
    .Q(\design_top.LEDFF[8] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14544_ (.D(_02629_),
    .Q(\design_top.LEDFF[9] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14545_ (.D(_02630_),
    .Q(\design_top.LEDFF[10] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14546_ (.D(_02631_),
    .Q(\design_top.LEDFF[11] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14547_ (.D(_02632_),
    .Q(\design_top.LEDFF[12] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14548_ (.D(_02633_),
    .Q(\design_top.LEDFF[13] ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14549_ (.D(_02634_),
    .Q(\design_top.LEDFF[14] ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14550_ (.D(_02635_),
    .Q(\design_top.LEDFF[15] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14551_ (.D(_02636_),
    .Q(io_out[15]),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14552_ (.D(_02637_),
    .Q(\design_top.GPIOFF[1] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14553_ (.D(_02638_),
    .Q(\design_top.GPIOFF[2] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14554_ (.D(_02639_),
    .Q(\design_top.GPIOFF[3] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14555_ (.D(_02640_),
    .Q(\design_top.GPIOFF[4] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14556_ (.D(_02641_),
    .Q(\design_top.GPIOFF[5] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14557_ (.D(_02642_),
    .Q(\design_top.GPIOFF[6] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14558_ (.D(_02643_),
    .Q(\design_top.GPIOFF[7] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14559_ (.D(_02644_),
    .Q(\design_top.GPIOFF[8] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14560_ (.D(_02645_),
    .Q(\design_top.GPIOFF[9] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14561_ (.D(_02646_),
    .Q(\design_top.GPIOFF[10] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14562_ (.D(_02647_),
    .Q(\design_top.GPIOFF[11] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14563_ (.D(_02648_),
    .Q(\design_top.GPIOFF[12] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14564_ (.D(_02649_),
    .Q(\design_top.GPIOFF[13] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14565_ (.D(_02650_),
    .Q(\design_top.GPIOFF[14] ),
    .CLK(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14566_ (.D(_02651_),
    .Q(\design_top.GPIOFF[15] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14567_ (.D(_02652_),
    .Q(\design_top.MEM[9][0] ),
    .CLK(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14568_ (.D(_02653_),
    .Q(\design_top.MEM[9][1] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14569_ (.D(_02654_),
    .Q(\design_top.MEM[9][2] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14570_ (.D(_02655_),
    .Q(\design_top.MEM[9][3] ),
    .CLK(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14571_ (.D(_02656_),
    .Q(\design_top.MEM[9][4] ),
    .CLK(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14572_ (.D(_02657_),
    .Q(\design_top.MEM[9][5] ),
    .CLK(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14573_ (.D(_02658_),
    .Q(\design_top.MEM[9][6] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14574_ (.D(_02659_),
    .Q(\design_top.MEM[9][7] ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14575_ (.D(_02660_),
    .Q(\design_top.MEM[8][0] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14576_ (.D(_02661_),
    .Q(\design_top.MEM[8][1] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14577_ (.D(_02662_),
    .Q(\design_top.MEM[8][2] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14578_ (.D(_02663_),
    .Q(\design_top.MEM[8][3] ),
    .CLK(clknet_leaf_235_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14579_ (.D(_02664_),
    .Q(\design_top.MEM[8][4] ),
    .CLK(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14580_ (.D(_02665_),
    .Q(\design_top.MEM[8][5] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14581_ (.D(_02666_),
    .Q(\design_top.MEM[8][6] ),
    .CLK(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14582_ (.D(_02667_),
    .Q(\design_top.MEM[8][7] ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14583_ (.D(_02668_),
    .Q(\design_top.core0.REG2[14][0] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14584_ (.D(_02669_),
    .Q(\design_top.core0.REG2[14][1] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14585_ (.D(_02670_),
    .Q(\design_top.core0.REG2[14][2] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14586_ (.D(_02671_),
    .Q(\design_top.core0.REG2[14][3] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14587_ (.D(_02672_),
    .Q(\design_top.core0.REG2[14][4] ),
    .CLK(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14588_ (.D(_02673_),
    .Q(\design_top.core0.REG2[14][5] ),
    .CLK(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14589_ (.D(_02674_),
    .Q(\design_top.core0.REG2[14][6] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14590_ (.D(_02675_),
    .Q(\design_top.core0.REG2[14][7] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14591_ (.D(_02676_),
    .Q(\design_top.core0.REG2[14][8] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14592_ (.D(_02677_),
    .Q(\design_top.core0.REG2[14][9] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14593_ (.D(_02678_),
    .Q(\design_top.core0.REG2[14][10] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14594_ (.D(_02679_),
    .Q(\design_top.core0.REG2[14][11] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14595_ (.D(_02680_),
    .Q(\design_top.core0.REG2[14][12] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14596_ (.D(_02681_),
    .Q(\design_top.core0.REG2[14][13] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14597_ (.D(_02682_),
    .Q(\design_top.core0.REG2[14][14] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14598_ (.D(_02683_),
    .Q(\design_top.core0.REG2[14][15] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14599_ (.D(_02684_),
    .Q(\design_top.core0.REG2[14][16] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14600_ (.D(_02685_),
    .Q(\design_top.core0.REG2[14][17] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14601_ (.D(_02686_),
    .Q(\design_top.core0.REG2[14][18] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14602_ (.D(_02687_),
    .Q(\design_top.core0.REG2[14][19] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14603_ (.D(_02688_),
    .Q(\design_top.core0.REG2[14][20] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14604_ (.D(_02689_),
    .Q(\design_top.core0.REG2[14][21] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14605_ (.D(_02690_),
    .Q(\design_top.core0.REG2[14][22] ),
    .CLK(clknet_leaf_76_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14606_ (.D(_02691_),
    .Q(\design_top.core0.REG2[14][23] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14607_ (.D(_02692_),
    .Q(\design_top.core0.REG2[14][24] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14608_ (.D(_02693_),
    .Q(\design_top.core0.REG2[14][25] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14609_ (.D(_02694_),
    .Q(\design_top.core0.REG2[14][26] ),
    .CLK(clknet_leaf_76_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14610_ (.D(_02695_),
    .Q(\design_top.core0.REG2[14][27] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14611_ (.D(_02696_),
    .Q(\design_top.core0.REG2[14][28] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14612_ (.D(_02697_),
    .Q(\design_top.core0.REG2[14][29] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14613_ (.D(_02698_),
    .Q(\design_top.core0.REG2[14][30] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14614_ (.D(_02699_),
    .Q(\design_top.core0.REG2[14][31] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14615_ (.D(_02700_),
    .Q(\design_top.core0.REG2[13][0] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14616_ (.D(_02701_),
    .Q(\design_top.core0.REG2[13][1] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14617_ (.D(_02702_),
    .Q(\design_top.core0.REG2[13][2] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14618_ (.D(_02703_),
    .Q(\design_top.core0.REG2[13][3] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14619_ (.D(_02704_),
    .Q(\design_top.core0.REG2[13][4] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14620_ (.D(_02705_),
    .Q(\design_top.core0.REG2[13][5] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14621_ (.D(_02706_),
    .Q(\design_top.core0.REG2[13][6] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14622_ (.D(_02707_),
    .Q(\design_top.core0.REG2[13][7] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14623_ (.D(_02708_),
    .Q(\design_top.core0.REG2[13][8] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14624_ (.D(_02709_),
    .Q(\design_top.core0.REG2[13][9] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14625_ (.D(_02710_),
    .Q(\design_top.core0.REG2[13][10] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14626_ (.D(_02711_),
    .Q(\design_top.core0.REG2[13][11] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14627_ (.D(_02712_),
    .Q(\design_top.core0.REG2[13][12] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14628_ (.D(_02713_),
    .Q(\design_top.core0.REG2[13][13] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14629_ (.D(_02714_),
    .Q(\design_top.core0.REG2[13][14] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14630_ (.D(_02715_),
    .Q(\design_top.core0.REG2[13][15] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14631_ (.D(_02716_),
    .Q(\design_top.core0.REG2[13][16] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14632_ (.D(_02717_),
    .Q(\design_top.core0.REG2[13][17] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14633_ (.D(_02718_),
    .Q(\design_top.core0.REG2[13][18] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14634_ (.D(_02719_),
    .Q(\design_top.core0.REG2[13][19] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14635_ (.D(_02720_),
    .Q(\design_top.core0.REG2[13][20] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14636_ (.D(_02721_),
    .Q(\design_top.core0.REG2[13][21] ),
    .CLK(clknet_leaf_76_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14637_ (.D(_02722_),
    .Q(\design_top.core0.REG2[13][22] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14638_ (.D(_02723_),
    .Q(\design_top.core0.REG2[13][23] ),
    .CLK(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14639_ (.D(_02724_),
    .Q(\design_top.core0.REG2[13][24] ),
    .CLK(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14640_ (.D(_02725_),
    .Q(\design_top.core0.REG2[13][25] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14641_ (.D(_02726_),
    .Q(\design_top.core0.REG2[13][26] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14642_ (.D(_02727_),
    .Q(\design_top.core0.REG2[13][27] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14643_ (.D(_02728_),
    .Q(\design_top.core0.REG2[13][28] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14644_ (.D(_02729_),
    .Q(\design_top.core0.REG2[13][29] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14645_ (.D(_02730_),
    .Q(\design_top.core0.REG2[13][30] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14646_ (.D(_02731_),
    .Q(\design_top.core0.REG2[13][31] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14647_ (.D(_02732_),
    .Q(\design_top.core0.REG2[12][0] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14648_ (.D(_02733_),
    .Q(\design_top.core0.REG2[12][1] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14649_ (.D(_02734_),
    .Q(\design_top.core0.REG2[12][2] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14650_ (.D(_02735_),
    .Q(\design_top.core0.REG2[12][3] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14651_ (.D(_02736_),
    .Q(\design_top.core0.REG2[12][4] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14652_ (.D(_02737_),
    .Q(\design_top.core0.REG2[12][5] ),
    .CLK(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14653_ (.D(_02738_),
    .Q(\design_top.core0.REG2[12][6] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14654_ (.D(_02739_),
    .Q(\design_top.core0.REG2[12][7] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14655_ (.D(_02740_),
    .Q(\design_top.core0.REG2[12][8] ),
    .CLK(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14656_ (.D(_02741_),
    .Q(\design_top.core0.REG2[12][9] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14657_ (.D(_02742_),
    .Q(\design_top.core0.REG2[12][10] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14658_ (.D(_02743_),
    .Q(\design_top.core0.REG2[12][11] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14659_ (.D(_02744_),
    .Q(\design_top.core0.REG2[12][12] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14660_ (.D(_02745_),
    .Q(\design_top.core0.REG2[12][13] ),
    .CLK(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14661_ (.D(_02746_),
    .Q(\design_top.core0.REG2[12][14] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14662_ (.D(_02747_),
    .Q(\design_top.core0.REG2[12][15] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14663_ (.D(_02748_),
    .Q(\design_top.core0.REG2[12][16] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14664_ (.D(_02749_),
    .Q(\design_top.core0.REG2[12][17] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14665_ (.D(_02750_),
    .Q(\design_top.core0.REG2[12][18] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14666_ (.D(_02751_),
    .Q(\design_top.core0.REG2[12][19] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14667_ (.D(_02752_),
    .Q(\design_top.core0.REG2[12][20] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14668_ (.D(_02753_),
    .Q(\design_top.core0.REG2[12][21] ),
    .CLK(clknet_leaf_76_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14669_ (.D(_02754_),
    .Q(\design_top.core0.REG2[12][22] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14670_ (.D(_02755_),
    .Q(\design_top.core0.REG2[12][23] ),
    .CLK(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14671_ (.D(_02756_),
    .Q(\design_top.core0.REG2[12][24] ),
    .CLK(clknet_leaf_76_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14672_ (.D(_02757_),
    .Q(\design_top.core0.REG2[12][25] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14673_ (.D(_02758_),
    .Q(\design_top.core0.REG2[12][26] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14674_ (.D(_02759_),
    .Q(\design_top.core0.REG2[12][27] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14675_ (.D(_02760_),
    .Q(\design_top.core0.REG2[12][28] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14676_ (.D(_02761_),
    .Q(\design_top.core0.REG2[12][29] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14677_ (.D(_02762_),
    .Q(\design_top.core0.REG2[12][30] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14678_ (.D(_02763_),
    .Q(\design_top.core0.REG2[12][31] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14679_ (.D(_02764_),
    .Q(\design_top.core0.REG2[11][0] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14680_ (.D(_02765_),
    .Q(\design_top.core0.REG2[11][1] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14681_ (.D(_02766_),
    .Q(\design_top.core0.REG2[11][2] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14682_ (.D(_02767_),
    .Q(\design_top.core0.REG2[11][3] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14683_ (.D(_02768_),
    .Q(\design_top.core0.REG2[11][4] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14684_ (.D(_02769_),
    .Q(\design_top.core0.REG2[11][5] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14685_ (.D(_02770_),
    .Q(\design_top.core0.REG2[11][6] ),
    .CLK(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14686_ (.D(_02771_),
    .Q(\design_top.core0.REG2[11][7] ),
    .CLK(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14687_ (.D(_02772_),
    .Q(\design_top.core0.REG2[11][8] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14688_ (.D(_02773_),
    .Q(\design_top.core0.REG2[11][9] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14689_ (.D(_02774_),
    .Q(\design_top.core0.REG2[11][10] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14690_ (.D(_02775_),
    .Q(\design_top.core0.REG2[11][11] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14691_ (.D(_02776_),
    .Q(\design_top.core0.REG2[11][12] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14692_ (.D(_02777_),
    .Q(\design_top.core0.REG2[11][13] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14693_ (.D(_02778_),
    .Q(\design_top.core0.REG2[11][14] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14694_ (.D(_02779_),
    .Q(\design_top.core0.REG2[11][15] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14695_ (.D(_02780_),
    .Q(\design_top.core0.REG2[11][16] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14696_ (.D(_02781_),
    .Q(\design_top.core0.REG2[11][17] ),
    .CLK(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14697_ (.D(_02782_),
    .Q(\design_top.core0.REG2[11][18] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14698_ (.D(_02783_),
    .Q(\design_top.core0.REG2[11][19] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14699_ (.D(_02784_),
    .Q(\design_top.core0.REG2[11][20] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14700_ (.D(_02785_),
    .Q(\design_top.core0.REG2[11][21] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14701_ (.D(_02786_),
    .Q(\design_top.core0.REG2[11][22] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14702_ (.D(_02787_),
    .Q(\design_top.core0.REG2[11][23] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14703_ (.D(_02788_),
    .Q(\design_top.core0.REG2[11][24] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14704_ (.D(_02789_),
    .Q(\design_top.core0.REG2[11][25] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14705_ (.D(_02790_),
    .Q(\design_top.core0.REG2[11][26] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14706_ (.D(_02791_),
    .Q(\design_top.core0.REG2[11][27] ),
    .CLK(clknet_leaf_48_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14707_ (.D(_02792_),
    .Q(\design_top.core0.REG2[11][28] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14708_ (.D(_02793_),
    .Q(\design_top.core0.REG2[11][29] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14709_ (.D(_02794_),
    .Q(\design_top.core0.REG2[11][30] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14710_ (.D(_02795_),
    .Q(\design_top.core0.REG2[11][31] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14711_ (.D(_02796_),
    .Q(\design_top.core0.REG2[10][0] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14712_ (.D(_02797_),
    .Q(\design_top.core0.REG2[10][1] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14713_ (.D(_02798_),
    .Q(\design_top.core0.REG2[10][2] ),
    .CLK(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14714_ (.D(_02799_),
    .Q(\design_top.core0.REG2[10][3] ),
    .CLK(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14715_ (.D(_02800_),
    .Q(\design_top.core0.REG2[10][4] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14716_ (.D(_02801_),
    .Q(\design_top.core0.REG2[10][5] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14717_ (.D(_02802_),
    .Q(\design_top.core0.REG2[10][6] ),
    .CLK(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14718_ (.D(_02803_),
    .Q(\design_top.core0.REG2[10][7] ),
    .CLK(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14719_ (.D(_02804_),
    .Q(\design_top.core0.REG2[10][8] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14720_ (.D(_02805_),
    .Q(\design_top.core0.REG2[10][9] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14721_ (.D(_02806_),
    .Q(\design_top.core0.REG2[10][10] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14722_ (.D(_02807_),
    .Q(\design_top.core0.REG2[10][11] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14723_ (.D(_02808_),
    .Q(\design_top.core0.REG2[10][12] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14724_ (.D(_02809_),
    .Q(\design_top.core0.REG2[10][13] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14725_ (.D(_02810_),
    .Q(\design_top.core0.REG2[10][14] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14726_ (.D(_02811_),
    .Q(\design_top.core0.REG2[10][15] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14727_ (.D(_02812_),
    .Q(\design_top.core0.REG2[10][16] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14728_ (.D(_02813_),
    .Q(\design_top.core0.REG2[10][17] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14729_ (.D(_02814_),
    .Q(\design_top.core0.REG2[10][18] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14730_ (.D(_02815_),
    .Q(\design_top.core0.REG2[10][19] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14731_ (.D(_02816_),
    .Q(\design_top.core0.REG2[10][20] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14732_ (.D(_02817_),
    .Q(\design_top.core0.REG2[10][21] ),
    .CLK(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14733_ (.D(_02818_),
    .Q(\design_top.core0.REG2[10][22] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14734_ (.D(_02819_),
    .Q(\design_top.core0.REG2[10][23] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14735_ (.D(_02820_),
    .Q(\design_top.core0.REG2[10][24] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14736_ (.D(_02821_),
    .Q(\design_top.core0.REG2[10][25] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14737_ (.D(_02822_),
    .Q(\design_top.core0.REG2[10][26] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14738_ (.D(_02823_),
    .Q(\design_top.core0.REG2[10][27] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14739_ (.D(_02824_),
    .Q(\design_top.core0.REG2[10][28] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14740_ (.D(_02825_),
    .Q(\design_top.core0.REG2[10][29] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14741_ (.D(_02826_),
    .Q(\design_top.core0.REG2[10][30] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14742_ (.D(_02827_),
    .Q(\design_top.core0.REG2[10][31] ),
    .CLK(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14743_ (.D(_02828_),
    .Q(\design_top.core0.REG2[0][0] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14744_ (.D(_02829_),
    .Q(\design_top.core0.REG2[0][1] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14745_ (.D(_02830_),
    .Q(\design_top.core0.REG2[0][2] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14746_ (.D(_02831_),
    .Q(\design_top.core0.REG2[0][3] ),
    .CLK(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14747_ (.D(_02832_),
    .Q(\design_top.core0.REG2[0][4] ),
    .CLK(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14748_ (.D(_02833_),
    .Q(\design_top.core0.REG2[0][5] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14749_ (.D(_02834_),
    .Q(\design_top.core0.REG2[0][6] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14750_ (.D(_02835_),
    .Q(\design_top.core0.REG2[0][7] ),
    .CLK(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14751_ (.D(_02836_),
    .Q(\design_top.core0.REG2[0][8] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14752_ (.D(_02837_),
    .Q(\design_top.core0.REG2[0][9] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14753_ (.D(_02838_),
    .Q(\design_top.core0.REG2[0][10] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14754_ (.D(_02839_),
    .Q(\design_top.core0.REG2[0][11] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14755_ (.D(_02840_),
    .Q(\design_top.core0.REG2[0][12] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14756_ (.D(_02841_),
    .Q(\design_top.core0.REG2[0][13] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14757_ (.D(_02842_),
    .Q(\design_top.core0.REG2[0][14] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14758_ (.D(_02843_),
    .Q(\design_top.core0.REG2[0][15] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14759_ (.D(_02844_),
    .Q(\design_top.core0.REG2[0][16] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14760_ (.D(_02845_),
    .Q(\design_top.core0.REG2[0][17] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14761_ (.D(_02846_),
    .Q(\design_top.core0.REG2[0][18] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14762_ (.D(_02847_),
    .Q(\design_top.core0.REG2[0][19] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14763_ (.D(_02848_),
    .Q(\design_top.core0.REG2[0][20] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14764_ (.D(_02849_),
    .Q(\design_top.core0.REG2[0][21] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14765_ (.D(_02850_),
    .Q(\design_top.core0.REG2[0][22] ),
    .CLK(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14766_ (.D(_02851_),
    .Q(\design_top.core0.REG2[0][23] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14767_ (.D(_02852_),
    .Q(\design_top.core0.REG2[0][24] ),
    .CLK(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14768_ (.D(_02853_),
    .Q(\design_top.core0.REG2[0][25] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14769_ (.D(_02854_),
    .Q(\design_top.core0.REG2[0][26] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14770_ (.D(_02855_),
    .Q(\design_top.core0.REG2[0][27] ),
    .CLK(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14771_ (.D(_02856_),
    .Q(\design_top.core0.REG2[0][28] ),
    .CLK(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14772_ (.D(_02857_),
    .Q(\design_top.core0.REG2[0][29] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14773_ (.D(_02858_),
    .Q(\design_top.core0.REG2[0][30] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14774_ (.D(_02859_),
    .Q(\design_top.core0.REG2[0][31] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14775_ (.D(_02860_),
    .Q(\design_top.core0.REG2[8][0] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14776_ (.D(_02861_),
    .Q(\design_top.core0.REG2[8][1] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14777_ (.D(_02862_),
    .Q(\design_top.core0.REG2[8][2] ),
    .CLK(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14778_ (.D(_02863_),
    .Q(\design_top.core0.REG2[8][3] ),
    .CLK(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14779_ (.D(_02864_),
    .Q(\design_top.core0.REG2[8][4] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14780_ (.D(_02865_),
    .Q(\design_top.core0.REG2[8][5] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14781_ (.D(_02866_),
    .Q(\design_top.core0.REG2[8][6] ),
    .CLK(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14782_ (.D(_02867_),
    .Q(\design_top.core0.REG2[8][7] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14783_ (.D(_02868_),
    .Q(\design_top.core0.REG2[8][8] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14784_ (.D(_02869_),
    .Q(\design_top.core0.REG2[8][9] ),
    .CLK(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14785_ (.D(_02870_),
    .Q(\design_top.core0.REG2[8][10] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14786_ (.D(_02871_),
    .Q(\design_top.core0.REG2[8][11] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14787_ (.D(_02872_),
    .Q(\design_top.core0.REG2[8][12] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14788_ (.D(_02873_),
    .Q(\design_top.core0.REG2[8][13] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14789_ (.D(_02874_),
    .Q(\design_top.core0.REG2[8][14] ),
    .CLK(clknet_leaf_37_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14790_ (.D(_02875_),
    .Q(\design_top.core0.REG2[8][15] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14791_ (.D(_02876_),
    .Q(\design_top.core0.REG2[8][16] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14792_ (.D(_02877_),
    .Q(\design_top.core0.REG2[8][17] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14793_ (.D(_02878_),
    .Q(\design_top.core0.REG2[8][18] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14794_ (.D(_02879_),
    .Q(\design_top.core0.REG2[8][19] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14795_ (.D(_02880_),
    .Q(\design_top.core0.REG2[8][20] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14796_ (.D(_02881_),
    .Q(\design_top.core0.REG2[8][21] ),
    .CLK(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14797_ (.D(_02882_),
    .Q(\design_top.core0.REG2[8][22] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14798_ (.D(_02883_),
    .Q(\design_top.core0.REG2[8][23] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14799_ (.D(_02884_),
    .Q(\design_top.core0.REG2[8][24] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14800_ (.D(_02885_),
    .Q(\design_top.core0.REG2[8][25] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14801_ (.D(_02886_),
    .Q(\design_top.core0.REG2[8][26] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14802_ (.D(_02887_),
    .Q(\design_top.core0.REG2[8][27] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14803_ (.D(_02888_),
    .Q(\design_top.core0.REG2[8][28] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14804_ (.D(_02889_),
    .Q(\design_top.core0.REG2[8][29] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14805_ (.D(_02890_),
    .Q(\design_top.core0.REG2[8][30] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14806_ (.D(_02891_),
    .Q(\design_top.core0.REG2[8][31] ),
    .CLK(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14807_ (.D(_02892_),
    .Q(\design_top.core0.REG2[7][0] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14808_ (.D(_02893_),
    .Q(\design_top.core0.REG2[7][1] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14809_ (.D(_02894_),
    .Q(\design_top.core0.REG2[7][2] ),
    .CLK(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14810_ (.D(_02895_),
    .Q(\design_top.core0.REG2[7][3] ),
    .CLK(clknet_leaf_48_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14811_ (.D(_02896_),
    .Q(\design_top.core0.REG2[7][4] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14812_ (.D(_02897_),
    .Q(\design_top.core0.REG2[7][5] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14813_ (.D(_02898_),
    .Q(\design_top.core0.REG2[7][6] ),
    .CLK(clknet_leaf_37_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14814_ (.D(_02899_),
    .Q(\design_top.core0.REG2[7][7] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14815_ (.D(_02900_),
    .Q(\design_top.core0.REG2[7][8] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14816_ (.D(_02901_),
    .Q(\design_top.core0.REG2[7][9] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14817_ (.D(_02902_),
    .Q(\design_top.core0.REG2[7][10] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14818_ (.D(_02903_),
    .Q(\design_top.core0.REG2[7][11] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14819_ (.D(_02904_),
    .Q(\design_top.core0.REG2[7][12] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14820_ (.D(_02905_),
    .Q(\design_top.core0.REG2[7][13] ),
    .CLK(clknet_leaf_79_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14821_ (.D(_02906_),
    .Q(\design_top.core0.REG2[7][14] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14822_ (.D(_02907_),
    .Q(\design_top.core0.REG2[7][15] ),
    .CLK(clknet_leaf_39_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14823_ (.D(_02908_),
    .Q(\design_top.core0.REG2[7][16] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14824_ (.D(_02909_),
    .Q(\design_top.core0.REG2[7][17] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14825_ (.D(_02910_),
    .Q(\design_top.core0.REG2[7][18] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14826_ (.D(_02911_),
    .Q(\design_top.core0.REG2[7][19] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14827_ (.D(_02912_),
    .Q(\design_top.core0.REG2[7][20] ),
    .CLK(clknet_leaf_84_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14828_ (.D(_02913_),
    .Q(\design_top.core0.REG2[7][21] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14829_ (.D(_02914_),
    .Q(\design_top.core0.REG2[7][22] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14830_ (.D(_02915_),
    .Q(\design_top.core0.REG2[7][23] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14831_ (.D(_02916_),
    .Q(\design_top.core0.REG2[7][24] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14832_ (.D(_02917_),
    .Q(\design_top.core0.REG2[7][25] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14833_ (.D(_02918_),
    .Q(\design_top.core0.REG2[7][26] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14834_ (.D(_02919_),
    .Q(\design_top.core0.REG2[7][27] ),
    .CLK(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14835_ (.D(_02920_),
    .Q(\design_top.core0.REG2[7][28] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14836_ (.D(_02921_),
    .Q(\design_top.core0.REG2[7][29] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14837_ (.D(_02922_),
    .Q(\design_top.core0.REG2[7][30] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14838_ (.D(_02923_),
    .Q(\design_top.core0.REG2[7][31] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14839_ (.D(_02924_),
    .Q(\design_top.core0.REG2[6][0] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14840_ (.D(_02925_),
    .Q(\design_top.core0.REG2[6][1] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14841_ (.D(_02926_),
    .Q(\design_top.core0.REG2[6][2] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14842_ (.D(_02927_),
    .Q(\design_top.core0.REG2[6][3] ),
    .CLK(clknet_leaf_48_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14843_ (.D(_02928_),
    .Q(\design_top.core0.REG2[6][4] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14844_ (.D(_02929_),
    .Q(\design_top.core0.REG2[6][5] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14845_ (.D(_02930_),
    .Q(\design_top.core0.REG2[6][6] ),
    .CLK(clknet_leaf_37_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14846_ (.D(_02931_),
    .Q(\design_top.core0.REG2[6][7] ),
    .CLK(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14847_ (.D(_02932_),
    .Q(\design_top.core0.REG2[6][8] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14848_ (.D(_02933_),
    .Q(\design_top.core0.REG2[6][9] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14849_ (.D(_02934_),
    .Q(\design_top.core0.REG2[6][10] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14850_ (.D(_02935_),
    .Q(\design_top.core0.REG2[6][11] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14851_ (.D(_02936_),
    .Q(\design_top.core0.REG2[6][12] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14852_ (.D(_02937_),
    .Q(\design_top.core0.REG2[6][13] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14853_ (.D(_02938_),
    .Q(\design_top.core0.REG2[6][14] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14854_ (.D(_02939_),
    .Q(\design_top.core0.REG2[6][15] ),
    .CLK(clknet_leaf_39_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14855_ (.D(_02940_),
    .Q(\design_top.core0.REG2[6][16] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14856_ (.D(_02941_),
    .Q(\design_top.core0.REG2[6][17] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14857_ (.D(_02942_),
    .Q(\design_top.core0.REG2[6][18] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14858_ (.D(_02943_),
    .Q(\design_top.core0.REG2[6][19] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14859_ (.D(_02944_),
    .Q(\design_top.core0.REG2[6][20] ),
    .CLK(clknet_leaf_84_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14860_ (.D(_02945_),
    .Q(\design_top.core0.REG2[6][21] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14861_ (.D(_02946_),
    .Q(\design_top.core0.REG2[6][22] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14862_ (.D(_02947_),
    .Q(\design_top.core0.REG2[6][23] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14863_ (.D(_02948_),
    .Q(\design_top.core0.REG2[6][24] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14864_ (.D(_02949_),
    .Q(\design_top.core0.REG2[6][25] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14865_ (.D(_02950_),
    .Q(\design_top.core0.REG2[6][26] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14866_ (.D(_02951_),
    .Q(\design_top.core0.REG2[6][27] ),
    .CLK(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14867_ (.D(_02952_),
    .Q(\design_top.core0.REG2[6][28] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14868_ (.D(_02953_),
    .Q(\design_top.core0.REG2[6][29] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14869_ (.D(_02954_),
    .Q(\design_top.core0.REG2[6][30] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14870_ (.D(_02955_),
    .Q(\design_top.core0.REG2[6][31] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14871_ (.D(_02956_),
    .Q(\design_top.core0.REG2[5][0] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14872_ (.D(_02957_),
    .Q(\design_top.core0.REG2[5][1] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14873_ (.D(_02958_),
    .Q(\design_top.core0.REG2[5][2] ),
    .CLK(clknet_leaf_48_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14874_ (.D(_02959_),
    .Q(\design_top.core0.REG2[5][3] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14875_ (.D(_02960_),
    .Q(\design_top.core0.REG2[5][4] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14876_ (.D(_02961_),
    .Q(\design_top.core0.REG2[5][5] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14877_ (.D(_02962_),
    .Q(\design_top.core0.REG2[5][6] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14878_ (.D(_02963_),
    .Q(\design_top.core0.REG2[5][7] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14879_ (.D(_02964_),
    .Q(\design_top.core0.REG2[5][8] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14880_ (.D(_02965_),
    .Q(\design_top.core0.REG2[5][9] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14881_ (.D(_02966_),
    .Q(\design_top.core0.REG2[5][10] ),
    .CLK(clknet_leaf_37_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14882_ (.D(_02967_),
    .Q(\design_top.core0.REG2[5][11] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14883_ (.D(_02968_),
    .Q(\design_top.core0.REG2[5][12] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14884_ (.D(_02969_),
    .Q(\design_top.core0.REG2[5][13] ),
    .CLK(clknet_leaf_79_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14885_ (.D(_02970_),
    .Q(\design_top.core0.REG2[5][14] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14886_ (.D(_02971_),
    .Q(\design_top.core0.REG2[5][15] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14887_ (.D(_02972_),
    .Q(\design_top.core0.REG2[5][16] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14888_ (.D(_02973_),
    .Q(\design_top.core0.REG2[5][17] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14889_ (.D(_02974_),
    .Q(\design_top.core0.REG2[5][18] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14890_ (.D(_02975_),
    .Q(\design_top.core0.REG2[5][19] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14891_ (.D(_02976_),
    .Q(\design_top.core0.REG2[5][20] ),
    .CLK(clknet_leaf_84_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14892_ (.D(_02977_),
    .Q(\design_top.core0.REG2[5][21] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14893_ (.D(_02978_),
    .Q(\design_top.core0.REG2[5][22] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14894_ (.D(_02979_),
    .Q(\design_top.core0.REG2[5][23] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14895_ (.D(_02980_),
    .Q(\design_top.core0.REG2[5][24] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14896_ (.D(_02981_),
    .Q(\design_top.core0.REG2[5][25] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14897_ (.D(_02982_),
    .Q(\design_top.core0.REG2[5][26] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14898_ (.D(_02983_),
    .Q(\design_top.core0.REG2[5][27] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14899_ (.D(_02984_),
    .Q(\design_top.core0.REG2[5][28] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14900_ (.D(_02985_),
    .Q(\design_top.core0.REG2[5][29] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14901_ (.D(_02986_),
    .Q(\design_top.core0.REG2[5][30] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14902_ (.D(_02987_),
    .Q(\design_top.core0.REG2[5][31] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14903_ (.D(_02988_),
    .Q(\design_top.MEM[7][0] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14904_ (.D(_02989_),
    .Q(\design_top.MEM[7][1] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14905_ (.D(_02990_),
    .Q(\design_top.MEM[7][2] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14906_ (.D(_02991_),
    .Q(\design_top.MEM[7][3] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14907_ (.D(_02992_),
    .Q(\design_top.MEM[7][4] ),
    .CLK(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14908_ (.D(_02993_),
    .Q(\design_top.MEM[7][5] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14909_ (.D(_02994_),
    .Q(\design_top.MEM[7][6] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14910_ (.D(_02995_),
    .Q(\design_top.MEM[7][7] ),
    .CLK(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14911_ (.D(_02996_),
    .Q(\design_top.core0.REG2[4][0] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14912_ (.D(_02997_),
    .Q(\design_top.core0.REG2[4][1] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14913_ (.D(_02998_),
    .Q(\design_top.core0.REG2[4][2] ),
    .CLK(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14914_ (.D(_02999_),
    .Q(\design_top.core0.REG2[4][3] ),
    .CLK(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14915_ (.D(_03000_),
    .Q(\design_top.core0.REG2[4][4] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14916_ (.D(_03001_),
    .Q(\design_top.core0.REG2[4][5] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14917_ (.D(_03002_),
    .Q(\design_top.core0.REG2[4][6] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14918_ (.D(_03003_),
    .Q(\design_top.core0.REG2[4][7] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14919_ (.D(_03004_),
    .Q(\design_top.core0.REG2[4][8] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14920_ (.D(_03005_),
    .Q(\design_top.core0.REG2[4][9] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14921_ (.D(_03006_),
    .Q(\design_top.core0.REG2[4][10] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14922_ (.D(_03007_),
    .Q(\design_top.core0.REG2[4][11] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14923_ (.D(_03008_),
    .Q(\design_top.core0.REG2[4][12] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14924_ (.D(_03009_),
    .Q(\design_top.core0.REG2[4][13] ),
    .CLK(clknet_leaf_79_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14925_ (.D(_03010_),
    .Q(\design_top.core0.REG2[4][14] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14926_ (.D(_03011_),
    .Q(\design_top.core0.REG2[4][15] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14927_ (.D(_03012_),
    .Q(\design_top.core0.REG2[4][16] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14928_ (.D(_03013_),
    .Q(\design_top.core0.REG2[4][17] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14929_ (.D(_03014_),
    .Q(\design_top.core0.REG2[4][18] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14930_ (.D(_03015_),
    .Q(\design_top.core0.REG2[4][19] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14931_ (.D(_03016_),
    .Q(\design_top.core0.REG2[4][20] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14932_ (.D(_03017_),
    .Q(\design_top.core0.REG2[4][21] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14933_ (.D(_03018_),
    .Q(\design_top.core0.REG2[4][22] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14934_ (.D(_03019_),
    .Q(\design_top.core0.REG2[4][23] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14935_ (.D(_03020_),
    .Q(\design_top.core0.REG2[4][24] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14936_ (.D(_03021_),
    .Q(\design_top.core0.REG2[4][25] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14937_ (.D(_03022_),
    .Q(\design_top.core0.REG2[4][26] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14938_ (.D(_03023_),
    .Q(\design_top.core0.REG2[4][27] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14939_ (.D(_03024_),
    .Q(\design_top.core0.REG2[4][28] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14940_ (.D(_03025_),
    .Q(\design_top.core0.REG2[4][29] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14941_ (.D(_03026_),
    .Q(\design_top.core0.REG2[4][30] ),
    .CLK(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14942_ (.D(_03027_),
    .Q(\design_top.core0.REG2[4][31] ),
    .CLK(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14943_ (.D(_03028_),
    .Q(\design_top.core0.REG2[3][0] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14944_ (.D(_03029_),
    .Q(\design_top.core0.REG2[3][1] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14945_ (.D(_03030_),
    .Q(\design_top.core0.REG2[3][2] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14946_ (.D(_03031_),
    .Q(\design_top.core0.REG2[3][3] ),
    .CLK(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14947_ (.D(_03032_),
    .Q(\design_top.core0.REG2[3][4] ),
    .CLK(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14948_ (.D(_03033_),
    .Q(\design_top.core0.REG2[3][5] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14949_ (.D(_03034_),
    .Q(\design_top.core0.REG2[3][6] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14950_ (.D(_03035_),
    .Q(\design_top.core0.REG2[3][7] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14951_ (.D(_03036_),
    .Q(\design_top.core0.REG2[3][8] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14952_ (.D(_03037_),
    .Q(\design_top.core0.REG2[3][9] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14953_ (.D(_03038_),
    .Q(\design_top.core0.REG2[3][10] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14954_ (.D(_03039_),
    .Q(\design_top.core0.REG2[3][11] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14955_ (.D(_03040_),
    .Q(\design_top.core0.REG2[3][12] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14956_ (.D(_03041_),
    .Q(\design_top.core0.REG2[3][13] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14957_ (.D(_03042_),
    .Q(\design_top.core0.REG2[3][14] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14958_ (.D(_03043_),
    .Q(\design_top.core0.REG2[3][15] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14959_ (.D(_03044_),
    .Q(\design_top.core0.REG2[3][16] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14960_ (.D(_03045_),
    .Q(\design_top.core0.REG2[3][17] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14961_ (.D(_03046_),
    .Q(\design_top.core0.REG2[3][18] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14962_ (.D(_03047_),
    .Q(\design_top.core0.REG2[3][19] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14963_ (.D(_03048_),
    .Q(\design_top.core0.REG2[3][20] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14964_ (.D(_03049_),
    .Q(\design_top.core0.REG2[3][21] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14965_ (.D(_03050_),
    .Q(\design_top.core0.REG2[3][22] ),
    .CLK(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14966_ (.D(_03051_),
    .Q(\design_top.core0.REG2[3][23] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14967_ (.D(_03052_),
    .Q(\design_top.core0.REG2[3][24] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14968_ (.D(_03053_),
    .Q(\design_top.core0.REG2[3][25] ),
    .CLK(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14969_ (.D(_03054_),
    .Q(\design_top.core0.REG2[3][26] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14970_ (.D(_03055_),
    .Q(\design_top.core0.REG2[3][27] ),
    .CLK(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14971_ (.D(_03056_),
    .Q(\design_top.core0.REG2[3][28] ),
    .CLK(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14972_ (.D(_03057_),
    .Q(\design_top.core0.REG2[3][29] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14973_ (.D(_03058_),
    .Q(\design_top.core0.REG2[3][30] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14974_ (.D(_03059_),
    .Q(\design_top.core0.REG2[3][31] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14975_ (.D(_03060_),
    .Q(\design_top.core0.REG2[2][0] ),
    .CLK(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14976_ (.D(_03061_),
    .Q(\design_top.core0.REG2[2][1] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14977_ (.D(_03062_),
    .Q(\design_top.core0.REG2[2][2] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14978_ (.D(_03063_),
    .Q(\design_top.core0.REG2[2][3] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14979_ (.D(_03064_),
    .Q(\design_top.core0.REG2[2][4] ),
    .CLK(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14980_ (.D(_03065_),
    .Q(\design_top.core0.REG2[2][5] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14981_ (.D(_03066_),
    .Q(\design_top.core0.REG2[2][6] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14982_ (.D(_03067_),
    .Q(\design_top.core0.REG2[2][7] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14983_ (.D(_03068_),
    .Q(\design_top.core0.REG2[2][8] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14984_ (.D(_03069_),
    .Q(\design_top.core0.REG2[2][9] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14985_ (.D(_03070_),
    .Q(\design_top.core0.REG2[2][10] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14986_ (.D(_03071_),
    .Q(\design_top.core0.REG2[2][11] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14987_ (.D(_03072_),
    .Q(\design_top.core0.REG2[2][12] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14988_ (.D(_03073_),
    .Q(\design_top.core0.REG2[2][13] ),
    .CLK(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14989_ (.D(_03074_),
    .Q(\design_top.core0.REG2[2][14] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14990_ (.D(_03075_),
    .Q(\design_top.core0.REG2[2][15] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14991_ (.D(_03076_),
    .Q(\design_top.core0.REG2[2][16] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14992_ (.D(_03077_),
    .Q(\design_top.core0.REG2[2][17] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14993_ (.D(_03078_),
    .Q(\design_top.core0.REG2[2][18] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14994_ (.D(_03079_),
    .Q(\design_top.core0.REG2[2][19] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14995_ (.D(_03080_),
    .Q(\design_top.core0.REG2[2][20] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14996_ (.D(_03081_),
    .Q(\design_top.core0.REG2[2][21] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14997_ (.D(_03082_),
    .Q(\design_top.core0.REG2[2][22] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14998_ (.D(_03083_),
    .Q(\design_top.core0.REG2[2][23] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _14999_ (.D(_03084_),
    .Q(\design_top.core0.REG2[2][24] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15000_ (.D(_03085_),
    .Q(\design_top.core0.REG2[2][25] ),
    .CLK(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15001_ (.D(_03086_),
    .Q(\design_top.core0.REG2[2][26] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15002_ (.D(_03087_),
    .Q(\design_top.core0.REG2[2][27] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15003_ (.D(_03088_),
    .Q(\design_top.core0.REG2[2][28] ),
    .CLK(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15004_ (.D(_03089_),
    .Q(\design_top.core0.REG2[2][29] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15005_ (.D(_03090_),
    .Q(\design_top.core0.REG2[2][30] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15006_ (.D(_03091_),
    .Q(\design_top.core0.REG2[2][31] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15007_ (.D(_03092_),
    .Q(\design_top.core0.REG2[1][0] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15008_ (.D(_03093_),
    .Q(\design_top.core0.REG2[1][1] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15009_ (.D(_03094_),
    .Q(\design_top.core0.REG2[1][2] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15010_ (.D(_03095_),
    .Q(\design_top.core0.REG2[1][3] ),
    .CLK(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15011_ (.D(_03096_),
    .Q(\design_top.core0.REG2[1][4] ),
    .CLK(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15012_ (.D(_03097_),
    .Q(\design_top.core0.REG2[1][5] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15013_ (.D(_03098_),
    .Q(\design_top.core0.REG2[1][6] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15014_ (.D(_03099_),
    .Q(\design_top.core0.REG2[1][7] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15015_ (.D(_03100_),
    .Q(\design_top.core0.REG2[1][8] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15016_ (.D(_03101_),
    .Q(\design_top.core0.REG2[1][9] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15017_ (.D(_03102_),
    .Q(\design_top.core0.REG2[1][10] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15018_ (.D(_03103_),
    .Q(\design_top.core0.REG2[1][11] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15019_ (.D(_03104_),
    .Q(\design_top.core0.REG2[1][12] ),
    .CLK(clknet_leaf_79_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15020_ (.D(_03105_),
    .Q(\design_top.core0.REG2[1][13] ),
    .CLK(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15021_ (.D(_03106_),
    .Q(\design_top.core0.REG2[1][14] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15022_ (.D(_03107_),
    .Q(\design_top.core0.REG2[1][15] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15023_ (.D(_03108_),
    .Q(\design_top.core0.REG2[1][16] ),
    .CLK(clknet_leaf_79_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15024_ (.D(_03109_),
    .Q(\design_top.core0.REG2[1][17] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15025_ (.D(_03110_),
    .Q(\design_top.core0.REG2[1][18] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15026_ (.D(_03111_),
    .Q(\design_top.core0.REG2[1][19] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15027_ (.D(_03112_),
    .Q(\design_top.core0.REG2[1][20] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15028_ (.D(_03113_),
    .Q(\design_top.core0.REG2[1][21] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15029_ (.D(_03114_),
    .Q(\design_top.core0.REG2[1][22] ),
    .CLK(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15030_ (.D(_03115_),
    .Q(\design_top.core0.REG2[1][23] ),
    .CLK(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15031_ (.D(_03116_),
    .Q(\design_top.core0.REG2[1][24] ),
    .CLK(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15032_ (.D(_03117_),
    .Q(\design_top.core0.REG2[1][25] ),
    .CLK(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15033_ (.D(_03118_),
    .Q(\design_top.core0.REG2[1][26] ),
    .CLK(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15034_ (.D(_03119_),
    .Q(\design_top.core0.REG2[1][27] ),
    .CLK(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15035_ (.D(_03120_),
    .Q(\design_top.core0.REG2[1][28] ),
    .CLK(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15036_ (.D(_03121_),
    .Q(\design_top.core0.REG2[1][29] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15037_ (.D(_03122_),
    .Q(\design_top.core0.REG2[1][30] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15038_ (.D(_03123_),
    .Q(\design_top.core0.REG2[1][31] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15039_ (.D(_03124_),
    .Q(\design_top.core0.REG2[15][0] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15040_ (.D(_03125_),
    .Q(\design_top.core0.REG2[15][1] ),
    .CLK(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15041_ (.D(_03126_),
    .Q(\design_top.core0.REG2[15][2] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15042_ (.D(_03127_),
    .Q(\design_top.core0.REG2[15][3] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15043_ (.D(_03128_),
    .Q(\design_top.core0.REG2[15][4] ),
    .CLK(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15044_ (.D(_03129_),
    .Q(\design_top.core0.REG2[15][5] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15045_ (.D(_03130_),
    .Q(\design_top.core0.REG2[15][6] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15046_ (.D(_03131_),
    .Q(\design_top.core0.REG2[15][7] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15047_ (.D(_03132_),
    .Q(\design_top.core0.REG2[15][8] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15048_ (.D(_03133_),
    .Q(\design_top.core0.REG2[15][9] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15049_ (.D(_03134_),
    .Q(\design_top.core0.REG2[15][10] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15050_ (.D(_03135_),
    .Q(\design_top.core0.REG2[15][11] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15051_ (.D(_03136_),
    .Q(\design_top.core0.REG2[15][12] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15052_ (.D(_03137_),
    .Q(\design_top.core0.REG2[15][13] ),
    .CLK(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15053_ (.D(_03138_),
    .Q(\design_top.core0.REG2[15][14] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15054_ (.D(_03139_),
    .Q(\design_top.core0.REG2[15][15] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15055_ (.D(_03140_),
    .Q(\design_top.core0.REG2[15][16] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15056_ (.D(_03141_),
    .Q(\design_top.core0.REG2[15][17] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15057_ (.D(_03142_),
    .Q(\design_top.core0.REG2[15][18] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15058_ (.D(_03143_),
    .Q(\design_top.core0.REG2[15][19] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15059_ (.D(_03144_),
    .Q(\design_top.core0.REG2[15][20] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15060_ (.D(_03145_),
    .Q(\design_top.core0.REG2[15][21] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15061_ (.D(_03146_),
    .Q(\design_top.core0.REG2[15][22] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15062_ (.D(_03147_),
    .Q(\design_top.core0.REG2[15][23] ),
    .CLK(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15063_ (.D(_03148_),
    .Q(\design_top.core0.REG2[15][24] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15064_ (.D(_03149_),
    .Q(\design_top.core0.REG2[15][25] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15065_ (.D(_03150_),
    .Q(\design_top.core0.REG2[15][26] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15066_ (.D(_03151_),
    .Q(\design_top.core0.REG2[15][27] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15067_ (.D(_03152_),
    .Q(\design_top.core0.REG2[15][28] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15068_ (.D(_03153_),
    .Q(\design_top.core0.REG2[15][29] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15069_ (.D(_03154_),
    .Q(\design_top.core0.REG2[15][30] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15070_ (.D(_03155_),
    .Q(\design_top.core0.REG2[15][31] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15071_ (.D(_03156_),
    .Q(\design_top.MEM[6][0] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15072_ (.D(_03157_),
    .Q(\design_top.MEM[6][1] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15073_ (.D(_03158_),
    .Q(\design_top.MEM[6][2] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15074_ (.D(_03159_),
    .Q(\design_top.MEM[6][3] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15075_ (.D(_03160_),
    .Q(\design_top.MEM[6][4] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15076_ (.D(_03161_),
    .Q(\design_top.MEM[6][5] ),
    .CLK(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15077_ (.D(_03162_),
    .Q(\design_top.MEM[6][6] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15078_ (.D(_03163_),
    .Q(\design_top.MEM[6][7] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15079_ (.D(_03164_),
    .Q(\design_top.MEM[5][0] ),
    .CLK(clknet_leaf_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15080_ (.D(_03165_),
    .Q(\design_top.MEM[5][1] ),
    .CLK(clknet_leaf_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15081_ (.D(_03166_),
    .Q(\design_top.MEM[5][2] ),
    .CLK(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15082_ (.D(_03167_),
    .Q(\design_top.MEM[5][3] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15083_ (.D(_03168_),
    .Q(\design_top.MEM[5][4] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15084_ (.D(_03169_),
    .Q(\design_top.MEM[5][5] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15085_ (.D(_03170_),
    .Q(\design_top.MEM[5][6] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15086_ (.D(_03171_),
    .Q(\design_top.MEM[5][7] ),
    .CLK(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15087_ (.D(_03172_),
    .Q(\design_top.core0.REG1[14][0] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15088_ (.D(_03173_),
    .Q(\design_top.core0.REG1[14][1] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15089_ (.D(_03174_),
    .Q(\design_top.core0.REG1[14][2] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15090_ (.D(_03175_),
    .Q(\design_top.core0.REG1[14][3] ),
    .CLK(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15091_ (.D(_03176_),
    .Q(\design_top.core0.REG1[14][4] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15092_ (.D(_03177_),
    .Q(\design_top.core0.REG1[14][5] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15093_ (.D(_03178_),
    .Q(\design_top.core0.REG1[14][6] ),
    .CLK(clknet_leaf_143_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15094_ (.D(_03179_),
    .Q(\design_top.core0.REG1[14][7] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15095_ (.D(_03180_),
    .Q(\design_top.core0.REG1[14][8] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15096_ (.D(_03181_),
    .Q(\design_top.core0.REG1[14][9] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15097_ (.D(_03182_),
    .Q(\design_top.core0.REG1[14][10] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15098_ (.D(_03183_),
    .Q(\design_top.core0.REG1[14][11] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15099_ (.D(_03184_),
    .Q(\design_top.core0.REG1[14][12] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15100_ (.D(_03185_),
    .Q(\design_top.core0.REG1[14][13] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15101_ (.D(_03186_),
    .Q(\design_top.core0.REG1[14][14] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15102_ (.D(_03187_),
    .Q(\design_top.core0.REG1[14][15] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15103_ (.D(_03188_),
    .Q(\design_top.core0.REG1[14][16] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15104_ (.D(_03189_),
    .Q(\design_top.core0.REG1[14][17] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15105_ (.D(_03190_),
    .Q(\design_top.core0.REG1[14][18] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15106_ (.D(_03191_),
    .Q(\design_top.core0.REG1[14][19] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15107_ (.D(_03192_),
    .Q(\design_top.core0.REG1[14][20] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15108_ (.D(_03193_),
    .Q(\design_top.core0.REG1[14][21] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15109_ (.D(_03194_),
    .Q(\design_top.core0.REG1[14][22] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15110_ (.D(_03195_),
    .Q(\design_top.core0.REG1[14][23] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15111_ (.D(_03196_),
    .Q(\design_top.core0.REG1[14][24] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15112_ (.D(_03197_),
    .Q(\design_top.core0.REG1[14][25] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15113_ (.D(_03198_),
    .Q(\design_top.core0.REG1[14][26] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15114_ (.D(_03199_),
    .Q(\design_top.core0.REG1[14][27] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15115_ (.D(_03200_),
    .Q(\design_top.core0.REG1[14][28] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15116_ (.D(_03201_),
    .Q(\design_top.core0.REG1[14][29] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15117_ (.D(_03202_),
    .Q(\design_top.core0.REG1[14][30] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15118_ (.D(_03203_),
    .Q(\design_top.core0.REG1[14][31] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15119_ (.D(_03204_),
    .Q(\design_top.core0.REG1[13][0] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15120_ (.D(_03205_),
    .Q(\design_top.core0.REG1[13][1] ),
    .CLK(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15121_ (.D(_03206_),
    .Q(\design_top.core0.REG1[13][2] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15122_ (.D(_03207_),
    .Q(\design_top.core0.REG1[13][3] ),
    .CLK(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15123_ (.D(_03208_),
    .Q(\design_top.core0.REG1[13][4] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15124_ (.D(_03209_),
    .Q(\design_top.core0.REG1[13][5] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15125_ (.D(_03210_),
    .Q(\design_top.core0.REG1[13][6] ),
    .CLK(clknet_leaf_143_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15126_ (.D(_03211_),
    .Q(\design_top.core0.REG1[13][7] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15127_ (.D(_03212_),
    .Q(\design_top.core0.REG1[13][8] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15128_ (.D(_03213_),
    .Q(\design_top.core0.REG1[13][9] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15129_ (.D(_03214_),
    .Q(\design_top.core0.REG1[13][10] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15130_ (.D(_03215_),
    .Q(\design_top.core0.REG1[13][11] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15131_ (.D(_03216_),
    .Q(\design_top.core0.REG1[13][12] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15132_ (.D(_03217_),
    .Q(\design_top.core0.REG1[13][13] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15133_ (.D(_03218_),
    .Q(\design_top.core0.REG1[13][14] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15134_ (.D(_03219_),
    .Q(\design_top.core0.REG1[13][15] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15135_ (.D(_03220_),
    .Q(\design_top.core0.REG1[13][16] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15136_ (.D(_03221_),
    .Q(\design_top.core0.REG1[13][17] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15137_ (.D(_03222_),
    .Q(\design_top.core0.REG1[13][18] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15138_ (.D(_03223_),
    .Q(\design_top.core0.REG1[13][19] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15139_ (.D(_03224_),
    .Q(\design_top.core0.REG1[13][20] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15140_ (.D(_03225_),
    .Q(\design_top.core0.REG1[13][21] ),
    .CLK(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15141_ (.D(_03226_),
    .Q(\design_top.core0.REG1[13][22] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15142_ (.D(_03227_),
    .Q(\design_top.core0.REG1[13][23] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15143_ (.D(_03228_),
    .Q(\design_top.core0.REG1[13][24] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15144_ (.D(_03229_),
    .Q(\design_top.core0.REG1[13][25] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15145_ (.D(_03230_),
    .Q(\design_top.core0.REG1[13][26] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15146_ (.D(_03231_),
    .Q(\design_top.core0.REG1[13][27] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15147_ (.D(_03232_),
    .Q(\design_top.core0.REG1[13][28] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15148_ (.D(_03233_),
    .Q(\design_top.core0.REG1[13][29] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15149_ (.D(_03234_),
    .Q(\design_top.core0.REG1[13][30] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15150_ (.D(_03235_),
    .Q(\design_top.core0.REG1[13][31] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15151_ (.D(_03236_),
    .Q(\design_top.core0.REG1[12][0] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15152_ (.D(_03237_),
    .Q(\design_top.core0.REG1[12][1] ),
    .CLK(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15153_ (.D(_03238_),
    .Q(\design_top.core0.REG1[12][2] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15154_ (.D(_03239_),
    .Q(\design_top.core0.REG1[12][3] ),
    .CLK(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15155_ (.D(_03240_),
    .Q(\design_top.core0.REG1[12][4] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15156_ (.D(_03241_),
    .Q(\design_top.core0.REG1[12][5] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15157_ (.D(_03242_),
    .Q(\design_top.core0.REG1[12][6] ),
    .CLK(clknet_leaf_143_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15158_ (.D(_03243_),
    .Q(\design_top.core0.REG1[12][7] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15159_ (.D(_03244_),
    .Q(\design_top.core0.REG1[12][8] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15160_ (.D(_03245_),
    .Q(\design_top.core0.REG1[12][9] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15161_ (.D(_03246_),
    .Q(\design_top.core0.REG1[12][10] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15162_ (.D(_03247_),
    .Q(\design_top.core0.REG1[12][11] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15163_ (.D(_03248_),
    .Q(\design_top.core0.REG1[12][12] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15164_ (.D(_03249_),
    .Q(\design_top.core0.REG1[12][13] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15165_ (.D(_03250_),
    .Q(\design_top.core0.REG1[12][14] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15166_ (.D(_03251_),
    .Q(\design_top.core0.REG1[12][15] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15167_ (.D(_03252_),
    .Q(\design_top.core0.REG1[12][16] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15168_ (.D(_03253_),
    .Q(\design_top.core0.REG1[12][17] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15169_ (.D(_03254_),
    .Q(\design_top.core0.REG1[12][18] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15170_ (.D(_03255_),
    .Q(\design_top.core0.REG1[12][19] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15171_ (.D(_03256_),
    .Q(\design_top.core0.REG1[12][20] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15172_ (.D(_03257_),
    .Q(\design_top.core0.REG1[12][21] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15173_ (.D(_03258_),
    .Q(\design_top.core0.REG1[12][22] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15174_ (.D(_03259_),
    .Q(\design_top.core0.REG1[12][23] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15175_ (.D(_03260_),
    .Q(\design_top.core0.REG1[12][24] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15176_ (.D(_03261_),
    .Q(\design_top.core0.REG1[12][25] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15177_ (.D(_03262_),
    .Q(\design_top.core0.REG1[12][26] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15178_ (.D(_03263_),
    .Q(\design_top.core0.REG1[12][27] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15179_ (.D(_03264_),
    .Q(\design_top.core0.REG1[12][28] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15180_ (.D(_03265_),
    .Q(\design_top.core0.REG1[12][29] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15181_ (.D(_03266_),
    .Q(\design_top.core0.REG1[12][30] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15182_ (.D(_03267_),
    .Q(\design_top.core0.REG1[12][31] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15183_ (.D(_03268_),
    .Q(\design_top.core0.REG1[11][0] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15184_ (.D(_03269_),
    .Q(\design_top.core0.REG1[11][1] ),
    .CLK(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15185_ (.D(_03270_),
    .Q(\design_top.core0.REG1[11][2] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15186_ (.D(_03271_),
    .Q(\design_top.core0.REG1[11][3] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15187_ (.D(_03272_),
    .Q(\design_top.core0.REG1[11][4] ),
    .CLK(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15188_ (.D(_03273_),
    .Q(\design_top.core0.REG1[11][5] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15189_ (.D(_03274_),
    .Q(\design_top.core0.REG1[11][6] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15190_ (.D(_03275_),
    .Q(\design_top.core0.REG1[11][7] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15191_ (.D(_03276_),
    .Q(\design_top.core0.REG1[11][8] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15192_ (.D(_03277_),
    .Q(\design_top.core0.REG1[11][9] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15193_ (.D(_03278_),
    .Q(\design_top.core0.REG1[11][10] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15194_ (.D(_03279_),
    .Q(\design_top.core0.REG1[11][11] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15195_ (.D(_03280_),
    .Q(\design_top.core0.REG1[11][12] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15196_ (.D(_03281_),
    .Q(\design_top.core0.REG1[11][13] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15197_ (.D(_03282_),
    .Q(\design_top.core0.REG1[11][14] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15198_ (.D(_03283_),
    .Q(\design_top.core0.REG1[11][15] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15199_ (.D(_03284_),
    .Q(\design_top.core0.REG1[11][16] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15200_ (.D(_03285_),
    .Q(\design_top.core0.REG1[11][17] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15201_ (.D(_03286_),
    .Q(\design_top.core0.REG1[11][18] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15202_ (.D(_03287_),
    .Q(\design_top.core0.REG1[11][19] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15203_ (.D(_03288_),
    .Q(\design_top.core0.REG1[11][20] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15204_ (.D(_03289_),
    .Q(\design_top.core0.REG1[11][21] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15205_ (.D(_03290_),
    .Q(\design_top.core0.REG1[11][22] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15206_ (.D(_03291_),
    .Q(\design_top.core0.REG1[11][23] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15207_ (.D(_03292_),
    .Q(\design_top.core0.REG1[11][24] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15208_ (.D(_03293_),
    .Q(\design_top.core0.REG1[11][25] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15209_ (.D(_03294_),
    .Q(\design_top.core0.REG1[11][26] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15210_ (.D(_03295_),
    .Q(\design_top.core0.REG1[11][27] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15211_ (.D(_03296_),
    .Q(\design_top.core0.REG1[11][28] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15212_ (.D(_03297_),
    .Q(\design_top.core0.REG1[11][29] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15213_ (.D(_03298_),
    .Q(\design_top.core0.REG1[11][30] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15214_ (.D(_03299_),
    .Q(\design_top.core0.REG1[11][31] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15215_ (.D(_03300_),
    .Q(\design_top.core0.REG1[10][0] ),
    .CLK(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15216_ (.D(_03301_),
    .Q(\design_top.core0.REG1[10][1] ),
    .CLK(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15217_ (.D(_03302_),
    .Q(\design_top.core0.REG1[10][2] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15218_ (.D(_03303_),
    .Q(\design_top.core0.REG1[10][3] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15219_ (.D(_03304_),
    .Q(\design_top.core0.REG1[10][4] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15220_ (.D(_03305_),
    .Q(\design_top.core0.REG1[10][5] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15221_ (.D(_03306_),
    .Q(\design_top.core0.REG1[10][6] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15222_ (.D(_03307_),
    .Q(\design_top.core0.REG1[10][7] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15223_ (.D(_03308_),
    .Q(\design_top.core0.REG1[10][8] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15224_ (.D(_03309_),
    .Q(\design_top.core0.REG1[10][9] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15225_ (.D(_03310_),
    .Q(\design_top.core0.REG1[10][10] ),
    .CLK(clknet_leaf_143_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15226_ (.D(_03311_),
    .Q(\design_top.core0.REG1[10][11] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15227_ (.D(_03312_),
    .Q(\design_top.core0.REG1[10][12] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15228_ (.D(_03313_),
    .Q(\design_top.core0.REG1[10][13] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15229_ (.D(_03314_),
    .Q(\design_top.core0.REG1[10][14] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15230_ (.D(_03315_),
    .Q(\design_top.core0.REG1[10][15] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15231_ (.D(_03316_),
    .Q(\design_top.core0.REG1[10][16] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15232_ (.D(_03317_),
    .Q(\design_top.core0.REG1[10][17] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15233_ (.D(_03318_),
    .Q(\design_top.core0.REG1[10][18] ),
    .CLK(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15234_ (.D(_03319_),
    .Q(\design_top.core0.REG1[10][19] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15235_ (.D(_03320_),
    .Q(\design_top.core0.REG1[10][20] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15236_ (.D(_03321_),
    .Q(\design_top.core0.REG1[10][21] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15237_ (.D(_03322_),
    .Q(\design_top.core0.REG1[10][22] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15238_ (.D(_03323_),
    .Q(\design_top.core0.REG1[10][23] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15239_ (.D(_03324_),
    .Q(\design_top.core0.REG1[10][24] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15240_ (.D(_03325_),
    .Q(\design_top.core0.REG1[10][25] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15241_ (.D(_03326_),
    .Q(\design_top.core0.REG1[10][26] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15242_ (.D(_03327_),
    .Q(\design_top.core0.REG1[10][27] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15243_ (.D(_03328_),
    .Q(\design_top.core0.REG1[10][28] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15244_ (.D(_03329_),
    .Q(\design_top.core0.REG1[10][29] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15245_ (.D(_03330_),
    .Q(\design_top.core0.REG1[10][30] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15246_ (.D(_03331_),
    .Q(\design_top.core0.REG1[10][31] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15247_ (.D(_03332_),
    .Q(\design_top.core0.REG1[0][0] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15248_ (.D(_03333_),
    .Q(\design_top.core0.REG1[0][1] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15249_ (.D(_03334_),
    .Q(\design_top.core0.REG1[0][2] ),
    .CLK(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15250_ (.D(_03335_),
    .Q(\design_top.core0.REG1[0][3] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15251_ (.D(_03336_),
    .Q(\design_top.core0.REG1[0][4] ),
    .CLK(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15252_ (.D(_03337_),
    .Q(\design_top.core0.REG1[0][5] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15253_ (.D(_03338_),
    .Q(\design_top.core0.REG1[0][6] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15254_ (.D(_03339_),
    .Q(\design_top.core0.REG1[0][7] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15255_ (.D(_03340_),
    .Q(\design_top.core0.REG1[0][8] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15256_ (.D(_03341_),
    .Q(\design_top.core0.REG1[0][9] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15257_ (.D(_03342_),
    .Q(\design_top.core0.REG1[0][10] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15258_ (.D(_03343_),
    .Q(\design_top.core0.REG1[0][11] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15259_ (.D(_03344_),
    .Q(\design_top.core0.REG1[0][12] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15260_ (.D(_03345_),
    .Q(\design_top.core0.REG1[0][13] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15261_ (.D(_03346_),
    .Q(\design_top.core0.REG1[0][14] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15262_ (.D(_03347_),
    .Q(\design_top.core0.REG1[0][15] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15263_ (.D(_03348_),
    .Q(\design_top.core0.REG1[0][16] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15264_ (.D(_03349_),
    .Q(\design_top.core0.REG1[0][17] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15265_ (.D(_03350_),
    .Q(\design_top.core0.REG1[0][18] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15266_ (.D(_03351_),
    .Q(\design_top.core0.REG1[0][19] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15267_ (.D(_03352_),
    .Q(\design_top.core0.REG1[0][20] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15268_ (.D(_03353_),
    .Q(\design_top.core0.REG1[0][21] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15269_ (.D(_03354_),
    .Q(\design_top.core0.REG1[0][22] ),
    .CLK(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15270_ (.D(_03355_),
    .Q(\design_top.core0.REG1[0][23] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15271_ (.D(_03356_),
    .Q(\design_top.core0.REG1[0][24] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15272_ (.D(_03357_),
    .Q(\design_top.core0.REG1[0][25] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15273_ (.D(_03358_),
    .Q(\design_top.core0.REG1[0][26] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15274_ (.D(_03359_),
    .Q(\design_top.core0.REG1[0][27] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15275_ (.D(_03360_),
    .Q(\design_top.core0.REG1[0][28] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15276_ (.D(_03361_),
    .Q(\design_top.core0.REG1[0][29] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15277_ (.D(_03362_),
    .Q(\design_top.core0.REG1[0][30] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15278_ (.D(_03363_),
    .Q(\design_top.core0.REG1[0][31] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15279_ (.D(_03364_),
    .Q(\design_top.core0.REG1[8][0] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15280_ (.D(_03365_),
    .Q(\design_top.core0.REG1[8][1] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15281_ (.D(_03366_),
    .Q(\design_top.core0.REG1[8][2] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15282_ (.D(_03367_),
    .Q(\design_top.core0.REG1[8][3] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15283_ (.D(_03368_),
    .Q(\design_top.core0.REG1[8][4] ),
    .CLK(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15284_ (.D(_03369_),
    .Q(\design_top.core0.REG1[8][5] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15285_ (.D(_03370_),
    .Q(\design_top.core0.REG1[8][6] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15286_ (.D(_03371_),
    .Q(\design_top.core0.REG1[8][7] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15287_ (.D(_03372_),
    .Q(\design_top.core0.REG1[8][8] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15288_ (.D(_03373_),
    .Q(\design_top.core0.REG1[8][9] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15289_ (.D(_03374_),
    .Q(\design_top.core0.REG1[8][10] ),
    .CLK(clknet_leaf_143_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15290_ (.D(_03375_),
    .Q(\design_top.core0.REG1[8][11] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15291_ (.D(_03376_),
    .Q(\design_top.core0.REG1[8][12] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15292_ (.D(_03377_),
    .Q(\design_top.core0.REG1[8][13] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15293_ (.D(_03378_),
    .Q(\design_top.core0.REG1[8][14] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15294_ (.D(_03379_),
    .Q(\design_top.core0.REG1[8][15] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15295_ (.D(_03380_),
    .Q(\design_top.core0.REG1[8][16] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15296_ (.D(_03381_),
    .Q(\design_top.core0.REG1[8][17] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15297_ (.D(_03382_),
    .Q(\design_top.core0.REG1[8][18] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15298_ (.D(_03383_),
    .Q(\design_top.core0.REG1[8][19] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15299_ (.D(_03384_),
    .Q(\design_top.core0.REG1[8][20] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15300_ (.D(_03385_),
    .Q(\design_top.core0.REG1[8][21] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15301_ (.D(_03386_),
    .Q(\design_top.core0.REG1[8][22] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15302_ (.D(_03387_),
    .Q(\design_top.core0.REG1[8][23] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15303_ (.D(_03388_),
    .Q(\design_top.core0.REG1[8][24] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15304_ (.D(_03389_),
    .Q(\design_top.core0.REG1[8][25] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15305_ (.D(_03390_),
    .Q(\design_top.core0.REG1[8][26] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15306_ (.D(_03391_),
    .Q(\design_top.core0.REG1[8][27] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15307_ (.D(_03392_),
    .Q(\design_top.core0.REG1[8][28] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15308_ (.D(_03393_),
    .Q(\design_top.core0.REG1[8][29] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15309_ (.D(_03394_),
    .Q(\design_top.core0.REG1[8][30] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15310_ (.D(_03395_),
    .Q(\design_top.core0.REG1[8][31] ),
    .CLK(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15311_ (.D(_03396_),
    .Q(\design_top.MEM[4][0] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15312_ (.D(_03397_),
    .Q(\design_top.MEM[4][1] ),
    .CLK(clknet_leaf_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15313_ (.D(_03398_),
    .Q(\design_top.MEM[4][2] ),
    .CLK(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15314_ (.D(_03399_),
    .Q(\design_top.MEM[4][3] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15315_ (.D(_03400_),
    .Q(\design_top.MEM[4][4] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15316_ (.D(_03401_),
    .Q(\design_top.MEM[4][5] ),
    .CLK(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15317_ (.D(_03402_),
    .Q(\design_top.MEM[4][6] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15318_ (.D(_03403_),
    .Q(\design_top.MEM[4][7] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15319_ (.D(_03404_),
    .Q(\design_top.core0.REG1[7][0] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15320_ (.D(_03405_),
    .Q(\design_top.core0.REG1[7][1] ),
    .CLK(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15321_ (.D(_03406_),
    .Q(\design_top.core0.REG1[7][2] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15322_ (.D(_03407_),
    .Q(\design_top.core0.REG1[7][3] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15323_ (.D(_03408_),
    .Q(\design_top.core0.REG1[7][4] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15324_ (.D(_03409_),
    .Q(\design_top.core0.REG1[7][5] ),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15325_ (.D(_03410_),
    .Q(\design_top.core0.REG1[7][6] ),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15326_ (.D(_03411_),
    .Q(\design_top.core0.REG1[7][7] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15327_ (.D(_03412_),
    .Q(\design_top.core0.REG1[7][8] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15328_ (.D(_03413_),
    .Q(\design_top.core0.REG1[7][9] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15329_ (.D(_03414_),
    .Q(\design_top.core0.REG1[7][10] ),
    .CLK(clknet_leaf_143_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15330_ (.D(_03415_),
    .Q(\design_top.core0.REG1[7][11] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15331_ (.D(_03416_),
    .Q(\design_top.core0.REG1[7][12] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15332_ (.D(_03417_),
    .Q(\design_top.core0.REG1[7][13] ),
    .CLK(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15333_ (.D(_03418_),
    .Q(\design_top.core0.REG1[7][14] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15334_ (.D(_03419_),
    .Q(\design_top.core0.REG1[7][15] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15335_ (.D(_03420_),
    .Q(\design_top.core0.REG1[7][16] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15336_ (.D(_03421_),
    .Q(\design_top.core0.REG1[7][17] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15337_ (.D(_03422_),
    .Q(\design_top.core0.REG1[7][18] ),
    .CLK(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15338_ (.D(_03423_),
    .Q(\design_top.core0.REG1[7][19] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15339_ (.D(_03424_),
    .Q(\design_top.core0.REG1[7][20] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15340_ (.D(_03425_),
    .Q(\design_top.core0.REG1[7][21] ),
    .CLK(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15341_ (.D(_03426_),
    .Q(\design_top.core0.REG1[7][22] ),
    .CLK(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15342_ (.D(_03427_),
    .Q(\design_top.core0.REG1[7][23] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15343_ (.D(_03428_),
    .Q(\design_top.core0.REG1[7][24] ),
    .CLK(clknet_leaf_84_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15344_ (.D(_03429_),
    .Q(\design_top.core0.REG1[7][25] ),
    .CLK(clknet_leaf_84_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15345_ (.D(_03430_),
    .Q(\design_top.core0.REG1[7][26] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15346_ (.D(_03431_),
    .Q(\design_top.core0.REG1[7][27] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15347_ (.D(_03432_),
    .Q(\design_top.core0.REG1[7][28] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15348_ (.D(_03433_),
    .Q(\design_top.core0.REG1[7][29] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15349_ (.D(_03434_),
    .Q(\design_top.core0.REG1[7][30] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15350_ (.D(_03435_),
    .Q(\design_top.core0.REG1[7][31] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15351_ (.D(_03436_),
    .Q(\design_top.core0.REG1[6][0] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15352_ (.D(_03437_),
    .Q(\design_top.core0.REG1[6][1] ),
    .CLK(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15353_ (.D(_03438_),
    .Q(\design_top.core0.REG1[6][2] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15354_ (.D(_03439_),
    .Q(\design_top.core0.REG1[6][3] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15355_ (.D(_03440_),
    .Q(\design_top.core0.REG1[6][4] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15356_ (.D(_03441_),
    .Q(\design_top.core0.REG1[6][5] ),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15357_ (.D(_03442_),
    .Q(\design_top.core0.REG1[6][6] ),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15358_ (.D(_03443_),
    .Q(\design_top.core0.REG1[6][7] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15359_ (.D(_03444_),
    .Q(\design_top.core0.REG1[6][8] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15360_ (.D(_03445_),
    .Q(\design_top.core0.REG1[6][9] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15361_ (.D(_03446_),
    .Q(\design_top.core0.REG1[6][10] ),
    .CLK(clknet_leaf_143_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15362_ (.D(_03447_),
    .Q(\design_top.core0.REG1[6][11] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15363_ (.D(_03448_),
    .Q(\design_top.core0.REG1[6][12] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15364_ (.D(_03449_),
    .Q(\design_top.core0.REG1[6][13] ),
    .CLK(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15365_ (.D(_03450_),
    .Q(\design_top.core0.REG1[6][14] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15366_ (.D(_03451_),
    .Q(\design_top.core0.REG1[6][15] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15367_ (.D(_03452_),
    .Q(\design_top.core0.REG1[6][16] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15368_ (.D(_03453_),
    .Q(\design_top.core0.REG1[6][17] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15369_ (.D(_03454_),
    .Q(\design_top.core0.REG1[6][18] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15370_ (.D(_03455_),
    .Q(\design_top.core0.REG1[6][19] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15371_ (.D(_03456_),
    .Q(\design_top.core0.REG1[6][20] ),
    .CLK(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15372_ (.D(_03457_),
    .Q(\design_top.core0.REG1[6][21] ),
    .CLK(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15373_ (.D(_03458_),
    .Q(\design_top.core0.REG1[6][22] ),
    .CLK(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15374_ (.D(_03459_),
    .Q(\design_top.core0.REG1[6][23] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15375_ (.D(_03460_),
    .Q(\design_top.core0.REG1[6][24] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15376_ (.D(_03461_),
    .Q(\design_top.core0.REG1[6][25] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15377_ (.D(_03462_),
    .Q(\design_top.core0.REG1[6][26] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15378_ (.D(_03463_),
    .Q(\design_top.core0.REG1[6][27] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15379_ (.D(_03464_),
    .Q(\design_top.core0.REG1[6][28] ),
    .CLK(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15380_ (.D(_03465_),
    .Q(\design_top.core0.REG1[6][29] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15381_ (.D(_03466_),
    .Q(\design_top.core0.REG1[6][30] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15382_ (.D(_03467_),
    .Q(\design_top.core0.REG1[6][31] ),
    .CLK(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15383_ (.D(_03468_),
    .Q(\design_top.core0.REG1[5][0] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15384_ (.D(_03469_),
    .Q(\design_top.core0.REG1[5][1] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15385_ (.D(_03470_),
    .Q(\design_top.core0.REG1[5][2] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15386_ (.D(_03471_),
    .Q(\design_top.core0.REG1[5][3] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15387_ (.D(_03472_),
    .Q(\design_top.core0.REG1[5][4] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15388_ (.D(_03473_),
    .Q(\design_top.core0.REG1[5][5] ),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15389_ (.D(_03474_),
    .Q(\design_top.core0.REG1[5][6] ),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15390_ (.D(_03475_),
    .Q(\design_top.core0.REG1[5][7] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15391_ (.D(_03476_),
    .Q(\design_top.core0.REG1[5][8] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15392_ (.D(_03477_),
    .Q(\design_top.core0.REG1[5][9] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15393_ (.D(_03478_),
    .Q(\design_top.core0.REG1[5][10] ),
    .CLK(clknet_leaf_143_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15394_ (.D(_03479_),
    .Q(\design_top.core0.REG1[5][11] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15395_ (.D(_03480_),
    .Q(\design_top.core0.REG1[5][12] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15396_ (.D(_03481_),
    .Q(\design_top.core0.REG1[5][13] ),
    .CLK(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15397_ (.D(_03482_),
    .Q(\design_top.core0.REG1[5][14] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15398_ (.D(_03483_),
    .Q(\design_top.core0.REG1[5][15] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15399_ (.D(_03484_),
    .Q(\design_top.core0.REG1[5][16] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15400_ (.D(_03485_),
    .Q(\design_top.core0.REG1[5][17] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15401_ (.D(_03486_),
    .Q(\design_top.core0.REG1[5][18] ),
    .CLK(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15402_ (.D(_03487_),
    .Q(\design_top.core0.REG1[5][19] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15403_ (.D(_03488_),
    .Q(\design_top.core0.REG1[5][20] ),
    .CLK(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15404_ (.D(_03489_),
    .Q(\design_top.core0.REG1[5][21] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15405_ (.D(_03490_),
    .Q(\design_top.core0.REG1[5][22] ),
    .CLK(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15406_ (.D(_03491_),
    .Q(\design_top.core0.REG1[5][23] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15407_ (.D(_03492_),
    .Q(\design_top.core0.REG1[5][24] ),
    .CLK(clknet_leaf_84_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15408_ (.D(_03493_),
    .Q(\design_top.core0.REG1[5][25] ),
    .CLK(clknet_leaf_84_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15409_ (.D(_03494_),
    .Q(\design_top.core0.REG1[5][26] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15410_ (.D(_03495_),
    .Q(\design_top.core0.REG1[5][27] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15411_ (.D(_03496_),
    .Q(\design_top.core0.REG1[5][28] ),
    .CLK(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15412_ (.D(_03497_),
    .Q(\design_top.core0.REG1[5][29] ),
    .CLK(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15413_ (.D(_03498_),
    .Q(\design_top.core0.REG1[5][30] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15414_ (.D(_03499_),
    .Q(\design_top.core0.REG1[5][31] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15415_ (.D(_03500_),
    .Q(\design_top.core0.REG1[4][0] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15416_ (.D(_03501_),
    .Q(\design_top.core0.REG1[4][1] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15417_ (.D(_03502_),
    .Q(\design_top.core0.REG1[4][2] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15418_ (.D(_03503_),
    .Q(\design_top.core0.REG1[4][3] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15419_ (.D(_03504_),
    .Q(\design_top.core0.REG1[4][4] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15420_ (.D(_03505_),
    .Q(\design_top.core0.REG1[4][5] ),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15421_ (.D(_03506_),
    .Q(\design_top.core0.REG1[4][6] ),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15422_ (.D(_03507_),
    .Q(\design_top.core0.REG1[4][7] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15423_ (.D(_03508_),
    .Q(\design_top.core0.REG1[4][8] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15424_ (.D(_03509_),
    .Q(\design_top.core0.REG1[4][9] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15425_ (.D(_03510_),
    .Q(\design_top.core0.REG1[4][10] ),
    .CLK(clknet_leaf_143_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15426_ (.D(_03511_),
    .Q(\design_top.core0.REG1[4][11] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15427_ (.D(_03512_),
    .Q(\design_top.core0.REG1[4][12] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15428_ (.D(_03513_),
    .Q(\design_top.core0.REG1[4][13] ),
    .CLK(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15429_ (.D(_03514_),
    .Q(\design_top.core0.REG1[4][14] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15430_ (.D(_03515_),
    .Q(\design_top.core0.REG1[4][15] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15431_ (.D(_03516_),
    .Q(\design_top.core0.REG1[4][16] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15432_ (.D(_03517_),
    .Q(\design_top.core0.REG1[4][17] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15433_ (.D(_03518_),
    .Q(\design_top.core0.REG1[4][18] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15434_ (.D(_03519_),
    .Q(\design_top.core0.REG1[4][19] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15435_ (.D(_03520_),
    .Q(\design_top.core0.REG1[4][20] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15436_ (.D(_03521_),
    .Q(\design_top.core0.REG1[4][21] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15437_ (.D(_03522_),
    .Q(\design_top.core0.REG1[4][22] ),
    .CLK(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15438_ (.D(_03523_),
    .Q(\design_top.core0.REG1[4][23] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15439_ (.D(_03524_),
    .Q(\design_top.core0.REG1[4][24] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15440_ (.D(_03525_),
    .Q(\design_top.core0.REG1[4][25] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15441_ (.D(_03526_),
    .Q(\design_top.core0.REG1[4][26] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15442_ (.D(_03527_),
    .Q(\design_top.core0.REG1[4][27] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15443_ (.D(_03528_),
    .Q(\design_top.core0.REG1[4][28] ),
    .CLK(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15444_ (.D(_03529_),
    .Q(\design_top.core0.REG1[4][29] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15445_ (.D(_03530_),
    .Q(\design_top.core0.REG1[4][30] ),
    .CLK(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15446_ (.D(_03531_),
    .Q(\design_top.core0.REG1[4][31] ),
    .CLK(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15447_ (.D(_03532_),
    .Q(\design_top.core0.REG1[3][0] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15448_ (.D(_03533_),
    .Q(\design_top.core0.REG1[3][1] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15449_ (.D(_03534_),
    .Q(\design_top.core0.REG1[3][2] ),
    .CLK(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15450_ (.D(_03535_),
    .Q(\design_top.core0.REG1[3][3] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15451_ (.D(_03536_),
    .Q(\design_top.core0.REG1[3][4] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15452_ (.D(_03537_),
    .Q(\design_top.core0.REG1[3][5] ),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15453_ (.D(_03538_),
    .Q(\design_top.core0.REG1[3][6] ),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15454_ (.D(_03539_),
    .Q(\design_top.core0.REG1[3][7] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15455_ (.D(_03540_),
    .Q(\design_top.core0.REG1[3][8] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15456_ (.D(_03541_),
    .Q(\design_top.core0.REG1[3][9] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15457_ (.D(_03542_),
    .Q(\design_top.core0.REG1[3][10] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15458_ (.D(_03543_),
    .Q(\design_top.core0.REG1[3][11] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15459_ (.D(_03544_),
    .Q(\design_top.core0.REG1[3][12] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15460_ (.D(_03545_),
    .Q(\design_top.core0.REG1[3][13] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15461_ (.D(_03546_),
    .Q(\design_top.core0.REG1[3][14] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15462_ (.D(_03547_),
    .Q(\design_top.core0.REG1[3][15] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15463_ (.D(_03548_),
    .Q(\design_top.core0.REG1[3][16] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15464_ (.D(_03549_),
    .Q(\design_top.core0.REG1[3][17] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15465_ (.D(_03550_),
    .Q(\design_top.core0.REG1[3][18] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15466_ (.D(_03551_),
    .Q(\design_top.core0.REG1[3][19] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15467_ (.D(_03552_),
    .Q(\design_top.core0.REG1[3][20] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15468_ (.D(_03553_),
    .Q(\design_top.core0.REG1[3][21] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15469_ (.D(_03554_),
    .Q(\design_top.core0.REG1[3][22] ),
    .CLK(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15470_ (.D(_03555_),
    .Q(\design_top.core0.REG1[3][23] ),
    .CLK(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15471_ (.D(_03556_),
    .Q(\design_top.core0.REG1[3][24] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15472_ (.D(_03557_),
    .Q(\design_top.core0.REG1[3][25] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15473_ (.D(_03558_),
    .Q(\design_top.core0.REG1[3][26] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15474_ (.D(_03559_),
    .Q(\design_top.core0.REG1[3][27] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15475_ (.D(_03560_),
    .Q(\design_top.core0.REG1[3][28] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15476_ (.D(_03561_),
    .Q(\design_top.core0.REG1[3][29] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15477_ (.D(_03562_),
    .Q(\design_top.core0.REG1[3][30] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15478_ (.D(_03563_),
    .Q(\design_top.core0.REG1[3][31] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15479_ (.D(_03564_),
    .Q(\design_top.core0.REG1[2][0] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15480_ (.D(_03565_),
    .Q(\design_top.core0.REG1[2][1] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15481_ (.D(_03566_),
    .Q(\design_top.core0.REG1[2][2] ),
    .CLK(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15482_ (.D(_03567_),
    .Q(\design_top.core0.REG1[2][3] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15483_ (.D(_03568_),
    .Q(\design_top.core0.REG1[2][4] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15484_ (.D(_03569_),
    .Q(\design_top.core0.REG1[2][5] ),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15485_ (.D(_03570_),
    .Q(\design_top.core0.REG1[2][6] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15486_ (.D(_03571_),
    .Q(\design_top.core0.REG1[2][7] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15487_ (.D(_03572_),
    .Q(\design_top.core0.REG1[2][8] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15488_ (.D(_03573_),
    .Q(\design_top.core0.REG1[2][9] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15489_ (.D(_03574_),
    .Q(\design_top.core0.REG1[2][10] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15490_ (.D(_03575_),
    .Q(\design_top.core0.REG1[2][11] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15491_ (.D(_03576_),
    .Q(\design_top.core0.REG1[2][12] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15492_ (.D(_03577_),
    .Q(\design_top.core0.REG1[2][13] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15493_ (.D(_03578_),
    .Q(\design_top.core0.REG1[2][14] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15494_ (.D(_03579_),
    .Q(\design_top.core0.REG1[2][15] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15495_ (.D(_03580_),
    .Q(\design_top.core0.REG1[2][16] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15496_ (.D(_03581_),
    .Q(\design_top.core0.REG1[2][17] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15497_ (.D(_03582_),
    .Q(\design_top.core0.REG1[2][18] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15498_ (.D(_03583_),
    .Q(\design_top.core0.REG1[2][19] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15499_ (.D(_03584_),
    .Q(\design_top.core0.REG1[2][20] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15500_ (.D(_03585_),
    .Q(\design_top.core0.REG1[2][21] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15501_ (.D(_03586_),
    .Q(\design_top.core0.REG1[2][22] ),
    .CLK(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15502_ (.D(_03587_),
    .Q(\design_top.core0.REG1[2][23] ),
    .CLK(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15503_ (.D(_03588_),
    .Q(\design_top.core0.REG1[2][24] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15504_ (.D(_03589_),
    .Q(\design_top.core0.REG1[2][25] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15505_ (.D(_03590_),
    .Q(\design_top.core0.REG1[2][26] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15506_ (.D(_03591_),
    .Q(\design_top.core0.REG1[2][27] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15507_ (.D(_03592_),
    .Q(\design_top.core0.REG1[2][28] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15508_ (.D(_03593_),
    .Q(\design_top.core0.REG1[2][29] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15509_ (.D(_03594_),
    .Q(\design_top.core0.REG1[2][30] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15510_ (.D(_03595_),
    .Q(\design_top.core0.REG1[2][31] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15511_ (.D(_03596_),
    .Q(\design_top.core0.REG1[1][0] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15512_ (.D(_03597_),
    .Q(\design_top.core0.REG1[1][1] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15513_ (.D(_03598_),
    .Q(\design_top.core0.REG1[1][2] ),
    .CLK(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15514_ (.D(_03599_),
    .Q(\design_top.core0.REG1[1][3] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15515_ (.D(_03600_),
    .Q(\design_top.core0.REG1[1][4] ),
    .CLK(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15516_ (.D(_03601_),
    .Q(\design_top.core0.REG1[1][5] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15517_ (.D(_03602_),
    .Q(\design_top.core0.REG1[1][6] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15518_ (.D(_03603_),
    .Q(\design_top.core0.REG1[1][7] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15519_ (.D(_03604_),
    .Q(\design_top.core0.REG1[1][8] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15520_ (.D(_03605_),
    .Q(\design_top.core0.REG1[1][9] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15521_ (.D(_03606_),
    .Q(\design_top.core0.REG1[1][10] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15522_ (.D(_03607_),
    .Q(\design_top.core0.REG1[1][11] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15523_ (.D(_03608_),
    .Q(\design_top.core0.REG1[1][12] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15524_ (.D(_03609_),
    .Q(\design_top.core0.REG1[1][13] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15525_ (.D(_03610_),
    .Q(\design_top.core0.REG1[1][14] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15526_ (.D(_03611_),
    .Q(\design_top.core0.REG1[1][15] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15527_ (.D(_03612_),
    .Q(\design_top.core0.REG1[1][16] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15528_ (.D(_03613_),
    .Q(\design_top.core0.REG1[1][17] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15529_ (.D(_03614_),
    .Q(\design_top.core0.REG1[1][18] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15530_ (.D(_03615_),
    .Q(\design_top.core0.REG1[1][19] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15531_ (.D(_03616_),
    .Q(\design_top.core0.REG1[1][20] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15532_ (.D(_03617_),
    .Q(\design_top.core0.REG1[1][21] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15533_ (.D(_03618_),
    .Q(\design_top.core0.REG1[1][22] ),
    .CLK(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15534_ (.D(_03619_),
    .Q(\design_top.core0.REG1[1][23] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15535_ (.D(_03620_),
    .Q(\design_top.core0.REG1[1][24] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15536_ (.D(_03621_),
    .Q(\design_top.core0.REG1[1][25] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15537_ (.D(_03622_),
    .Q(\design_top.core0.REG1[1][26] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15538_ (.D(_03623_),
    .Q(\design_top.core0.REG1[1][27] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15539_ (.D(_03624_),
    .Q(\design_top.core0.REG1[1][28] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15540_ (.D(_03625_),
    .Q(\design_top.core0.REG1[1][29] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15541_ (.D(_03626_),
    .Q(\design_top.core0.REG1[1][30] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15542_ (.D(_03627_),
    .Q(\design_top.core0.REG1[1][31] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15543_ (.D(_03628_),
    .Q(\design_top.core0.REG1[15][0] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15544_ (.D(_03629_),
    .Q(\design_top.core0.REG1[15][1] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15545_ (.D(_03630_),
    .Q(\design_top.core0.REG1[15][2] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15546_ (.D(_03631_),
    .Q(\design_top.core0.REG1[15][3] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15547_ (.D(_03632_),
    .Q(\design_top.core0.REG1[15][4] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15548_ (.D(_03633_),
    .Q(\design_top.core0.REG1[15][5] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15549_ (.D(_03634_),
    .Q(\design_top.core0.REG1[15][6] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15550_ (.D(_03635_),
    .Q(\design_top.core0.REG1[15][7] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15551_ (.D(_03636_),
    .Q(\design_top.core0.REG1[15][8] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15552_ (.D(_03637_),
    .Q(\design_top.core0.REG1[15][9] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15553_ (.D(_03638_),
    .Q(\design_top.core0.REG1[15][10] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15554_ (.D(_03639_),
    .Q(\design_top.core0.REG1[15][11] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15555_ (.D(_03640_),
    .Q(\design_top.core0.REG1[15][12] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15556_ (.D(_03641_),
    .Q(\design_top.core0.REG1[15][13] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15557_ (.D(_03642_),
    .Q(\design_top.core0.REG1[15][14] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15558_ (.D(_03643_),
    .Q(\design_top.core0.REG1[15][15] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15559_ (.D(_03644_),
    .Q(\design_top.core0.REG1[15][16] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15560_ (.D(_03645_),
    .Q(\design_top.core0.REG1[15][17] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15561_ (.D(_03646_),
    .Q(\design_top.core0.REG1[15][18] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15562_ (.D(_03647_),
    .Q(\design_top.core0.REG1[15][19] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15563_ (.D(_03648_),
    .Q(\design_top.core0.REG1[15][20] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15564_ (.D(_03649_),
    .Q(\design_top.core0.REG1[15][21] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15565_ (.D(_03650_),
    .Q(\design_top.core0.REG1[15][22] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15566_ (.D(_03651_),
    .Q(\design_top.core0.REG1[15][23] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15567_ (.D(_03652_),
    .Q(\design_top.core0.REG1[15][24] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15568_ (.D(_03653_),
    .Q(\design_top.core0.REG1[15][25] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15569_ (.D(_03654_),
    .Q(\design_top.core0.REG1[15][26] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15570_ (.D(_03655_),
    .Q(\design_top.core0.REG1[15][27] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15571_ (.D(_03656_),
    .Q(\design_top.core0.REG1[15][28] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15572_ (.D(_03657_),
    .Q(\design_top.core0.REG1[15][29] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15573_ (.D(_03658_),
    .Q(\design_top.core0.REG1[15][30] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15574_ (.D(_03659_),
    .Q(\design_top.core0.REG1[15][31] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15575_ (.D(_03660_),
    .Q(\design_top.MEM[3][0] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15576_ (.D(_03661_),
    .Q(\design_top.MEM[3][1] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15577_ (.D(_03662_),
    .Q(\design_top.MEM[3][2] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15578_ (.D(_03663_),
    .Q(\design_top.MEM[3][3] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15579_ (.D(_03664_),
    .Q(\design_top.MEM[3][4] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15580_ (.D(_03665_),
    .Q(\design_top.MEM[3][5] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15581_ (.D(_03666_),
    .Q(\design_top.MEM[3][6] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15582_ (.D(_03667_),
    .Q(\design_top.MEM[3][7] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15583_ (.D(_03668_),
    .Q(\design_top.MEM[2][0] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15584_ (.D(_03669_),
    .Q(\design_top.MEM[2][1] ),
    .CLK(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15585_ (.D(_03670_),
    .Q(\design_top.MEM[2][2] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15586_ (.D(_03671_),
    .Q(\design_top.MEM[2][3] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15587_ (.D(_03672_),
    .Q(\design_top.MEM[2][4] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15588_ (.D(_03673_),
    .Q(\design_top.MEM[2][5] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15589_ (.D(_03674_),
    .Q(\design_top.MEM[2][6] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15590_ (.D(_03675_),
    .Q(\design_top.MEM[2][7] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15591_ (.D(_03676_),
    .Q(\design_top.MEM[1][0] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15592_ (.D(_03677_),
    .Q(\design_top.MEM[1][1] ),
    .CLK(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15593_ (.D(_03678_),
    .Q(\design_top.MEM[1][2] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15594_ (.D(_03679_),
    .Q(\design_top.MEM[1][3] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15595_ (.D(_03680_),
    .Q(\design_top.MEM[1][4] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15596_ (.D(_03681_),
    .Q(\design_top.MEM[1][5] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15597_ (.D(_03682_),
    .Q(\design_top.MEM[1][6] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15598_ (.D(_03683_),
    .Q(\design_top.MEM[1][7] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15599_ (.D(_03684_),
    .Q(\design_top.MEM[15][0] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15600_ (.D(_03685_),
    .Q(\design_top.MEM[15][1] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15601_ (.D(_03686_),
    .Q(\design_top.MEM[15][2] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15602_ (.D(_03687_),
    .Q(\design_top.MEM[15][3] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15603_ (.D(_03688_),
    .Q(\design_top.MEM[15][4] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15604_ (.D(_03689_),
    .Q(\design_top.MEM[15][5] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15605_ (.D(_03690_),
    .Q(\design_top.MEM[15][6] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15606_ (.D(_03691_),
    .Q(\design_top.MEM[15][7] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15607_ (.D(_03692_),
    .Q(\design_top.core0.REG1[9][0] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15608_ (.D(_03693_),
    .Q(\design_top.core0.REG1[9][1] ),
    .CLK(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15609_ (.D(_03694_),
    .Q(\design_top.core0.REG1[9][2] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15610_ (.D(_03695_),
    .Q(\design_top.core0.REG1[9][3] ),
    .CLK(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15611_ (.D(_03696_),
    .Q(\design_top.core0.REG1[9][4] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15612_ (.D(_03697_),
    .Q(\design_top.core0.REG1[9][5] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15613_ (.D(_03698_),
    .Q(\design_top.core0.REG1[9][6] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15614_ (.D(_03699_),
    .Q(\design_top.core0.REG1[9][7] ),
    .CLK(clknet_leaf_143_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15615_ (.D(_03700_),
    .Q(\design_top.core0.REG1[9][8] ),
    .CLK(clknet_leaf_143_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15616_ (.D(_03701_),
    .Q(\design_top.core0.REG1[9][9] ),
    .CLK(clknet_leaf_143_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15617_ (.D(_03702_),
    .Q(\design_top.core0.REG1[9][10] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15618_ (.D(_03703_),
    .Q(\design_top.core0.REG1[9][11] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15619_ (.D(_03704_),
    .Q(\design_top.core0.REG1[9][12] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15620_ (.D(_03705_),
    .Q(\design_top.core0.REG1[9][13] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15621_ (.D(_03706_),
    .Q(\design_top.core0.REG1[9][14] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15622_ (.D(_03707_),
    .Q(\design_top.core0.REG1[9][15] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15623_ (.D(_03708_),
    .Q(\design_top.core0.REG1[9][16] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15624_ (.D(_03709_),
    .Q(\design_top.core0.REG1[9][17] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15625_ (.D(_03710_),
    .Q(\design_top.core0.REG1[9][18] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15626_ (.D(_03711_),
    .Q(\design_top.core0.REG1[9][19] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15627_ (.D(_03712_),
    .Q(\design_top.core0.REG1[9][20] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15628_ (.D(_03713_),
    .Q(\design_top.core0.REG1[9][21] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15629_ (.D(_03714_),
    .Q(\design_top.core0.REG1[9][22] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15630_ (.D(_03715_),
    .Q(\design_top.core0.REG1[9][23] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15631_ (.D(_03716_),
    .Q(\design_top.core0.REG1[9][24] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15632_ (.D(_03717_),
    .Q(\design_top.core0.REG1[9][25] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15633_ (.D(_03718_),
    .Q(\design_top.core0.REG1[9][26] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15634_ (.D(_03719_),
    .Q(\design_top.core0.REG1[9][27] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15635_ (.D(_03720_),
    .Q(\design_top.core0.REG1[9][28] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15636_ (.D(_03721_),
    .Q(\design_top.core0.REG1[9][29] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15637_ (.D(_03722_),
    .Q(\design_top.core0.REG1[9][30] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15638_ (.D(_03723_),
    .Q(\design_top.core0.REG1[9][31] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15639_ (.D(_03724_),
    .Q(\design_top.MEM[13][0] ),
    .CLK(clknet_leaf_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15640_ (.D(_03725_),
    .Q(\design_top.MEM[13][1] ),
    .CLK(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15641_ (.D(_03726_),
    .Q(\design_top.MEM[13][2] ),
    .CLK(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15642_ (.D(_03727_),
    .Q(\design_top.MEM[13][3] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15643_ (.D(_03728_),
    .Q(\design_top.MEM[13][4] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15644_ (.D(_03729_),
    .Q(\design_top.MEM[13][5] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15645_ (.D(_03730_),
    .Q(\design_top.MEM[13][6] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15646_ (.D(_03731_),
    .Q(\design_top.MEM[13][7] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15647_ (.D(_03732_),
    .Q(io_out[14]),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15648_ (.D(_03733_),
    .Q(\design_top.TIMER[0] ),
    .CLK(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15649_ (.D(_03734_),
    .Q(\design_top.TIMER[1] ),
    .CLK(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15650_ (.D(_03735_),
    .Q(\design_top.TIMER[2] ),
    .CLK(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15651_ (.D(_03736_),
    .Q(\design_top.TIMER[3] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15652_ (.D(_03737_),
    .Q(\design_top.TIMER[4] ),
    .CLK(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15653_ (.D(_03738_),
    .Q(\design_top.TIMER[5] ),
    .CLK(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15654_ (.D(_03739_),
    .Q(\design_top.TIMER[6] ),
    .CLK(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15655_ (.D(_03740_),
    .Q(\design_top.TIMER[7] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15656_ (.D(_03741_),
    .Q(\design_top.TIMER[8] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15657_ (.D(_03742_),
    .Q(\design_top.TIMER[9] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15658_ (.D(_03743_),
    .Q(\design_top.TIMER[10] ),
    .CLK(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15659_ (.D(_03744_),
    .Q(\design_top.TIMER[11] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15660_ (.D(_03745_),
    .Q(\design_top.TIMER[12] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15661_ (.D(_03746_),
    .Q(\design_top.TIMER[13] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15662_ (.D(_03747_),
    .Q(\design_top.TIMER[14] ),
    .CLK(clknet_leaf_172_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15663_ (.D(_03748_),
    .Q(\design_top.TIMER[15] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15664_ (.D(_03749_),
    .Q(\design_top.TIMER[16] ),
    .CLK(clknet_leaf_172_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15665_ (.D(_03750_),
    .Q(\design_top.TIMER[17] ),
    .CLK(clknet_leaf_172_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15666_ (.D(_03751_),
    .Q(\design_top.TIMER[18] ),
    .CLK(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15667_ (.D(_03752_),
    .Q(\design_top.TIMER[19] ),
    .CLK(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15668_ (.D(_03753_),
    .Q(\design_top.TIMER[20] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15669_ (.D(_03754_),
    .Q(\design_top.TIMER[21] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15670_ (.D(_03755_),
    .Q(\design_top.TIMER[22] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15671_ (.D(_03756_),
    .Q(\design_top.TIMER[23] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15672_ (.D(_03757_),
    .Q(\design_top.TIMER[24] ),
    .CLK(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15673_ (.D(_03758_),
    .Q(\design_top.TIMER[25] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15674_ (.D(_03759_),
    .Q(\design_top.TIMER[26] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15675_ (.D(_03760_),
    .Q(\design_top.TIMER[27] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15676_ (.D(_03761_),
    .Q(\design_top.TIMER[28] ),
    .CLK(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15677_ (.D(_03762_),
    .Q(\design_top.TIMER[29] ),
    .CLK(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15678_ (.D(_03763_),
    .Q(\design_top.TIMER[30] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15679_ (.D(_03764_),
    .Q(\design_top.TIMER[31] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15680_ (.D(_03765_),
    .Q(\design_top.MEM[12][0] ),
    .CLK(clknet_leaf_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15681_ (.D(_03766_),
    .Q(\design_top.MEM[12][1] ),
    .CLK(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15682_ (.D(_03767_),
    .Q(\design_top.MEM[12][2] ),
    .CLK(clknet_leaf_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15683_ (.D(_03768_),
    .Q(\design_top.MEM[12][3] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15684_ (.D(_03769_),
    .Q(\design_top.MEM[12][4] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15685_ (.D(_03770_),
    .Q(\design_top.MEM[12][5] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15686_ (.D(_03771_),
    .Q(\design_top.MEM[12][6] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15687_ (.D(_03772_),
    .Q(\design_top.MEM[12][7] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15688_ (.D(_03773_),
    .Q(\design_top.MEM[11][0] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15689_ (.D(_03774_),
    .Q(\design_top.MEM[11][1] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15690_ (.D(_03775_),
    .Q(\design_top.MEM[11][2] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15691_ (.D(_03776_),
    .Q(\design_top.MEM[11][3] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15692_ (.D(_03777_),
    .Q(\design_top.MEM[11][4] ),
    .CLK(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15693_ (.D(_03778_),
    .Q(\design_top.MEM[11][5] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15694_ (.D(_03779_),
    .Q(\design_top.MEM[11][6] ),
    .CLK(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15695_ (.D(_03780_),
    .Q(\design_top.MEM[11][7] ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15696_ (.D(_03781_),
    .Q(\design_top.MEM[10][0] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15697_ (.D(_03782_),
    .Q(\design_top.MEM[10][1] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15698_ (.D(_03783_),
    .Q(\design_top.MEM[10][2] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15699_ (.D(_03784_),
    .Q(\design_top.MEM[10][3] ),
    .CLK(clknet_leaf_235_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15700_ (.D(_03785_),
    .Q(\design_top.MEM[10][4] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15701_ (.D(_03786_),
    .Q(\design_top.MEM[10][5] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15702_ (.D(_03787_),
    .Q(\design_top.MEM[10][6] ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15703_ (.D(_03788_),
    .Q(\design_top.MEM[10][7] ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15704_ (.D(_03789_),
    .Q(\design_top.MEM[0][0] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15705_ (.D(_03790_),
    .Q(\design_top.MEM[0][1] ),
    .CLK(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15706_ (.D(_03791_),
    .Q(\design_top.MEM[0][2] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15707_ (.D(_03792_),
    .Q(\design_top.MEM[0][3] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15708_ (.D(_03793_),
    .Q(\design_top.MEM[0][4] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15709_ (.D(_03794_),
    .Q(\design_top.MEM[0][5] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15710_ (.D(_03795_),
    .Q(\design_top.MEM[0][6] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15711_ (.D(_03796_),
    .Q(\design_top.MEM[0][7] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15712_ (.D(_03797_),
    .Q(\design_top.uart0.UART_XFIFO[0] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15713_ (.D(_03798_),
    .Q(\design_top.uart0.UART_XFIFO[1] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15714_ (.D(_03799_),
    .Q(\design_top.uart0.UART_XFIFO[2] ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15715_ (.D(_03800_),
    .Q(\design_top.uart0.UART_XFIFO[3] ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15716_ (.D(_03801_),
    .Q(\design_top.uart0.UART_XFIFO[4] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15717_ (.D(_03802_),
    .Q(\design_top.uart0.UART_XFIFO[5] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15718_ (.D(_03803_),
    .Q(\design_top.uart0.UART_XFIFO[6] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15719_ (.D(_03804_),
    .Q(\design_top.uart0.UART_XFIFO[7] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15720_ (.D(_03805_),
    .Q(\design_top.uart0.UART_XREQ ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15721_ (.D(_03806_),
    .Q(\design_top.uart0.UART_RACK ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15722_ (.D(_03807_),
    .Q(\design_top.MEM[14][0] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15723_ (.D(_03808_),
    .Q(\design_top.MEM[14][1] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15724_ (.D(_03809_),
    .Q(\design_top.MEM[14][2] ),
    .CLK(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15725_ (.D(_03810_),
    .Q(\design_top.MEM[14][3] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15726_ (.D(_03811_),
    .Q(\design_top.MEM[14][4] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15727_ (.D(_03812_),
    .Q(\design_top.MEM[14][5] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15728_ (.D(_03813_),
    .Q(\design_top.MEM[14][6] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15729_ (.D(_03814_),
    .Q(\design_top.MEM[14][7] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15730_ (.D(_03815_),
    .Q(\design_top.core0.REG2[9][0] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15731_ (.D(_03816_),
    .Q(\design_top.core0.REG2[9][1] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15732_ (.D(_03817_),
    .Q(\design_top.core0.REG2[9][2] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15733_ (.D(_03818_),
    .Q(\design_top.core0.REG2[9][3] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15734_ (.D(_03819_),
    .Q(\design_top.core0.REG2[9][4] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15735_ (.D(_03820_),
    .Q(\design_top.core0.REG2[9][5] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15736_ (.D(_03821_),
    .Q(\design_top.core0.REG2[9][6] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15737_ (.D(_03822_),
    .Q(\design_top.core0.REG2[9][7] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15738_ (.D(_03823_),
    .Q(\design_top.core0.REG2[9][8] ),
    .CLK(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15739_ (.D(_03824_),
    .Q(\design_top.core0.REG2[9][9] ),
    .CLK(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15740_ (.D(_03825_),
    .Q(\design_top.core0.REG2[9][10] ),
    .CLK(clknet_leaf_37_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15741_ (.D(_03826_),
    .Q(\design_top.core0.REG2[9][11] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15742_ (.D(_03827_),
    .Q(\design_top.core0.REG2[9][12] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15743_ (.D(_03828_),
    .Q(\design_top.core0.REG2[9][13] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15744_ (.D(_03829_),
    .Q(\design_top.core0.REG2[9][14] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15745_ (.D(_03830_),
    .Q(\design_top.core0.REG2[9][15] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15746_ (.D(_03831_),
    .Q(\design_top.core0.REG2[9][16] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15747_ (.D(_03832_),
    .Q(\design_top.core0.REG2[9][17] ),
    .CLK(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15748_ (.D(_03833_),
    .Q(\design_top.core0.REG2[9][18] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15749_ (.D(_03834_),
    .Q(\design_top.core0.REG2[9][19] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15750_ (.D(_03835_),
    .Q(\design_top.core0.REG2[9][20] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15751_ (.D(_03836_),
    .Q(\design_top.core0.REG2[9][21] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15752_ (.D(_03837_),
    .Q(\design_top.core0.REG2[9][22] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15753_ (.D(_03838_),
    .Q(\design_top.core0.REG2[9][23] ),
    .CLK(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15754_ (.D(_03839_),
    .Q(\design_top.core0.REG2[9][24] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15755_ (.D(_03840_),
    .Q(\design_top.core0.REG2[9][25] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15756_ (.D(_03841_),
    .Q(\design_top.core0.REG2[9][26] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15757_ (.D(_03842_),
    .Q(\design_top.core0.REG2[9][27] ),
    .CLK(clknet_leaf_48_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15758_ (.D(_03843_),
    .Q(\design_top.core0.REG2[9][28] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15759_ (.D(_03844_),
    .Q(\design_top.core0.REG2[9][29] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15760_ (.D(_03845_),
    .Q(\design_top.core0.REG2[9][30] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15761_ (.D(_03846_),
    .Q(\design_top.core0.REG2[9][31] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15762_ (.D(_03847_),
    .Q(\design_top.IRES[0] ),
    .CLK(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15763_ (.D(_03848_),
    .Q(\design_top.IRES[1] ),
    .CLK(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15764_ (.D(_03849_),
    .Q(\design_top.IRES[2] ),
    .CLK(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15765_ (.D(_03850_),
    .Q(\design_top.IRES[3] ),
    .CLK(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15766_ (.D(_03851_),
    .Q(\design_top.IRES[4] ),
    .CLK(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15767_ (.D(_03852_),
    .Q(\design_top.IRES[5] ),
    .CLK(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15768_ (.D(_03853_),
    .Q(\design_top.IRES[6] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15769_ (.D(_03854_),
    .Q(\design_top.IRES[7] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15770_ (.D(_03855_),
    .Q(\design_top.core0.RESMODE[0] ),
    .CLK(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15771_ (.D(_03856_),
    .Q(\design_top.core0.RESMODE[1] ),
    .CLK(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15772_ (.D(_03857_),
    .Q(\design_top.core0.RESMODE[2] ),
    .CLK(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15773_ (.D(_03858_),
    .Q(\design_top.core0.RESMODE[3] ),
    .CLK(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15774_ (.D(_03859_),
    .Q(\design_top.uart0.UART_RBAUD[1] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15775_ (.D(_03860_),
    .Q(\design_top.uart0.UART_RBAUD[2] ),
    .CLK(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15776_ (.D(_03861_),
    .Q(\design_top.uart0.UART_RBAUD[4] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15777_ (.D(_03862_),
    .Q(\design_top.uart0.UART_RBAUD[6] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15778_ (.D(_03863_),
    .Q(\design_top.uart0.UART_RBAUD[7] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15779_ (.D(_03864_),
    .Q(\design_top.uart0.UART_RBAUD[9] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15780_ (.D(_03865_),
    .Q(\design_top.uart0.UART_RSTATE[0] ),
    .CLK(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15781_ (.D(_03866_),
    .Q(\design_top.uart0.UART_RSTATE[1] ),
    .CLK(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15782_ (.D(_03867_),
    .Q(\design_top.uart0.UART_RSTATE[2] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15783_ (.D(_03868_),
    .Q(\design_top.uart0.UART_RSTATE[3] ),
    .CLK(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15784_ (.D(_03869_),
    .Q(\design_top.uart0.UART_XSTATE[0] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15785_ (.D(_03870_),
    .Q(\design_top.uart0.UART_XSTATE[1] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15786_ (.D(_03871_),
    .Q(\design_top.uart0.UART_XSTATE[2] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15787_ (.D(_03872_),
    .Q(\design_top.uart0.UART_XSTATE[3] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15788_ (.D(_03873_),
    .Q(\design_top.DACK[0] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15789_ (.D(_03874_),
    .Q(\design_top.DACK[1] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15790_ (.D(_03875_),
    .Q(_00301_),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15791_ (.D(_03876_),
    .Q(_00302_),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15792_ (.D(_03877_),
    .Q(_00303_),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15793_ (.D(_03878_),
    .Q(_00304_),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15794_ (.D(_03879_),
    .Q(\design_top.uart0.UART_XBAUD[0] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15795_ (.D(_03880_),
    .Q(\design_top.uart0.UART_XBAUD[1] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15796_ (.D(_03881_),
    .Q(\design_top.uart0.UART_XBAUD[2] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15797_ (.D(_03882_),
    .Q(\design_top.uart0.UART_XBAUD[3] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15798_ (.D(_03883_),
    .Q(\design_top.uart0.UART_XBAUD[4] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15799_ (.D(_03884_),
    .Q(\design_top.uart0.UART_XBAUD[5] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15800_ (.D(_03885_),
    .Q(\design_top.uart0.UART_XBAUD[6] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15801_ (.D(_03886_),
    .Q(\design_top.uart0.UART_XBAUD[7] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15802_ (.D(_03887_),
    .Q(\design_top.uart0.UART_XBAUD[8] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15803_ (.D(_03888_),
    .Q(\design_top.uart0.UART_XBAUD[9] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15804_ (.D(_03889_),
    .Q(\design_top.uart0.UART_XBAUD[10] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15805_ (.D(_03890_),
    .Q(\design_top.uart0.UART_XBAUD[11] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15806_ (.D(_03891_),
    .Q(\design_top.uart0.UART_XBAUD[12] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15807_ (.D(_03892_),
    .Q(\design_top.uart0.UART_XBAUD[13] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15808_ (.D(_03893_),
    .Q(\design_top.uart0.UART_XBAUD[14] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15809_ (.D(_03894_),
    .Q(\design_top.uart0.UART_XBAUD[15] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15810_ (.D(_03895_),
    .Q(\design_top.uart0.UART_RBAUD[0] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15811_ (.D(_03896_),
    .Q(\design_top.uart0.UART_RBAUD[3] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15812_ (.D(_03897_),
    .Q(\design_top.uart0.UART_RBAUD[5] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15813_ (.D(_03898_),
    .Q(\design_top.uart0.UART_RBAUD[8] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15814_ (.D(_03899_),
    .Q(\design_top.uart0.UART_RBAUD[10] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15815_ (.D(_03900_),
    .Q(\design_top.uart0.UART_RBAUD[11] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15816_ (.D(_03901_),
    .Q(\design_top.uart0.UART_RBAUD[12] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15817_ (.D(_03902_),
    .Q(\design_top.uart0.UART_RBAUD[13] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15818_ (.D(_03903_),
    .Q(\design_top.uart0.UART_RBAUD[14] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15819_ (.D(_03904_),
    .Q(\design_top.uart0.UART_RBAUD[15] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15820_ (.D(_03905_),
    .Q(_00305_),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15821_ (.D(_03906_),
    .Q(_00306_),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15822_ (.D(_03907_),
    .Q(_00307_),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15823_ (.D(_03908_),
    .Q(_00308_),
    .CLK(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15824_ (.D(_03909_),
    .Q(\design_top.core0.FLUSH[0] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15825_ (.D(_03910_),
    .Q(\design_top.core0.FLUSH[1] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15826_ (.D(_03911_),
    .Q(io_out[18]),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15827_ (.D(_03912_),
    .Q(io_out[19]),
    .CLK(clknet_leaf_29_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15828_ (.D(_03913_),
    .Q(\design_top.IADDR[4] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15829_ (.D(_03914_),
    .Q(\design_top.IADDR[5] ),
    .CLK(clknet_leaf_29_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15830_ (.D(_03915_),
    .Q(\design_top.IADDR[6] ),
    .CLK(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15831_ (.D(_03916_),
    .Q(\design_top.IADDR[7] ),
    .CLK(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15832_ (.D(_03917_),
    .Q(\design_top.IADDR[8] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15833_ (.D(_03918_),
    .Q(\design_top.IADDR[9] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15834_ (.D(_03919_),
    .Q(\design_top.IADDR[10] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15835_ (.D(_03920_),
    .Q(\design_top.IADDR[11] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15836_ (.D(_03921_),
    .Q(\design_top.IADDR[12] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15837_ (.D(_03922_),
    .Q(\design_top.IADDR[13] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15838_ (.D(_03923_),
    .Q(\design_top.IADDR[14] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15839_ (.D(_03924_),
    .Q(\design_top.IADDR[15] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15840_ (.D(_03925_),
    .Q(\design_top.IADDR[16] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15841_ (.D(_03926_),
    .Q(\design_top.IADDR[17] ),
    .CLK(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15842_ (.D(_03927_),
    .Q(\design_top.IADDR[18] ),
    .CLK(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15843_ (.D(_03928_),
    .Q(\design_top.IADDR[19] ),
    .CLK(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15844_ (.D(_03929_),
    .Q(\design_top.IADDR[20] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15845_ (.D(_03930_),
    .Q(\design_top.IADDR[21] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15846_ (.D(_03931_),
    .Q(\design_top.IADDR[22] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15847_ (.D(_03932_),
    .Q(\design_top.IADDR[23] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15848_ (.D(_03933_),
    .Q(\design_top.IADDR[24] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15849_ (.D(_03934_),
    .Q(\design_top.IADDR[25] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15850_ (.D(_03935_),
    .Q(\design_top.IADDR[26] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15851_ (.D(_03936_),
    .Q(\design_top.IADDR[27] ),
    .CLK(clknet_leaf_39_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15852_ (.D(_03937_),
    .Q(\design_top.IADDR[28] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15853_ (.D(_03938_),
    .Q(\design_top.IADDR[29] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15854_ (.D(_03939_),
    .Q(\design_top.IADDR[30] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15855_ (.D(_03940_),
    .Q(\design_top.IADDR[31] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15856_ (.D(_03941_),
    .Q(\design_top.core0.XIDATA[7] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15857_ (.D(_03942_),
    .Q(\design_top.core0.XIDATA[8] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15858_ (.D(_03943_),
    .Q(\design_top.core0.XIDATA[9] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15859_ (.D(_03944_),
    .Q(\design_top.core0.XIDATA[10] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15860_ (.D(_03945_),
    .Q(\design_top.core0.FCT3[0] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15861_ (.D(_03946_),
    .Q(\design_top.core0.FCT3[1] ),
    .CLK(clknet_5_13_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15862_ (.D(_03947_),
    .Q(\design_top.core0.FCT3[2] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15863_ (.D(_03948_),
    .Q(\design_top.core0.S1PTR[0] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15864_ (.D(_03949_),
    .Q(\design_top.core0.S1PTR[1] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15865_ (.D(_03950_),
    .Q(\design_top.core0.S1PTR[2] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15866_ (.D(_03951_),
    .Q(\design_top.core0.S1PTR[3] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15867_ (.D(_03952_),
    .Q(\design_top.core0.S2PTR[0] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15868_ (.D(_03953_),
    .Q(\design_top.core0.S2PTR[1] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15869_ (.D(_03954_),
    .Q(\design_top.core0.S2PTR[2] ),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15870_ (.D(_03955_),
    .Q(\design_top.core0.S2PTR[3] ),
    .CLK(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15871_ (.D(_03956_),
    .Q(\design_top.core0.FCT7[5] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15872_ (.D(_03957_),
    .Q(\design_top.core0.XLUI ),
    .CLK(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15873_ (.D(_03958_),
    .Q(\design_top.core0.XAUIPC ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15874_ (.D(_03959_),
    .Q(\design_top.core0.XJAL ),
    .CLK(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15875_ (.D(_03960_),
    .Q(\design_top.core0.XJALR ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15876_ (.D(_03961_),
    .Q(\design_top.core0.XBCC ),
    .CLK(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15877_ (.D(_03962_),
    .Q(\design_top.core0.XLCC ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15878_ (.D(_03963_),
    .Q(\design_top.core0.XSCC ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15879_ (.D(_03964_),
    .Q(\design_top.core0.XMCC ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15880_ (.D(_03965_),
    .Q(\design_top.core0.XRCC ),
    .CLK(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15881_ (.D(_03966_),
    .Q(\design_top.core0.SIMM[12] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15882_ (.D(_03967_),
    .Q(\design_top.core0.SIMM[13] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15883_ (.D(_03968_),
    .Q(\design_top.core0.SIMM[14] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15884_ (.D(_03969_),
    .Q(\design_top.core0.SIMM[15] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15885_ (.D(_03970_),
    .Q(\design_top.core0.SIMM[16] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15886_ (.D(_03971_),
    .Q(\design_top.core0.SIMM[17] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15887_ (.D(_03972_),
    .Q(\design_top.core0.SIMM[18] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15888_ (.D(_03973_),
    .Q(\design_top.core0.SIMM[19] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15889_ (.D(_03974_),
    .Q(\design_top.core0.SIMM[20] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15890_ (.D(_03975_),
    .Q(\design_top.core0.SIMM[21] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15891_ (.D(_03976_),
    .Q(\design_top.core0.SIMM[22] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15892_ (.D(_03977_),
    .Q(\design_top.core0.SIMM[23] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15893_ (.D(_03978_),
    .Q(\design_top.core0.SIMM[24] ),
    .CLK(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15894_ (.D(_03979_),
    .Q(\design_top.core0.SIMM[25] ),
    .CLK(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15895_ (.D(_03980_),
    .Q(\design_top.core0.SIMM[26] ),
    .CLK(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15896_ (.D(_03981_),
    .Q(\design_top.core0.SIMM[27] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15897_ (.D(_03982_),
    .Q(\design_top.core0.SIMM[28] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15898_ (.D(_03983_),
    .Q(\design_top.core0.SIMM[29] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15899_ (.D(_03984_),
    .Q(\design_top.core0.SIMM[30] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15900_ (.D(_03985_),
    .Q(\design_top.core0.SIMM[31] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15901_ (.D(_03986_),
    .Q(\design_top.core0.SIMM[0] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15902_ (.D(_03987_),
    .Q(\design_top.core0.SIMM[1] ),
    .CLK(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15903_ (.D(_03988_),
    .Q(\design_top.core0.SIMM[2] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15904_ (.D(_03989_),
    .Q(\design_top.core0.SIMM[3] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15905_ (.D(_03990_),
    .Q(\design_top.core0.SIMM[4] ),
    .CLK(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15906_ (.D(_03991_),
    .Q(\design_top.core0.SIMM[5] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15907_ (.D(_03992_),
    .Q(\design_top.core0.SIMM[6] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15908_ (.D(_03993_),
    .Q(\design_top.core0.SIMM[7] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15909_ (.D(_03994_),
    .Q(\design_top.core0.SIMM[8] ),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15910_ (.D(_03995_),
    .Q(\design_top.core0.SIMM[9] ),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15911_ (.D(_03996_),
    .Q(\design_top.core0.SIMM[10] ),
    .CLK(clknet_leaf_31_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15912_ (.D(_03997_),
    .Q(\design_top.core0.SIMM[11] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15913_ (.D(_03998_),
    .Q(\design_top.core0.UIMM[12] ),
    .CLK(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15914_ (.D(_03999_),
    .Q(\design_top.core0.UIMM[13] ),
    .CLK(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15915_ (.D(_04000_),
    .Q(\design_top.core0.UIMM[14] ),
    .CLK(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15916_ (.D(_04001_),
    .Q(\design_top.core0.UIMM[15] ),
    .CLK(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15917_ (.D(_04002_),
    .Q(\design_top.core0.UIMM[16] ),
    .CLK(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15918_ (.D(_04003_),
    .Q(\design_top.core0.UIMM[17] ),
    .CLK(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15919_ (.D(_04004_),
    .Q(\design_top.core0.UIMM[18] ),
    .CLK(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15920_ (.D(_04005_),
    .Q(\design_top.core0.UIMM[19] ),
    .CLK(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15921_ (.D(_04006_),
    .Q(\design_top.core0.UIMM[20] ),
    .CLK(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15922_ (.D(_04007_),
    .Q(\design_top.core0.UIMM[21] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15923_ (.D(_04008_),
    .Q(\design_top.core0.UIMM[22] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15924_ (.D(_04009_),
    .Q(\design_top.core0.UIMM[23] ),
    .CLK(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15925_ (.D(_04010_),
    .Q(\design_top.core0.UIMM[24] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15926_ (.D(_04011_),
    .Q(\design_top.core0.UIMM[25] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15927_ (.D(_04012_),
    .Q(\design_top.core0.UIMM[26] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15928_ (.D(_04013_),
    .Q(\design_top.core0.UIMM[27] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15929_ (.D(_04014_),
    .Q(\design_top.core0.UIMM[28] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15930_ (.D(_04015_),
    .Q(\design_top.core0.UIMM[29] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15931_ (.D(_04016_),
    .Q(\design_top.core0.UIMM[30] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15932_ (.D(_04017_),
    .Q(\design_top.core0.UIMM[31] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15933_ (.D(_04018_),
    .Q(\design_top.IOMUX[3][0] ),
    .CLK(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15934_ (.D(_04019_),
    .Q(\design_top.IOMUX[3][1] ),
    .CLK(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15935_ (.D(_04020_),
    .Q(\design_top.IOMUX[3][2] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15936_ (.D(_04021_),
    .Q(\design_top.IOMUX[3][3] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15937_ (.D(_04022_),
    .Q(\design_top.IOMUX[3][4] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15938_ (.D(_04023_),
    .Q(\design_top.IOMUX[3][5] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15939_ (.D(_04024_),
    .Q(\design_top.IOMUX[3][6] ),
    .CLK(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15940_ (.D(_04025_),
    .Q(\design_top.IOMUX[3][7] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15941_ (.D(_04026_),
    .Q(\design_top.IOMUX[3][8] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15942_ (.D(_04027_),
    .Q(\design_top.IOMUX[3][9] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15943_ (.D(_04028_),
    .Q(\design_top.IOMUX[3][10] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15944_ (.D(_04029_),
    .Q(\design_top.IOMUX[3][11] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15945_ (.D(_04030_),
    .Q(\design_top.IOMUX[3][12] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15946_ (.D(_04031_),
    .Q(\design_top.IOMUX[3][13] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15947_ (.D(_04032_),
    .Q(\design_top.IOMUX[3][14] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15948_ (.D(_04033_),
    .Q(\design_top.IOMUX[3][15] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15949_ (.D(_04034_),
    .Q(\design_top.IOMUX[3][16] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15950_ (.D(_04035_),
    .Q(\design_top.IOMUX[3][17] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15951_ (.D(_04036_),
    .Q(\design_top.IOMUX[3][18] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15952_ (.D(_04037_),
    .Q(\design_top.IOMUX[3][19] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15953_ (.D(_04038_),
    .Q(\design_top.IOMUX[3][20] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15954_ (.D(_04039_),
    .Q(\design_top.IOMUX[3][21] ),
    .CLK(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15955_ (.D(_04040_),
    .Q(\design_top.IOMUX[3][22] ),
    .CLK(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15956_ (.D(_04041_),
    .Q(\design_top.IOMUX[3][23] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15957_ (.D(_04042_),
    .Q(\design_top.IOMUX[3][24] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15958_ (.D(_04043_),
    .Q(\design_top.IOMUX[3][25] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15959_ (.D(_04044_),
    .Q(\design_top.IOMUX[3][26] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15960_ (.D(_04045_),
    .Q(\design_top.IOMUX[3][27] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15961_ (.D(_04046_),
    .Q(\design_top.IOMUX[3][28] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15962_ (.D(_04047_),
    .Q(\design_top.IOMUX[3][29] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15963_ (.D(_04048_),
    .Q(\design_top.IOMUX[3][30] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15964_ (.D(_04049_),
    .Q(\design_top.IOMUX[3][31] ),
    .CLK(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15965_ (.D(_04050_),
    .Q(\design_top.MEM[13][24] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15966_ (.D(_04051_),
    .Q(\design_top.MEM[13][25] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15967_ (.D(_04052_),
    .Q(\design_top.MEM[13][26] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15968_ (.D(_04053_),
    .Q(\design_top.MEM[13][27] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15969_ (.D(_04054_),
    .Q(\design_top.MEM[13][28] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15970_ (.D(_04055_),
    .Q(\design_top.MEM[13][29] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15971_ (.D(_04056_),
    .Q(\design_top.MEM[13][30] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15972_ (.D(_04057_),
    .Q(\design_top.MEM[13][31] ),
    .CLK(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15973_ (.D(_04058_),
    .Q(\design_top.MEM[9][16] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15974_ (.D(_04059_),
    .Q(\design_top.MEM[9][17] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15975_ (.D(_04060_),
    .Q(\design_top.MEM[9][18] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15976_ (.D(_04061_),
    .Q(\design_top.MEM[9][19] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15977_ (.D(_04062_),
    .Q(\design_top.MEM[9][20] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15978_ (.D(_04063_),
    .Q(\design_top.MEM[9][21] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15979_ (.D(_04064_),
    .Q(\design_top.MEM[9][22] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15980_ (.D(_04065_),
    .Q(\design_top.MEM[9][23] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15981_ (.D(_04066_),
    .Q(\design_top.MEM[9][8] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15982_ (.D(_04067_),
    .Q(\design_top.MEM[9][9] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15983_ (.D(_04068_),
    .Q(\design_top.MEM[9][10] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15984_ (.D(_04069_),
    .Q(\design_top.MEM[9][11] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15985_ (.D(_04070_),
    .Q(\design_top.MEM[9][12] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15986_ (.D(_04071_),
    .Q(\design_top.MEM[9][13] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15987_ (.D(_04072_),
    .Q(\design_top.MEM[9][14] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15988_ (.D(_04073_),
    .Q(\design_top.MEM[9][15] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15989_ (.D(_04074_),
    .Q(\design_top.MEM[8][24] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15990_ (.D(_04075_),
    .Q(\design_top.MEM[8][25] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15991_ (.D(_04076_),
    .Q(\design_top.MEM[8][26] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15992_ (.D(_04077_),
    .Q(\design_top.MEM[8][27] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15993_ (.D(_04078_),
    .Q(\design_top.MEM[8][28] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15994_ (.D(_04079_),
    .Q(\design_top.MEM[8][29] ),
    .CLK(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15995_ (.D(_04080_),
    .Q(\design_top.MEM[8][30] ),
    .CLK(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15996_ (.D(_04081_),
    .Q(\design_top.MEM[8][31] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15997_ (.D(_04082_),
    .Q(\design_top.MEM[8][16] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15998_ (.D(_04083_),
    .Q(\design_top.MEM[8][17] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _15999_ (.D(_04084_),
    .Q(\design_top.MEM[8][18] ),
    .CLK(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16000_ (.D(_04085_),
    .Q(\design_top.MEM[8][19] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16001_ (.D(_04086_),
    .Q(\design_top.MEM[8][20] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16002_ (.D(_04087_),
    .Q(\design_top.MEM[8][21] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16003_ (.D(_04088_),
    .Q(\design_top.MEM[8][22] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16004_ (.D(_04089_),
    .Q(\design_top.MEM[8][23] ),
    .CLK(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16005_ (.D(_04090_),
    .Q(\design_top.MEM[8][8] ),
    .CLK(clknet_leaf_235_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16006_ (.D(_04091_),
    .Q(\design_top.MEM[8][9] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16007_ (.D(_04092_),
    .Q(\design_top.MEM[8][10] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16008_ (.D(_04093_),
    .Q(\design_top.MEM[8][11] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16009_ (.D(_04094_),
    .Q(\design_top.MEM[8][12] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16010_ (.D(_04095_),
    .Q(\design_top.MEM[8][13] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16011_ (.D(_04096_),
    .Q(\design_top.MEM[8][14] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16012_ (.D(_04097_),
    .Q(\design_top.MEM[8][15] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16013_ (.D(_04098_),
    .Q(\design_top.MEM[7][24] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16014_ (.D(_04099_),
    .Q(\design_top.MEM[7][25] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16015_ (.D(_04100_),
    .Q(\design_top.MEM[7][26] ),
    .CLK(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16016_ (.D(_04101_),
    .Q(\design_top.MEM[7][27] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16017_ (.D(_04102_),
    .Q(\design_top.MEM[7][28] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16018_ (.D(_04103_),
    .Q(\design_top.MEM[7][29] ),
    .CLK(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16019_ (.D(_04104_),
    .Q(\design_top.MEM[7][30] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16020_ (.D(_04105_),
    .Q(\design_top.MEM[7][31] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16021_ (.D(_04106_),
    .Q(\design_top.MEM[7][16] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16022_ (.D(_04107_),
    .Q(\design_top.MEM[7][17] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16023_ (.D(_04108_),
    .Q(\design_top.MEM[7][18] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16024_ (.D(_04109_),
    .Q(\design_top.MEM[7][19] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16025_ (.D(_04110_),
    .Q(\design_top.MEM[7][20] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16026_ (.D(_04111_),
    .Q(\design_top.MEM[7][21] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16027_ (.D(_04112_),
    .Q(\design_top.MEM[7][22] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16028_ (.D(_04113_),
    .Q(\design_top.MEM[7][23] ),
    .CLK(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16029_ (.D(_04114_),
    .Q(\design_top.MEM[7][8] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16030_ (.D(_04115_),
    .Q(\design_top.MEM[7][9] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16031_ (.D(_04116_),
    .Q(\design_top.MEM[7][10] ),
    .CLK(clknet_leaf_235_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16032_ (.D(_04117_),
    .Q(\design_top.MEM[7][11] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16033_ (.D(_04118_),
    .Q(\design_top.MEM[7][12] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16034_ (.D(_04119_),
    .Q(\design_top.MEM[7][13] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16035_ (.D(_04120_),
    .Q(\design_top.MEM[7][14] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16036_ (.D(_04121_),
    .Q(\design_top.MEM[7][15] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16037_ (.D(_04122_),
    .Q(\design_top.MEM[6][24] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16038_ (.D(_04123_),
    .Q(\design_top.MEM[6][25] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16039_ (.D(_04124_),
    .Q(\design_top.MEM[6][26] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16040_ (.D(_04125_),
    .Q(\design_top.MEM[6][27] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16041_ (.D(_04126_),
    .Q(\design_top.MEM[6][28] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16042_ (.D(_04127_),
    .Q(\design_top.MEM[6][29] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16043_ (.D(_04128_),
    .Q(\design_top.MEM[6][30] ),
    .CLK(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16044_ (.D(_04129_),
    .Q(\design_top.MEM[6][31] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16045_ (.D(_04130_),
    .Q(\design_top.MEM[6][16] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16046_ (.D(_04131_),
    .Q(\design_top.MEM[6][17] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16047_ (.D(_04132_),
    .Q(\design_top.MEM[6][18] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16048_ (.D(_04133_),
    .Q(\design_top.MEM[6][19] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16049_ (.D(_04134_),
    .Q(\design_top.MEM[6][20] ),
    .CLK(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16050_ (.D(_04135_),
    .Q(\design_top.MEM[6][21] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16051_ (.D(_04136_),
    .Q(\design_top.MEM[6][22] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16052_ (.D(_04137_),
    .Q(\design_top.MEM[6][23] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16053_ (.D(_04138_),
    .Q(\design_top.MEM[6][8] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16054_ (.D(_04139_),
    .Q(\design_top.MEM[6][9] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16055_ (.D(_04140_),
    .Q(\design_top.MEM[6][10] ),
    .CLK(clknet_leaf_235_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16056_ (.D(_04141_),
    .Q(\design_top.MEM[6][11] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16057_ (.D(_04142_),
    .Q(\design_top.MEM[6][12] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16058_ (.D(_04143_),
    .Q(\design_top.MEM[6][13] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16059_ (.D(_04144_),
    .Q(\design_top.MEM[6][14] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16060_ (.D(_04145_),
    .Q(\design_top.MEM[6][15] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16061_ (.D(_04146_),
    .Q(\design_top.MEM[5][24] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16062_ (.D(_04147_),
    .Q(\design_top.MEM[5][25] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16063_ (.D(_04148_),
    .Q(\design_top.MEM[5][26] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16064_ (.D(_04149_),
    .Q(\design_top.MEM[5][27] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16065_ (.D(_04150_),
    .Q(\design_top.MEM[5][28] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16066_ (.D(_04151_),
    .Q(\design_top.MEM[5][29] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16067_ (.D(_04152_),
    .Q(\design_top.MEM[5][30] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16068_ (.D(_04153_),
    .Q(\design_top.MEM[5][31] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16069_ (.D(_04154_),
    .Q(\design_top.MEM[5][16] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16070_ (.D(_04155_),
    .Q(\design_top.MEM[5][17] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16071_ (.D(_04156_),
    .Q(\design_top.MEM[5][18] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16072_ (.D(_04157_),
    .Q(\design_top.MEM[5][19] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16073_ (.D(_04158_),
    .Q(\design_top.MEM[5][20] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16074_ (.D(_04159_),
    .Q(\design_top.MEM[5][21] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16075_ (.D(_04160_),
    .Q(\design_top.MEM[5][22] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16076_ (.D(_04161_),
    .Q(\design_top.MEM[5][23] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16077_ (.D(_04162_),
    .Q(\design_top.MEM[5][8] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16078_ (.D(_04163_),
    .Q(\design_top.MEM[5][9] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16079_ (.D(_04164_),
    .Q(\design_top.MEM[5][10] ),
    .CLK(clknet_leaf_235_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16080_ (.D(_04165_),
    .Q(\design_top.MEM[5][11] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16081_ (.D(_04166_),
    .Q(\design_top.MEM[5][12] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16082_ (.D(_04167_),
    .Q(\design_top.MEM[5][13] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16083_ (.D(_04168_),
    .Q(\design_top.MEM[5][14] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16084_ (.D(_04169_),
    .Q(\design_top.MEM[5][15] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16085_ (.D(_04170_),
    .Q(\design_top.MEM[4][24] ),
    .CLK(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16086_ (.D(_04171_),
    .Q(\design_top.MEM[4][25] ),
    .CLK(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16087_ (.D(_04172_),
    .Q(\design_top.MEM[4][26] ),
    .CLK(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16088_ (.D(_04173_),
    .Q(\design_top.MEM[4][27] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16089_ (.D(_04174_),
    .Q(\design_top.MEM[4][28] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16090_ (.D(_04175_),
    .Q(\design_top.MEM[4][29] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16091_ (.D(_04176_),
    .Q(\design_top.MEM[4][30] ),
    .CLK(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16092_ (.D(_04177_),
    .Q(\design_top.MEM[4][31] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16093_ (.D(_04178_),
    .Q(\design_top.MEM[4][16] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16094_ (.D(_04179_),
    .Q(\design_top.MEM[4][17] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16095_ (.D(_04180_),
    .Q(\design_top.MEM[4][18] ),
    .CLK(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16096_ (.D(_04181_),
    .Q(\design_top.MEM[4][19] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16097_ (.D(_04182_),
    .Q(\design_top.MEM[4][20] ),
    .CLK(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16098_ (.D(_04183_),
    .Q(\design_top.MEM[4][21] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16099_ (.D(_04184_),
    .Q(\design_top.MEM[4][22] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16100_ (.D(_04185_),
    .Q(\design_top.MEM[4][23] ),
    .CLK(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16101_ (.D(_04186_),
    .Q(\design_top.MEM[4][8] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16102_ (.D(_04187_),
    .Q(\design_top.MEM[4][9] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16103_ (.D(_04188_),
    .Q(\design_top.MEM[4][10] ),
    .CLK(clknet_leaf_235_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16104_ (.D(_04189_),
    .Q(\design_top.MEM[4][11] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16105_ (.D(_04190_),
    .Q(\design_top.MEM[4][12] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16106_ (.D(_04191_),
    .Q(\design_top.MEM[4][13] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16107_ (.D(_04192_),
    .Q(\design_top.MEM[4][14] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16108_ (.D(_04193_),
    .Q(\design_top.MEM[4][15] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16109_ (.D(_04194_),
    .Q(\design_top.MEM[3][24] ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16110_ (.D(_04195_),
    .Q(\design_top.MEM[3][25] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16111_ (.D(_04196_),
    .Q(\design_top.MEM[3][26] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16112_ (.D(_04197_),
    .Q(\design_top.MEM[3][27] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16113_ (.D(_04198_),
    .Q(\design_top.MEM[3][28] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16114_ (.D(_04199_),
    .Q(\design_top.MEM[3][29] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16115_ (.D(_04200_),
    .Q(\design_top.MEM[3][30] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16116_ (.D(_04201_),
    .Q(\design_top.MEM[3][31] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16117_ (.D(_04202_),
    .Q(\design_top.MEM[3][16] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16118_ (.D(_04203_),
    .Q(\design_top.MEM[3][17] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16119_ (.D(_04204_),
    .Q(\design_top.MEM[3][18] ),
    .CLK(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16120_ (.D(_04205_),
    .Q(\design_top.MEM[3][19] ),
    .CLK(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16121_ (.D(_04206_),
    .Q(\design_top.MEM[3][20] ),
    .CLK(clknet_leaf_187_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16122_ (.D(_04207_),
    .Q(\design_top.MEM[3][21] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16123_ (.D(_04208_),
    .Q(\design_top.MEM[3][22] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16124_ (.D(_04209_),
    .Q(\design_top.MEM[3][23] ),
    .CLK(clknet_leaf_187_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16125_ (.D(_04210_),
    .Q(\design_top.MEM[3][8] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16126_ (.D(_04211_),
    .Q(\design_top.MEM[3][9] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16127_ (.D(_04212_),
    .Q(\design_top.MEM[3][10] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16128_ (.D(_04213_),
    .Q(\design_top.MEM[3][11] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16129_ (.D(_04214_),
    .Q(\design_top.MEM[3][12] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16130_ (.D(_04215_),
    .Q(\design_top.MEM[3][13] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16131_ (.D(_04216_),
    .Q(\design_top.MEM[3][14] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16132_ (.D(_04217_),
    .Q(\design_top.MEM[3][15] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16133_ (.D(_04218_),
    .Q(\design_top.MEM[2][24] ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16134_ (.D(_04219_),
    .Q(\design_top.MEM[2][25] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16135_ (.D(_04220_),
    .Q(\design_top.MEM[2][26] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16136_ (.D(_04221_),
    .Q(\design_top.MEM[2][27] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16137_ (.D(_04222_),
    .Q(\design_top.MEM[2][28] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16138_ (.D(_04223_),
    .Q(\design_top.MEM[2][29] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16139_ (.D(_04224_),
    .Q(\design_top.MEM[2][30] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16140_ (.D(_04225_),
    .Q(\design_top.MEM[2][31] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16141_ (.D(_04226_),
    .Q(\design_top.MEM[2][16] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16142_ (.D(_04227_),
    .Q(\design_top.MEM[2][17] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16143_ (.D(_04228_),
    .Q(\design_top.MEM[2][18] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16144_ (.D(_04229_),
    .Q(\design_top.MEM[2][19] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16145_ (.D(_04230_),
    .Q(\design_top.MEM[2][20] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16146_ (.D(_04231_),
    .Q(\design_top.MEM[2][21] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16147_ (.D(_04232_),
    .Q(\design_top.MEM[2][22] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16148_ (.D(_04233_),
    .Q(\design_top.MEM[2][23] ),
    .CLK(clknet_leaf_187_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16149_ (.D(_04234_),
    .Q(\design_top.MEM[2][8] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16150_ (.D(_04235_),
    .Q(\design_top.MEM[2][9] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16151_ (.D(_04236_),
    .Q(\design_top.MEM[2][10] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16152_ (.D(_04237_),
    .Q(\design_top.MEM[2][11] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16153_ (.D(_04238_),
    .Q(\design_top.MEM[2][12] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16154_ (.D(_04239_),
    .Q(\design_top.MEM[2][13] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16155_ (.D(_04240_),
    .Q(\design_top.MEM[2][14] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16156_ (.D(_04241_),
    .Q(\design_top.MEM[2][15] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16157_ (.D(_04242_),
    .Q(\design_top.MEM[1][8] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16158_ (.D(_04243_),
    .Q(\design_top.MEM[1][9] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16159_ (.D(_04244_),
    .Q(\design_top.MEM[1][10] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16160_ (.D(_04245_),
    .Q(\design_top.MEM[1][11] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16161_ (.D(_04246_),
    .Q(\design_top.MEM[1][12] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16162_ (.D(_04247_),
    .Q(\design_top.MEM[1][13] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16163_ (.D(_04248_),
    .Q(\design_top.MEM[1][14] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16164_ (.D(_04249_),
    .Q(\design_top.MEM[1][15] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16165_ (.D(_04250_),
    .Q(\design_top.MEM[1][24] ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16166_ (.D(_04251_),
    .Q(\design_top.MEM[1][25] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16167_ (.D(_04252_),
    .Q(\design_top.MEM[1][26] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16168_ (.D(_04253_),
    .Q(\design_top.MEM[1][27] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16169_ (.D(_04254_),
    .Q(\design_top.MEM[1][28] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16170_ (.D(_04255_),
    .Q(\design_top.MEM[1][29] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16171_ (.D(_04256_),
    .Q(\design_top.MEM[1][30] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16172_ (.D(_04257_),
    .Q(\design_top.MEM[1][31] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16173_ (.D(_04258_),
    .Q(\design_top.MEM[1][16] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16174_ (.D(_04259_),
    .Q(\design_top.MEM[1][17] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16175_ (.D(_04260_),
    .Q(\design_top.MEM[1][18] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16176_ (.D(_04261_),
    .Q(\design_top.MEM[1][19] ),
    .CLK(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16177_ (.D(_04262_),
    .Q(\design_top.MEM[1][20] ),
    .CLK(clknet_leaf_187_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16178_ (.D(_04263_),
    .Q(\design_top.MEM[1][21] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16179_ (.D(_04264_),
    .Q(\design_top.MEM[1][22] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16180_ (.D(_04265_),
    .Q(\design_top.MEM[1][23] ),
    .CLK(clknet_leaf_187_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16181_ (.D(_04266_),
    .Q(\design_top.MEM[15][24] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16182_ (.D(_04267_),
    .Q(\design_top.MEM[15][25] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16183_ (.D(_04268_),
    .Q(\design_top.MEM[15][26] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16184_ (.D(_04269_),
    .Q(\design_top.MEM[15][27] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16185_ (.D(_04270_),
    .Q(\design_top.MEM[15][28] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16186_ (.D(_04271_),
    .Q(\design_top.MEM[15][29] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16187_ (.D(_04272_),
    .Q(\design_top.MEM[15][30] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16188_ (.D(_04273_),
    .Q(\design_top.MEM[15][31] ),
    .CLK(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16189_ (.D(_04274_),
    .Q(\design_top.MEM[15][16] ),
    .CLK(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16190_ (.D(_04275_),
    .Q(\design_top.MEM[15][17] ),
    .CLK(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16191_ (.D(_04276_),
    .Q(\design_top.MEM[15][18] ),
    .CLK(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16192_ (.D(_04277_),
    .Q(\design_top.MEM[15][19] ),
    .CLK(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16193_ (.D(_04278_),
    .Q(\design_top.MEM[15][20] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16194_ (.D(_04279_),
    .Q(\design_top.MEM[15][21] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16195_ (.D(_04280_),
    .Q(\design_top.MEM[15][22] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16196_ (.D(_04281_),
    .Q(\design_top.MEM[15][23] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16197_ (.D(_04282_),
    .Q(\design_top.MEM[15][8] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16198_ (.D(_04283_),
    .Q(\design_top.MEM[15][9] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16199_ (.D(_04284_),
    .Q(\design_top.MEM[15][10] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16200_ (.D(_04285_),
    .Q(\design_top.MEM[15][11] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16201_ (.D(_04286_),
    .Q(\design_top.MEM[15][12] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16202_ (.D(_04287_),
    .Q(\design_top.MEM[15][13] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16203_ (.D(_04288_),
    .Q(\design_top.MEM[15][14] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16204_ (.D(_04289_),
    .Q(\design_top.MEM[15][15] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16205_ (.D(_04290_),
    .Q(\design_top.MEM[13][16] ),
    .CLK(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16206_ (.D(_04291_),
    .Q(\design_top.MEM[13][17] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16207_ (.D(_04292_),
    .Q(\design_top.MEM[13][18] ),
    .CLK(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16208_ (.D(_04293_),
    .Q(\design_top.MEM[13][19] ),
    .CLK(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16209_ (.D(_04294_),
    .Q(\design_top.MEM[13][20] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16210_ (.D(_04295_),
    .Q(\design_top.MEM[13][21] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16211_ (.D(_04296_),
    .Q(\design_top.MEM[13][22] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16212_ (.D(_04297_),
    .Q(\design_top.MEM[13][23] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16213_ (.D(_04298_),
    .Q(\design_top.MEM[13][8] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16214_ (.D(_04299_),
    .Q(\design_top.MEM[13][9] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16215_ (.D(_04300_),
    .Q(\design_top.MEM[13][10] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16216_ (.D(_04301_),
    .Q(\design_top.MEM[13][11] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16217_ (.D(_04302_),
    .Q(\design_top.MEM[13][12] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16218_ (.D(_04303_),
    .Q(\design_top.MEM[13][13] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16219_ (.D(_04304_),
    .Q(\design_top.MEM[13][14] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16220_ (.D(_04305_),
    .Q(\design_top.MEM[13][15] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16221_ (.D(_04306_),
    .Q(\design_top.MEM[12][24] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16222_ (.D(_04307_),
    .Q(\design_top.MEM[12][25] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16223_ (.D(_04308_),
    .Q(\design_top.MEM[12][26] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16224_ (.D(_04309_),
    .Q(\design_top.MEM[12][27] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16225_ (.D(_04310_),
    .Q(\design_top.MEM[12][28] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16226_ (.D(_04311_),
    .Q(\design_top.MEM[12][29] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16227_ (.D(_04312_),
    .Q(\design_top.MEM[12][30] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16228_ (.D(_04313_),
    .Q(\design_top.MEM[12][31] ),
    .CLK(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16229_ (.D(_04314_),
    .Q(\design_top.MEM[12][16] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16230_ (.D(_04315_),
    .Q(\design_top.MEM[12][17] ),
    .CLK(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16231_ (.D(_04316_),
    .Q(\design_top.MEM[12][18] ),
    .CLK(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16232_ (.D(_04317_),
    .Q(\design_top.MEM[12][19] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16233_ (.D(_04318_),
    .Q(\design_top.MEM[12][20] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16234_ (.D(_04319_),
    .Q(\design_top.MEM[12][21] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16235_ (.D(_04320_),
    .Q(\design_top.MEM[12][22] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16236_ (.D(_04321_),
    .Q(\design_top.MEM[12][23] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16237_ (.D(_04322_),
    .Q(\design_top.IREQ[7] ),
    .CLK(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16238_ (.D(_04323_),
    .Q(\design_top.IACK[7] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16239_ (.D(_04324_),
    .Q(\design_top.MEM[12][8] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16240_ (.D(_04325_),
    .Q(\design_top.MEM[12][9] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16241_ (.D(_04326_),
    .Q(\design_top.MEM[12][10] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16242_ (.D(_04327_),
    .Q(\design_top.MEM[12][11] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16243_ (.D(_04328_),
    .Q(\design_top.MEM[12][12] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16244_ (.D(_04329_),
    .Q(\design_top.MEM[12][13] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16245_ (.D(_04330_),
    .Q(\design_top.MEM[12][14] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16246_ (.D(_04331_),
    .Q(\design_top.MEM[12][15] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16247_ (.D(_04332_),
    .Q(\design_top.MEM[11][8] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16248_ (.D(_04333_),
    .Q(\design_top.MEM[11][9] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16249_ (.D(_04334_),
    .Q(\design_top.MEM[11][10] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16250_ (.D(_04335_),
    .Q(\design_top.MEM[11][11] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16251_ (.D(_04336_),
    .Q(\design_top.MEM[11][12] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16252_ (.D(_04337_),
    .Q(\design_top.MEM[11][13] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16253_ (.D(_04338_),
    .Q(\design_top.MEM[11][14] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16254_ (.D(_04339_),
    .Q(\design_top.MEM[11][15] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16255_ (.D(_04340_),
    .Q(\design_top.MEM[11][24] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16256_ (.D(_04341_),
    .Q(\design_top.MEM[11][25] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16257_ (.D(_04342_),
    .Q(\design_top.MEM[11][26] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16258_ (.D(_04343_),
    .Q(\design_top.MEM[11][27] ),
    .CLK(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16259_ (.D(_04344_),
    .Q(\design_top.MEM[11][28] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16260_ (.D(_04345_),
    .Q(\design_top.MEM[11][29] ),
    .CLK(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16261_ (.D(_04346_),
    .Q(\design_top.MEM[11][30] ),
    .CLK(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16262_ (.D(_04347_),
    .Q(\design_top.MEM[11][31] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16263_ (.D(_04348_),
    .Q(\design_top.MEM[11][16] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16264_ (.D(_04349_),
    .Q(\design_top.MEM[11][17] ),
    .CLK(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16265_ (.D(_04350_),
    .Q(\design_top.MEM[11][18] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16266_ (.D(_04351_),
    .Q(\design_top.MEM[11][19] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16267_ (.D(_04352_),
    .Q(\design_top.MEM[11][20] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16268_ (.D(_04353_),
    .Q(\design_top.MEM[11][21] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16269_ (.D(_04354_),
    .Q(\design_top.MEM[11][22] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16270_ (.D(_04355_),
    .Q(\design_top.MEM[11][23] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16271_ (.D(_04356_),
    .Q(\design_top.MEM[10][24] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16272_ (.D(_04357_),
    .Q(\design_top.MEM[10][25] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16273_ (.D(_04358_),
    .Q(\design_top.MEM[10][26] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16274_ (.D(_04359_),
    .Q(\design_top.MEM[10][27] ),
    .CLK(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16275_ (.D(_04360_),
    .Q(\design_top.MEM[10][28] ),
    .CLK(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16276_ (.D(_04361_),
    .Q(\design_top.MEM[10][29] ),
    .CLK(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16277_ (.D(_04362_),
    .Q(\design_top.MEM[10][30] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16278_ (.D(_04363_),
    .Q(\design_top.MEM[10][31] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16279_ (.D(_04364_),
    .Q(\design_top.MEM[10][16] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16280_ (.D(_04365_),
    .Q(\design_top.MEM[10][17] ),
    .CLK(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16281_ (.D(_04366_),
    .Q(\design_top.MEM[10][18] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16282_ (.D(_04367_),
    .Q(\design_top.MEM[10][19] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16283_ (.D(_04368_),
    .Q(\design_top.MEM[10][20] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16284_ (.D(_04369_),
    .Q(\design_top.MEM[10][21] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16285_ (.D(_04370_),
    .Q(\design_top.MEM[10][22] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16286_ (.D(_04371_),
    .Q(\design_top.MEM[10][23] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16287_ (.D(_04372_),
    .Q(\design_top.MEM[10][8] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16288_ (.D(_04373_),
    .Q(\design_top.MEM[10][9] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16289_ (.D(_04374_),
    .Q(\design_top.MEM[10][10] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16290_ (.D(_04375_),
    .Q(\design_top.MEM[10][11] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16291_ (.D(_04376_),
    .Q(\design_top.MEM[10][12] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16292_ (.D(_04377_),
    .Q(\design_top.MEM[10][13] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16293_ (.D(_04378_),
    .Q(\design_top.MEM[10][14] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16294_ (.D(_04379_),
    .Q(\design_top.MEM[10][15] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16295_ (.D(_04380_),
    .Q(\design_top.MEM[0][8] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16296_ (.D(_04381_),
    .Q(\design_top.MEM[0][9] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16297_ (.D(_04382_),
    .Q(\design_top.MEM[0][10] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16298_ (.D(_04383_),
    .Q(\design_top.MEM[0][11] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16299_ (.D(_04384_),
    .Q(\design_top.MEM[0][12] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16300_ (.D(_04385_),
    .Q(\design_top.MEM[0][13] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16301_ (.D(_04386_),
    .Q(\design_top.MEM[0][14] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16302_ (.D(_04387_),
    .Q(\design_top.MEM[0][15] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16303_ (.D(_04388_),
    .Q(\design_top.MEM[0][16] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16304_ (.D(_04389_),
    .Q(\design_top.MEM[0][17] ),
    .CLK(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16305_ (.D(_04390_),
    .Q(\design_top.MEM[0][18] ),
    .CLK(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16306_ (.D(_04391_),
    .Q(\design_top.MEM[0][19] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16307_ (.D(_04392_),
    .Q(\design_top.MEM[0][20] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16308_ (.D(_04393_),
    .Q(\design_top.MEM[0][21] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16309_ (.D(_04394_),
    .Q(\design_top.MEM[0][22] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16310_ (.D(_04395_),
    .Q(\design_top.MEM[0][23] ),
    .CLK(clknet_leaf_187_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16311_ (.D(_04396_),
    .Q(\design_top.MEM[0][24] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16312_ (.D(_04397_),
    .Q(\design_top.MEM[0][25] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16313_ (.D(_04398_),
    .Q(\design_top.MEM[0][26] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16314_ (.D(_04399_),
    .Q(\design_top.MEM[0][27] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16315_ (.D(_04400_),
    .Q(\design_top.MEM[0][28] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16316_ (.D(_04401_),
    .Q(\design_top.MEM[0][29] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16317_ (.D(_04402_),
    .Q(\design_top.MEM[0][30] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16318_ (.D(_04403_),
    .Q(\design_top.MEM[0][31] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16319_ (.D(_04404_),
    .Q(\design_top.MEM[14][16] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16320_ (.D(_04405_),
    .Q(\design_top.MEM[14][17] ),
    .CLK(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16321_ (.D(_04406_),
    .Q(\design_top.MEM[14][18] ),
    .CLK(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16322_ (.D(_04407_),
    .Q(\design_top.MEM[14][19] ),
    .CLK(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16323_ (.D(_04408_),
    .Q(\design_top.MEM[14][20] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16324_ (.D(_04409_),
    .Q(\design_top.MEM[14][21] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16325_ (.D(_04410_),
    .Q(\design_top.MEM[14][22] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16326_ (.D(_04411_),
    .Q(\design_top.MEM[14][23] ),
    .CLK(clknet_leaf_187_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16327_ (.D(_04412_),
    .Q(\design_top.MEM[14][24] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16328_ (.D(_04413_),
    .Q(\design_top.MEM[14][25] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16329_ (.D(_04414_),
    .Q(\design_top.MEM[14][26] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16330_ (.D(_04415_),
    .Q(\design_top.MEM[14][27] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16331_ (.D(_04416_),
    .Q(\design_top.MEM[14][28] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16332_ (.D(_04417_),
    .Q(\design_top.MEM[14][29] ),
    .CLK(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16333_ (.D(_04418_),
    .Q(\design_top.MEM[14][30] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16334_ (.D(_04419_),
    .Q(\design_top.MEM[14][31] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16335_ (.D(_04420_),
    .Q(\design_top.MEM[14][8] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16336_ (.D(_04421_),
    .Q(\design_top.MEM[14][9] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16337_ (.D(_04422_),
    .Q(\design_top.MEM[14][10] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16338_ (.D(_04423_),
    .Q(\design_top.MEM[14][11] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16339_ (.D(_04424_),
    .Q(\design_top.MEM[14][12] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16340_ (.D(_04425_),
    .Q(\design_top.MEM[14][13] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16341_ (.D(_04426_),
    .Q(\design_top.MEM[14][14] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16342_ (.D(_04427_),
    .Q(\design_top.MEM[14][15] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16343_ (.D(_04428_),
    .Q(\design_top.MEM[9][24] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16344_ (.D(_04429_),
    .Q(\design_top.MEM[9][25] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16345_ (.D(_04430_),
    .Q(\design_top.MEM[9][26] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16346_ (.D(_04431_),
    .Q(\design_top.MEM[9][27] ),
    .CLK(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16347_ (.D(_04432_),
    .Q(\design_top.MEM[9][28] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16348_ (.D(_04433_),
    .Q(\design_top.MEM[9][29] ),
    .CLK(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16349_ (.D(_04434_),
    .Q(\design_top.MEM[9][30] ),
    .CLK(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16350_ (.D(_04435_),
    .Q(\design_top.MEM[9][31] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16351_ (.D(_04436_),
    .Q(io_out[16]),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _16352_ (.D(_04437_),
    .Q(io_out[17]),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_29_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_user_clock2 (.A(clknet_opt_1_user_clock2),
    .X(clknet_leaf_31_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_37_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_39_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_48_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_76_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_79_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_84_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_user_clock2 (.A(clknet_opt_3_user_clock2),
    .X(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_user_clock2 (.A(clknet_opt_5_user_clock2),
    .X(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_user_clock2 (.A(clknet_opt_6_user_clock2),
    .X(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_user_clock2 (.A(clknet_opt_4_user_clock2),
    .X(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_user_clock2 (.A(clknet_opt_2_user_clock2),
    .X(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_143_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_user_clock2 (.A(clknet_opt_0_user_clock2),
    .X(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_user_clock2 (.A(clknet_5_14_0_user_clock2),
    .X(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_user_clock2 (.A(clknet_5_14_0_user_clock2),
    .X(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_user_clock2 (.A(clknet_5_14_0_user_clock2),
    .X(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_user_clock2 (.A(clknet_5_14_0_user_clock2),
    .X(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_user_clock2 (.A(clknet_5_14_0_user_clock2),
    .X(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_172_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_user_clock2 (.A(clknet_5_14_0_user_clock2),
    .X(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_187_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_193_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_194_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_195_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_196_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_197_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_198_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_199_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_200_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_201_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_202_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_203_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_204_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_205_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_206_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_207_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_208_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_209_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_210_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_211_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_212_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_213_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_214_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_215_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_216_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_217_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_218_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_219_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_220_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_221_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_222_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_223_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_224_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_225_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_226_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_227_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_228_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_229_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_230_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_231_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_232_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_233_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_234_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_235_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_235_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_236_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_237_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_238_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_239_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_240_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_241_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_242_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_243_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_user_clock2 (.A(user_clock2),
    .X(clknet_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_0_user_clock2 (.A(clknet_0_user_clock2),
    .X(clknet_1_0_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_1_user_clock2 (.A(clknet_1_0_0_user_clock2),
    .X(clknet_1_0_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_0_user_clock2 (.A(clknet_0_user_clock2),
    .X(clknet_1_1_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_1_user_clock2 (.A(clknet_1_1_0_user_clock2),
    .X(clknet_1_1_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_0_0_user_clock2 (.A(clknet_1_0_1_user_clock2),
    .X(clknet_2_0_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_0_1_user_clock2 (.A(clknet_2_0_0_user_clock2),
    .X(clknet_2_0_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_1_0_user_clock2 (.A(clknet_1_0_1_user_clock2),
    .X(clknet_2_1_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_1_1_user_clock2 (.A(clknet_2_1_0_user_clock2),
    .X(clknet_2_1_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_2_0_user_clock2 (.A(clknet_1_1_1_user_clock2),
    .X(clknet_2_2_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_2_1_user_clock2 (.A(clknet_2_2_0_user_clock2),
    .X(clknet_2_2_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_3_0_user_clock2 (.A(clknet_1_1_1_user_clock2),
    .X(clknet_2_3_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_3_1_user_clock2 (.A(clknet_2_3_0_user_clock2),
    .X(clknet_2_3_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_0_0_user_clock2 (.A(clknet_2_0_1_user_clock2),
    .X(clknet_3_0_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_1_0_user_clock2 (.A(clknet_2_0_1_user_clock2),
    .X(clknet_3_1_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_2_0_user_clock2 (.A(clknet_2_1_1_user_clock2),
    .X(clknet_3_2_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_3_0_user_clock2 (.A(clknet_2_1_1_user_clock2),
    .X(clknet_3_3_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_4_0_user_clock2 (.A(clknet_2_2_1_user_clock2),
    .X(clknet_3_4_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_5_0_user_clock2 (.A(clknet_2_2_1_user_clock2),
    .X(clknet_3_5_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_6_0_user_clock2 (.A(clknet_2_3_1_user_clock2),
    .X(clknet_3_6_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_7_0_user_clock2 (.A(clknet_2_3_1_user_clock2),
    .X(clknet_3_7_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_0_0_user_clock2 (.A(clknet_3_0_0_user_clock2),
    .X(clknet_4_0_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_1_0_user_clock2 (.A(clknet_3_0_0_user_clock2),
    .X(clknet_4_1_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_2_0_user_clock2 (.A(clknet_3_1_0_user_clock2),
    .X(clknet_4_2_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_3_0_user_clock2 (.A(clknet_3_1_0_user_clock2),
    .X(clknet_4_3_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_4_0_user_clock2 (.A(clknet_3_2_0_user_clock2),
    .X(clknet_4_4_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_5_0_user_clock2 (.A(clknet_3_2_0_user_clock2),
    .X(clknet_4_5_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_6_0_user_clock2 (.A(clknet_3_3_0_user_clock2),
    .X(clknet_4_6_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_7_0_user_clock2 (.A(clknet_3_3_0_user_clock2),
    .X(clknet_4_7_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_8_0_user_clock2 (.A(clknet_3_4_0_user_clock2),
    .X(clknet_4_8_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_9_0_user_clock2 (.A(clknet_3_4_0_user_clock2),
    .X(clknet_4_9_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_10_0_user_clock2 (.A(clknet_3_5_0_user_clock2),
    .X(clknet_4_10_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_11_0_user_clock2 (.A(clknet_3_5_0_user_clock2),
    .X(clknet_4_11_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_12_0_user_clock2 (.A(clknet_3_6_0_user_clock2),
    .X(clknet_4_12_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_13_0_user_clock2 (.A(clknet_3_6_0_user_clock2),
    .X(clknet_4_13_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_14_0_user_clock2 (.A(clknet_3_7_0_user_clock2),
    .X(clknet_4_14_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_15_0_user_clock2 (.A(clknet_3_7_0_user_clock2),
    .X(clknet_4_15_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_0_0_user_clock2 (.A(clknet_4_0_0_user_clock2),
    .X(clknet_5_0_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_1_0_user_clock2 (.A(clknet_4_0_0_user_clock2),
    .X(clknet_5_1_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_2_0_user_clock2 (.A(clknet_4_1_0_user_clock2),
    .X(clknet_5_2_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_3_0_user_clock2 (.A(clknet_4_1_0_user_clock2),
    .X(clknet_5_3_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_4_0_user_clock2 (.A(clknet_4_2_0_user_clock2),
    .X(clknet_5_4_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_5_0_user_clock2 (.A(clknet_4_2_0_user_clock2),
    .X(clknet_5_5_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_6_0_user_clock2 (.A(clknet_4_3_0_user_clock2),
    .X(clknet_5_6_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_7_0_user_clock2 (.A(clknet_4_3_0_user_clock2),
    .X(clknet_5_7_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_8_0_user_clock2 (.A(clknet_4_4_0_user_clock2),
    .X(clknet_5_8_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_9_0_user_clock2 (.A(clknet_4_4_0_user_clock2),
    .X(clknet_5_9_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_10_0_user_clock2 (.A(clknet_4_5_0_user_clock2),
    .X(clknet_5_10_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_11_0_user_clock2 (.A(clknet_4_5_0_user_clock2),
    .X(clknet_5_11_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_12_0_user_clock2 (.A(clknet_4_6_0_user_clock2),
    .X(clknet_5_12_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_13_0_user_clock2 (.A(clknet_4_6_0_user_clock2),
    .X(clknet_5_13_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_14_0_user_clock2 (.A(clknet_4_7_0_user_clock2),
    .X(clknet_5_14_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_15_0_user_clock2 (.A(clknet_4_7_0_user_clock2),
    .X(clknet_5_15_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_16_0_user_clock2 (.A(clknet_4_8_0_user_clock2),
    .X(clknet_5_16_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_17_0_user_clock2 (.A(clknet_4_8_0_user_clock2),
    .X(clknet_5_17_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_18_0_user_clock2 (.A(clknet_4_9_0_user_clock2),
    .X(clknet_5_18_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_19_0_user_clock2 (.A(clknet_4_9_0_user_clock2),
    .X(clknet_5_19_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_20_0_user_clock2 (.A(clknet_4_10_0_user_clock2),
    .X(clknet_5_20_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_21_0_user_clock2 (.A(clknet_4_10_0_user_clock2),
    .X(clknet_5_21_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_22_0_user_clock2 (.A(clknet_4_11_0_user_clock2),
    .X(clknet_5_22_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_23_0_user_clock2 (.A(clknet_4_11_0_user_clock2),
    .X(clknet_5_23_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_24_0_user_clock2 (.A(clknet_4_12_0_user_clock2),
    .X(clknet_5_24_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_25_0_user_clock2 (.A(clknet_4_12_0_user_clock2),
    .X(clknet_5_25_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_26_0_user_clock2 (.A(clknet_4_13_0_user_clock2),
    .X(clknet_5_26_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_27_0_user_clock2 (.A(clknet_4_13_0_user_clock2),
    .X(clknet_5_27_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_28_0_user_clock2 (.A(clknet_4_14_0_user_clock2),
    .X(clknet_5_28_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_29_0_user_clock2 (.A(clknet_4_14_0_user_clock2),
    .X(clknet_5_29_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_30_0_user_clock2 (.A(clknet_4_15_0_user_clock2),
    .X(clknet_5_30_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_31_0_user_clock2 (.A(clknet_4_15_0_user_clock2),
    .X(clknet_5_31_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_0_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_opt_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_opt_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_opt_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_3_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_opt_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_4_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_opt_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_5_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_opt_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_6_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_opt_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
endmodule
