magic
tech sky130A
magscale 1 2
timestamp 1622195742
<< obsli1 >>
rect 1225 2261 120307 121091
<< obsm1 >>
rect 1104 2128 121058 121440
<< metal2 >>
rect 478 123200 534 124000
rect 938 123200 994 124000
rect 1858 123200 1914 124000
rect 2318 123200 2374 124000
rect 2778 123200 2834 124000
rect 3698 123200 3754 124000
rect 4158 123200 4214 124000
rect 4618 123200 4674 124000
rect 5538 123200 5594 124000
rect 5998 123200 6054 124000
rect 6918 123200 6974 124000
rect 7378 123200 7434 124000
rect 7838 123200 7894 124000
rect 8758 123200 8814 124000
rect 9218 123200 9274 124000
rect 10138 123200 10194 124000
rect 10598 123200 10654 124000
rect 11058 123200 11114 124000
rect 11978 123200 12034 124000
rect 12438 123200 12494 124000
rect 13358 123200 13414 124000
rect 13818 123200 13874 124000
rect 14278 123200 14334 124000
rect 15198 123200 15254 124000
rect 15658 123200 15714 124000
rect 16578 123200 16634 124000
rect 17038 123200 17094 124000
rect 17498 123200 17554 124000
rect 18418 123200 18474 124000
rect 18878 123200 18934 124000
rect 19798 123200 19854 124000
rect 20258 123200 20314 124000
rect 20718 123200 20774 124000
rect 21638 123200 21694 124000
rect 22098 123200 22154 124000
rect 23018 123200 23074 124000
rect 23478 123200 23534 124000
rect 23938 123200 23994 124000
rect 24858 123200 24914 124000
rect 25318 123200 25374 124000
rect 25778 123200 25834 124000
rect 26698 123200 26754 124000
rect 27158 123200 27214 124000
rect 28078 123200 28134 124000
rect 28538 123200 28594 124000
rect 28998 123200 29054 124000
rect 29918 123200 29974 124000
rect 30378 123200 30434 124000
rect 31298 123200 31354 124000
rect 31758 123200 31814 124000
rect 32218 123200 32274 124000
rect 33138 123200 33194 124000
rect 33598 123200 33654 124000
rect 34518 123200 34574 124000
rect 34978 123200 35034 124000
rect 35438 123200 35494 124000
rect 36358 123200 36414 124000
rect 36818 123200 36874 124000
rect 37738 123200 37794 124000
rect 38198 123200 38254 124000
rect 38658 123200 38714 124000
rect 39578 123200 39634 124000
rect 40038 123200 40094 124000
rect 40958 123200 41014 124000
rect 41418 123200 41474 124000
rect 41878 123200 41934 124000
rect 42798 123200 42854 124000
rect 43258 123200 43314 124000
rect 44178 123200 44234 124000
rect 44638 123200 44694 124000
rect 45098 123200 45154 124000
rect 46018 123200 46074 124000
rect 46478 123200 46534 124000
rect 46938 123200 46994 124000
rect 47858 123200 47914 124000
rect 48318 123200 48374 124000
rect 49238 123200 49294 124000
rect 49698 123200 49754 124000
rect 50158 123200 50214 124000
rect 51078 123200 51134 124000
rect 51538 123200 51594 124000
rect 52458 123200 52514 124000
rect 52918 123200 52974 124000
rect 53378 123200 53434 124000
rect 54298 123200 54354 124000
rect 54758 123200 54814 124000
rect 55678 123200 55734 124000
rect 56138 123200 56194 124000
rect 56598 123200 56654 124000
rect 57518 123200 57574 124000
rect 57978 123200 58034 124000
rect 58898 123200 58954 124000
rect 59358 123200 59414 124000
rect 59818 123200 59874 124000
rect 60738 123200 60794 124000
rect 61198 123200 61254 124000
rect 62118 123200 62174 124000
rect 62578 123200 62634 124000
rect 63038 123200 63094 124000
rect 63958 123200 64014 124000
rect 64418 123200 64474 124000
rect 65338 123200 65394 124000
rect 65798 123200 65854 124000
rect 66258 123200 66314 124000
rect 67178 123200 67234 124000
rect 67638 123200 67694 124000
rect 68098 123200 68154 124000
rect 69018 123200 69074 124000
rect 69478 123200 69534 124000
rect 70398 123200 70454 124000
rect 70858 123200 70914 124000
rect 71318 123200 71374 124000
rect 72238 123200 72294 124000
rect 72698 123200 72754 124000
rect 73618 123200 73674 124000
rect 74078 123200 74134 124000
rect 74538 123200 74594 124000
rect 75458 123200 75514 124000
rect 75918 123200 75974 124000
rect 76838 123200 76894 124000
rect 77298 123200 77354 124000
rect 77758 123200 77814 124000
rect 78678 123200 78734 124000
rect 79138 123200 79194 124000
rect 80058 123200 80114 124000
rect 80518 123200 80574 124000
rect 80978 123200 81034 124000
rect 81898 123200 81954 124000
rect 82358 123200 82414 124000
rect 83278 123200 83334 124000
rect 83738 123200 83794 124000
rect 84198 123200 84254 124000
rect 85118 123200 85174 124000
rect 85578 123200 85634 124000
rect 86498 123200 86554 124000
rect 86958 123200 87014 124000
rect 87418 123200 87474 124000
rect 88338 123200 88394 124000
rect 88798 123200 88854 124000
rect 89258 123200 89314 124000
rect 90178 123200 90234 124000
rect 90638 123200 90694 124000
rect 91558 123200 91614 124000
rect 92018 123200 92074 124000
rect 92478 123200 92534 124000
rect 93398 123200 93454 124000
rect 93858 123200 93914 124000
rect 94778 123200 94834 124000
rect 95238 123200 95294 124000
rect 95698 123200 95754 124000
rect 96618 123200 96674 124000
rect 97078 123200 97134 124000
rect 97998 123200 98054 124000
rect 98458 123200 98514 124000
rect 98918 123200 98974 124000
rect 99838 123200 99894 124000
rect 100298 123200 100354 124000
rect 101218 123200 101274 124000
rect 101678 123200 101734 124000
rect 102138 123200 102194 124000
rect 103058 123200 103114 124000
rect 103518 123200 103574 124000
rect 104438 123200 104494 124000
rect 104898 123200 104954 124000
rect 105358 123200 105414 124000
rect 106278 123200 106334 124000
rect 106738 123200 106794 124000
rect 107658 123200 107714 124000
rect 108118 123200 108174 124000
rect 108578 123200 108634 124000
rect 109498 123200 109554 124000
rect 109958 123200 110014 124000
rect 110418 123200 110474 124000
rect 111338 123200 111394 124000
rect 111798 123200 111854 124000
rect 112718 123200 112774 124000
rect 113178 123200 113234 124000
rect 113638 123200 113694 124000
rect 114558 123200 114614 124000
rect 115018 123200 115074 124000
rect 115938 123200 115994 124000
rect 116398 123200 116454 124000
rect 116858 123200 116914 124000
rect 117778 123200 117834 124000
rect 118238 123200 118294 124000
rect 119158 123200 119214 124000
rect 119618 123200 119674 124000
rect 120078 123200 120134 124000
rect 120998 123200 121054 124000
rect 478 0 534 800
rect 938 0 994 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3238 0 3294 800
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 7378 0 7434 800
rect 7838 0 7894 800
rect 8758 0 8814 800
rect 9218 0 9274 800
rect 9678 0 9734 800
rect 10598 0 10654 800
rect 11058 0 11114 800
rect 11978 0 12034 800
rect 12438 0 12494 800
rect 12898 0 12954 800
rect 13818 0 13874 800
rect 14278 0 14334 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 18418 0 18474 800
rect 18878 0 18934 800
rect 19338 0 19394 800
rect 20258 0 20314 800
rect 20718 0 20774 800
rect 21638 0 21694 800
rect 22098 0 22154 800
rect 22558 0 22614 800
rect 23478 0 23534 800
rect 23938 0 23994 800
rect 24398 0 24454 800
rect 25318 0 25374 800
rect 25778 0 25834 800
rect 26698 0 26754 800
rect 27158 0 27214 800
rect 27618 0 27674 800
rect 28538 0 28594 800
rect 28998 0 29054 800
rect 29918 0 29974 800
rect 30378 0 30434 800
rect 30838 0 30894 800
rect 31758 0 31814 800
rect 32218 0 32274 800
rect 33138 0 33194 800
rect 33598 0 33654 800
rect 34058 0 34114 800
rect 34978 0 35034 800
rect 35438 0 35494 800
rect 36358 0 36414 800
rect 36818 0 36874 800
rect 37278 0 37334 800
rect 38198 0 38254 800
rect 38658 0 38714 800
rect 39578 0 39634 800
rect 40038 0 40094 800
rect 40498 0 40554 800
rect 41418 0 41474 800
rect 41878 0 41934 800
rect 42798 0 42854 800
rect 43258 0 43314 800
rect 43718 0 43774 800
rect 44638 0 44694 800
rect 45098 0 45154 800
rect 45558 0 45614 800
rect 46478 0 46534 800
rect 46938 0 46994 800
rect 47858 0 47914 800
rect 48318 0 48374 800
rect 48778 0 48834 800
rect 49698 0 49754 800
rect 50158 0 50214 800
rect 51078 0 51134 800
rect 51538 0 51594 800
rect 51998 0 52054 800
rect 52918 0 52974 800
rect 53378 0 53434 800
rect 54298 0 54354 800
rect 54758 0 54814 800
rect 55218 0 55274 800
rect 56138 0 56194 800
rect 56598 0 56654 800
rect 57518 0 57574 800
rect 57978 0 58034 800
rect 58438 0 58494 800
rect 59358 0 59414 800
rect 59818 0 59874 800
rect 60738 0 60794 800
rect 61198 0 61254 800
rect 61658 0 61714 800
rect 62578 0 62634 800
rect 63038 0 63094 800
rect 63958 0 64014 800
rect 64418 0 64474 800
rect 64878 0 64934 800
rect 65798 0 65854 800
rect 66258 0 66314 800
rect 66718 0 66774 800
rect 67638 0 67694 800
rect 68098 0 68154 800
rect 69018 0 69074 800
rect 69478 0 69534 800
rect 69938 0 69994 800
rect 70858 0 70914 800
rect 71318 0 71374 800
rect 72238 0 72294 800
rect 72698 0 72754 800
rect 73158 0 73214 800
rect 74078 0 74134 800
rect 74538 0 74594 800
rect 75458 0 75514 800
rect 75918 0 75974 800
rect 76378 0 76434 800
rect 77298 0 77354 800
rect 77758 0 77814 800
rect 78678 0 78734 800
rect 79138 0 79194 800
rect 79598 0 79654 800
rect 80518 0 80574 800
rect 80978 0 81034 800
rect 81898 0 81954 800
rect 82358 0 82414 800
rect 82818 0 82874 800
rect 83738 0 83794 800
rect 84198 0 84254 800
rect 85118 0 85174 800
rect 85578 0 85634 800
rect 86038 0 86094 800
rect 86958 0 87014 800
rect 87418 0 87474 800
rect 87878 0 87934 800
rect 88798 0 88854 800
rect 89258 0 89314 800
rect 90178 0 90234 800
rect 90638 0 90694 800
rect 91098 0 91154 800
rect 92018 0 92074 800
rect 92478 0 92534 800
rect 93398 0 93454 800
rect 93858 0 93914 800
rect 94318 0 94374 800
rect 95238 0 95294 800
rect 95698 0 95754 800
rect 96618 0 96674 800
rect 97078 0 97134 800
rect 97538 0 97594 800
rect 98458 0 98514 800
rect 98918 0 98974 800
rect 99838 0 99894 800
rect 100298 0 100354 800
rect 100758 0 100814 800
rect 101678 0 101734 800
rect 102138 0 102194 800
rect 103058 0 103114 800
rect 103518 0 103574 800
rect 103978 0 104034 800
rect 104898 0 104954 800
rect 105358 0 105414 800
rect 106278 0 106334 800
rect 106738 0 106794 800
rect 107198 0 107254 800
rect 108118 0 108174 800
rect 108578 0 108634 800
rect 109038 0 109094 800
rect 109958 0 110014 800
rect 110418 0 110474 800
rect 111338 0 111394 800
rect 111798 0 111854 800
rect 112258 0 112314 800
rect 113178 0 113234 800
rect 113638 0 113694 800
rect 114558 0 114614 800
rect 115018 0 115074 800
rect 115478 0 115534 800
rect 116398 0 116454 800
rect 116858 0 116914 800
rect 117778 0 117834 800
rect 118238 0 118294 800
rect 118698 0 118754 800
rect 119618 0 119674 800
rect 120078 0 120134 800
rect 120998 0 121054 800
<< obsm2 >>
rect 1216 123144 1802 123200
rect 1970 123144 2262 123200
rect 2430 123144 2722 123200
rect 2890 123144 3642 123200
rect 3810 123144 4102 123200
rect 4270 123144 4562 123200
rect 4730 123144 5482 123200
rect 5650 123144 5942 123200
rect 6110 123144 6862 123200
rect 7030 123144 7322 123200
rect 7490 123144 7782 123200
rect 7950 123144 8702 123200
rect 8870 123144 9162 123200
rect 9330 123144 10082 123200
rect 10250 123144 10542 123200
rect 10710 123144 11002 123200
rect 11170 123144 11922 123200
rect 12090 123144 12382 123200
rect 12550 123144 13302 123200
rect 13470 123144 13762 123200
rect 13930 123144 14222 123200
rect 14390 123144 15142 123200
rect 15310 123144 15602 123200
rect 15770 123144 16522 123200
rect 16690 123144 16982 123200
rect 17150 123144 17442 123200
rect 17610 123144 18362 123200
rect 18530 123144 18822 123200
rect 18990 123144 19742 123200
rect 19910 123144 20202 123200
rect 20370 123144 20662 123200
rect 20830 123144 21582 123200
rect 21750 123144 22042 123200
rect 22210 123144 22962 123200
rect 23130 123144 23422 123200
rect 23590 123144 23882 123200
rect 24050 123144 24802 123200
rect 24970 123144 25262 123200
rect 25430 123144 25722 123200
rect 25890 123144 26642 123200
rect 26810 123144 27102 123200
rect 27270 123144 28022 123200
rect 28190 123144 28482 123200
rect 28650 123144 28942 123200
rect 29110 123144 29862 123200
rect 30030 123144 30322 123200
rect 30490 123144 31242 123200
rect 31410 123144 31702 123200
rect 31870 123144 32162 123200
rect 32330 123144 33082 123200
rect 33250 123144 33542 123200
rect 33710 123144 34462 123200
rect 34630 123144 34922 123200
rect 35090 123144 35382 123200
rect 35550 123144 36302 123200
rect 36470 123144 36762 123200
rect 36930 123144 37682 123200
rect 37850 123144 38142 123200
rect 38310 123144 38602 123200
rect 38770 123144 39522 123200
rect 39690 123144 39982 123200
rect 40150 123144 40902 123200
rect 41070 123144 41362 123200
rect 41530 123144 41822 123200
rect 41990 123144 42742 123200
rect 42910 123144 43202 123200
rect 43370 123144 44122 123200
rect 44290 123144 44582 123200
rect 44750 123144 45042 123200
rect 45210 123144 45962 123200
rect 46130 123144 46422 123200
rect 46590 123144 46882 123200
rect 47050 123144 47802 123200
rect 47970 123144 48262 123200
rect 48430 123144 49182 123200
rect 49350 123144 49642 123200
rect 49810 123144 50102 123200
rect 50270 123144 51022 123200
rect 51190 123144 51482 123200
rect 51650 123144 52402 123200
rect 52570 123144 52862 123200
rect 53030 123144 53322 123200
rect 53490 123144 54242 123200
rect 54410 123144 54702 123200
rect 54870 123144 55622 123200
rect 55790 123144 56082 123200
rect 56250 123144 56542 123200
rect 56710 123144 57462 123200
rect 57630 123144 57922 123200
rect 58090 123144 58842 123200
rect 59010 123144 59302 123200
rect 59470 123144 59762 123200
rect 59930 123144 60682 123200
rect 60850 123144 61142 123200
rect 61310 123144 62062 123200
rect 62230 123144 62522 123200
rect 62690 123144 62982 123200
rect 63150 123144 63902 123200
rect 64070 123144 64362 123200
rect 64530 123144 65282 123200
rect 65450 123144 65742 123200
rect 65910 123144 66202 123200
rect 66370 123144 67122 123200
rect 67290 123144 67582 123200
rect 67750 123144 68042 123200
rect 68210 123144 68962 123200
rect 69130 123144 69422 123200
rect 69590 123144 70342 123200
rect 70510 123144 70802 123200
rect 70970 123144 71262 123200
rect 71430 123144 72182 123200
rect 72350 123144 72642 123200
rect 72810 123144 73562 123200
rect 73730 123144 74022 123200
rect 74190 123144 74482 123200
rect 74650 123144 75402 123200
rect 75570 123144 75862 123200
rect 76030 123144 76782 123200
rect 76950 123144 77242 123200
rect 77410 123144 77702 123200
rect 77870 123144 78622 123200
rect 78790 123144 79082 123200
rect 79250 123144 80002 123200
rect 80170 123144 80462 123200
rect 80630 123144 80922 123200
rect 81090 123144 81842 123200
rect 82010 123144 82302 123200
rect 82470 123144 83222 123200
rect 83390 123144 83682 123200
rect 83850 123144 84142 123200
rect 84310 123144 85062 123200
rect 85230 123144 85522 123200
rect 85690 123144 86442 123200
rect 86610 123144 86902 123200
rect 87070 123144 87362 123200
rect 87530 123144 88282 123200
rect 88450 123144 88742 123200
rect 88910 123144 89202 123200
rect 89370 123144 90122 123200
rect 90290 123144 90582 123200
rect 90750 123144 91502 123200
rect 91670 123144 91962 123200
rect 92130 123144 92422 123200
rect 92590 123144 93342 123200
rect 93510 123144 93802 123200
rect 93970 123144 94722 123200
rect 94890 123144 95182 123200
rect 95350 123144 95642 123200
rect 95810 123144 96562 123200
rect 96730 123144 97022 123200
rect 97190 123144 97942 123200
rect 98110 123144 98402 123200
rect 98570 123144 98862 123200
rect 99030 123144 99782 123200
rect 99950 123144 100242 123200
rect 100410 123144 101162 123200
rect 101330 123144 101622 123200
rect 101790 123144 102082 123200
rect 102250 123144 103002 123200
rect 103170 123144 103462 123200
rect 103630 123144 104382 123200
rect 104550 123144 104842 123200
rect 105010 123144 105302 123200
rect 105470 123144 106222 123200
rect 106390 123144 106682 123200
rect 106850 123144 107602 123200
rect 107770 123144 108062 123200
rect 108230 123144 108522 123200
rect 108690 123144 109442 123200
rect 109610 123144 109902 123200
rect 110070 123144 110362 123200
rect 110530 123144 111282 123200
rect 111450 123144 111742 123200
rect 111910 123144 112662 123200
rect 112830 123144 113122 123200
rect 113290 123144 113582 123200
rect 113750 123144 114502 123200
rect 114670 123144 114962 123200
rect 115130 123144 115882 123200
rect 116050 123144 116342 123200
rect 116510 123144 116802 123200
rect 116970 123144 117722 123200
rect 117890 123144 118182 123200
rect 118350 123144 119102 123200
rect 119270 123144 119562 123200
rect 119730 123144 120022 123200
rect 120190 123144 120942 123200
rect 1216 856 121052 123144
rect 1216 711 1342 856
rect 1510 711 2262 856
rect 2430 711 2722 856
rect 2890 711 3182 856
rect 3350 711 4102 856
rect 4270 711 4562 856
rect 4730 711 5482 856
rect 5650 711 5942 856
rect 6110 711 6402 856
rect 6570 711 7322 856
rect 7490 711 7782 856
rect 7950 711 8702 856
rect 8870 711 9162 856
rect 9330 711 9622 856
rect 9790 711 10542 856
rect 10710 711 11002 856
rect 11170 711 11922 856
rect 12090 711 12382 856
rect 12550 711 12842 856
rect 13010 711 13762 856
rect 13930 711 14222 856
rect 14390 711 15142 856
rect 15310 711 15602 856
rect 15770 711 16062 856
rect 16230 711 16982 856
rect 17150 711 17442 856
rect 17610 711 18362 856
rect 18530 711 18822 856
rect 18990 711 19282 856
rect 19450 711 20202 856
rect 20370 711 20662 856
rect 20830 711 21582 856
rect 21750 711 22042 856
rect 22210 711 22502 856
rect 22670 711 23422 856
rect 23590 711 23882 856
rect 24050 711 24342 856
rect 24510 711 25262 856
rect 25430 711 25722 856
rect 25890 711 26642 856
rect 26810 711 27102 856
rect 27270 711 27562 856
rect 27730 711 28482 856
rect 28650 711 28942 856
rect 29110 711 29862 856
rect 30030 711 30322 856
rect 30490 711 30782 856
rect 30950 711 31702 856
rect 31870 711 32162 856
rect 32330 711 33082 856
rect 33250 711 33542 856
rect 33710 711 34002 856
rect 34170 711 34922 856
rect 35090 711 35382 856
rect 35550 711 36302 856
rect 36470 711 36762 856
rect 36930 711 37222 856
rect 37390 711 38142 856
rect 38310 711 38602 856
rect 38770 711 39522 856
rect 39690 711 39982 856
rect 40150 711 40442 856
rect 40610 711 41362 856
rect 41530 711 41822 856
rect 41990 711 42742 856
rect 42910 711 43202 856
rect 43370 711 43662 856
rect 43830 711 44582 856
rect 44750 711 45042 856
rect 45210 711 45502 856
rect 45670 711 46422 856
rect 46590 711 46882 856
rect 47050 711 47802 856
rect 47970 711 48262 856
rect 48430 711 48722 856
rect 48890 711 49642 856
rect 49810 711 50102 856
rect 50270 711 51022 856
rect 51190 711 51482 856
rect 51650 711 51942 856
rect 52110 711 52862 856
rect 53030 711 53322 856
rect 53490 711 54242 856
rect 54410 711 54702 856
rect 54870 711 55162 856
rect 55330 711 56082 856
rect 56250 711 56542 856
rect 56710 711 57462 856
rect 57630 711 57922 856
rect 58090 711 58382 856
rect 58550 711 59302 856
rect 59470 711 59762 856
rect 59930 711 60682 856
rect 60850 711 61142 856
rect 61310 711 61602 856
rect 61770 711 62522 856
rect 62690 711 62982 856
rect 63150 711 63902 856
rect 64070 711 64362 856
rect 64530 711 64822 856
rect 64990 711 65742 856
rect 65910 711 66202 856
rect 66370 711 66662 856
rect 66830 711 67582 856
rect 67750 711 68042 856
rect 68210 711 68962 856
rect 69130 711 69422 856
rect 69590 711 69882 856
rect 70050 711 70802 856
rect 70970 711 71262 856
rect 71430 711 72182 856
rect 72350 711 72642 856
rect 72810 711 73102 856
rect 73270 711 74022 856
rect 74190 711 74482 856
rect 74650 711 75402 856
rect 75570 711 75862 856
rect 76030 711 76322 856
rect 76490 711 77242 856
rect 77410 711 77702 856
rect 77870 711 78622 856
rect 78790 711 79082 856
rect 79250 711 79542 856
rect 79710 711 80462 856
rect 80630 711 80922 856
rect 81090 711 81842 856
rect 82010 711 82302 856
rect 82470 711 82762 856
rect 82930 711 83682 856
rect 83850 711 84142 856
rect 84310 711 85062 856
rect 85230 711 85522 856
rect 85690 711 85982 856
rect 86150 711 86902 856
rect 87070 711 87362 856
rect 87530 711 87822 856
rect 87990 711 88742 856
rect 88910 711 89202 856
rect 89370 711 90122 856
rect 90290 711 90582 856
rect 90750 711 91042 856
rect 91210 711 91962 856
rect 92130 711 92422 856
rect 92590 711 93342 856
rect 93510 711 93802 856
rect 93970 711 94262 856
rect 94430 711 95182 856
rect 95350 711 95642 856
rect 95810 711 96562 856
rect 96730 711 97022 856
rect 97190 711 97482 856
rect 97650 711 98402 856
rect 98570 711 98862 856
rect 99030 711 99782 856
rect 99950 711 100242 856
rect 100410 711 100702 856
rect 100870 711 101622 856
rect 101790 711 102082 856
rect 102250 711 103002 856
rect 103170 711 103462 856
rect 103630 711 103922 856
rect 104090 711 104842 856
rect 105010 711 105302 856
rect 105470 711 106222 856
rect 106390 711 106682 856
rect 106850 711 107142 856
rect 107310 711 108062 856
rect 108230 711 108522 856
rect 108690 711 108982 856
rect 109150 711 109902 856
rect 110070 711 110362 856
rect 110530 711 111282 856
rect 111450 711 111742 856
rect 111910 711 112202 856
rect 112370 711 113122 856
rect 113290 711 113582 856
rect 113750 711 114502 856
rect 114670 711 114962 856
rect 115130 711 115422 856
rect 115590 711 116342 856
rect 116510 711 116802 856
rect 116970 711 117722 856
rect 117890 711 118182 856
rect 118350 711 118642 856
rect 118810 711 119562 856
rect 119730 711 120022 856
rect 120190 711 120942 856
<< metal3 >>
rect 121056 123088 121856 123208
rect 0 122408 800 122528
rect 0 121728 800 121848
rect 121056 121728 121856 121848
rect 0 121048 800 121168
rect 121056 121048 121856 121168
rect 121056 120368 121856 120488
rect 0 119688 800 119808
rect 0 119008 800 119128
rect 121056 119008 121856 119128
rect 121056 118328 121856 118448
rect 0 117648 800 117768
rect 0 116968 800 117088
rect 121056 116968 121856 117088
rect 0 116288 800 116408
rect 121056 116288 121856 116408
rect 121056 115608 121856 115728
rect 0 114928 800 115048
rect 0 114248 800 114368
rect 121056 114248 121856 114368
rect 121056 113568 121856 113688
rect 0 112888 800 113008
rect 0 112208 800 112328
rect 121056 112208 121856 112328
rect 0 111528 800 111648
rect 121056 111528 121856 111648
rect 121056 110848 121856 110968
rect 0 110168 800 110288
rect 0 109488 800 109608
rect 121056 109488 121856 109608
rect 121056 108808 121856 108928
rect 0 108128 800 108248
rect 0 107448 800 107568
rect 121056 107448 121856 107568
rect 0 106768 800 106888
rect 121056 106768 121856 106888
rect 121056 106088 121856 106208
rect 0 105408 800 105528
rect 0 104728 800 104848
rect 121056 104728 121856 104848
rect 121056 104048 121856 104168
rect 0 103368 800 103488
rect 121056 103368 121856 103488
rect 0 102688 800 102808
rect 0 102008 800 102128
rect 121056 102008 121856 102128
rect 121056 101328 121856 101448
rect 0 100648 800 100768
rect 0 99968 800 100088
rect 121056 99968 121856 100088
rect 121056 99288 121856 99408
rect 0 98608 800 98728
rect 121056 98608 121856 98728
rect 0 97928 800 98048
rect 0 97248 800 97368
rect 121056 97248 121856 97368
rect 121056 96568 121856 96688
rect 0 95888 800 96008
rect 0 95208 800 95328
rect 121056 95208 121856 95328
rect 0 94528 800 94648
rect 121056 94528 121856 94648
rect 121056 93848 121856 93968
rect 0 93168 800 93288
rect 0 92488 800 92608
rect 121056 92488 121856 92608
rect 121056 91808 121856 91928
rect 0 91128 800 91248
rect 0 90448 800 90568
rect 121056 90448 121856 90568
rect 0 89768 800 89888
rect 121056 89768 121856 89888
rect 121056 89088 121856 89208
rect 0 88408 800 88528
rect 0 87728 800 87848
rect 121056 87728 121856 87848
rect 121056 87048 121856 87168
rect 0 86368 800 86488
rect 0 85688 800 85808
rect 121056 85688 121856 85808
rect 0 85008 800 85128
rect 121056 85008 121856 85128
rect 121056 84328 121856 84448
rect 0 83648 800 83768
rect 0 82968 800 83088
rect 121056 82968 121856 83088
rect 121056 82288 121856 82408
rect 0 81608 800 81728
rect 0 80928 800 81048
rect 121056 80928 121856 81048
rect 0 80248 800 80368
rect 121056 80248 121856 80368
rect 121056 79568 121856 79688
rect 0 78888 800 79008
rect 0 78208 800 78328
rect 121056 78208 121856 78328
rect 121056 77528 121856 77648
rect 0 76848 800 76968
rect 0 76168 800 76288
rect 121056 76168 121856 76288
rect 0 75488 800 75608
rect 121056 75488 121856 75608
rect 121056 74808 121856 74928
rect 0 74128 800 74248
rect 0 73448 800 73568
rect 121056 73448 121856 73568
rect 121056 72768 121856 72888
rect 0 72088 800 72208
rect 121056 72088 121856 72208
rect 0 71408 800 71528
rect 0 70728 800 70848
rect 121056 70728 121856 70848
rect 121056 70048 121856 70168
rect 0 69368 800 69488
rect 0 68688 800 68808
rect 121056 68688 121856 68808
rect 121056 68008 121856 68128
rect 0 67328 800 67448
rect 121056 67328 121856 67448
rect 0 66648 800 66768
rect 0 65968 800 66088
rect 121056 65968 121856 66088
rect 121056 65288 121856 65408
rect 0 64608 800 64728
rect 0 63928 800 64048
rect 121056 63928 121856 64048
rect 0 63248 800 63368
rect 121056 63248 121856 63368
rect 121056 62568 121856 62688
rect 0 61888 800 62008
rect 0 61208 800 61328
rect 121056 61208 121856 61328
rect 121056 60528 121856 60648
rect 0 59848 800 59968
rect 0 59168 800 59288
rect 121056 59168 121856 59288
rect 0 58488 800 58608
rect 121056 58488 121856 58608
rect 121056 57808 121856 57928
rect 0 57128 800 57248
rect 0 56448 800 56568
rect 121056 56448 121856 56568
rect 121056 55768 121856 55888
rect 0 55088 800 55208
rect 0 54408 800 54528
rect 121056 54408 121856 54528
rect 0 53728 800 53848
rect 121056 53728 121856 53848
rect 121056 53048 121856 53168
rect 0 52368 800 52488
rect 0 51688 800 51808
rect 121056 51688 121856 51808
rect 121056 51008 121856 51128
rect 0 50328 800 50448
rect 0 49648 800 49768
rect 121056 49648 121856 49768
rect 0 48968 800 49088
rect 121056 48968 121856 49088
rect 121056 48288 121856 48408
rect 0 47608 800 47728
rect 0 46928 800 47048
rect 121056 46928 121856 47048
rect 121056 46248 121856 46368
rect 0 45568 800 45688
rect 0 44888 800 45008
rect 121056 44888 121856 45008
rect 0 44208 800 44328
rect 121056 44208 121856 44328
rect 121056 43528 121856 43648
rect 0 42848 800 42968
rect 0 42168 800 42288
rect 121056 42168 121856 42288
rect 121056 41488 121856 41608
rect 0 40808 800 40928
rect 121056 40808 121856 40928
rect 0 40128 800 40248
rect 0 39448 800 39568
rect 121056 39448 121856 39568
rect 121056 38768 121856 38888
rect 0 38088 800 38208
rect 0 37408 800 37528
rect 121056 37408 121856 37528
rect 121056 36728 121856 36848
rect 0 36048 800 36168
rect 121056 36048 121856 36168
rect 0 35368 800 35488
rect 0 34688 800 34808
rect 121056 34688 121856 34808
rect 121056 34008 121856 34128
rect 0 33328 800 33448
rect 0 32648 800 32768
rect 121056 32648 121856 32768
rect 0 31968 800 32088
rect 121056 31968 121856 32088
rect 121056 31288 121856 31408
rect 0 30608 800 30728
rect 0 29928 800 30048
rect 121056 29928 121856 30048
rect 121056 29248 121856 29368
rect 0 28568 800 28688
rect 0 27888 800 28008
rect 121056 27888 121856 28008
rect 0 27208 800 27328
rect 121056 27208 121856 27328
rect 121056 26528 121856 26648
rect 0 25848 800 25968
rect 0 25168 800 25288
rect 121056 25168 121856 25288
rect 121056 24488 121856 24608
rect 0 23808 800 23928
rect 0 23128 800 23248
rect 121056 23128 121856 23248
rect 0 22448 800 22568
rect 121056 22448 121856 22568
rect 121056 21768 121856 21888
rect 0 21088 800 21208
rect 0 20408 800 20528
rect 121056 20408 121856 20528
rect 121056 19728 121856 19848
rect 0 19048 800 19168
rect 0 18368 800 18488
rect 121056 18368 121856 18488
rect 0 17688 800 17808
rect 121056 17688 121856 17808
rect 121056 17008 121856 17128
rect 0 16328 800 16448
rect 0 15648 800 15768
rect 121056 15648 121856 15768
rect 121056 14968 121856 15088
rect 0 14288 800 14408
rect 0 13608 800 13728
rect 121056 13608 121856 13728
rect 0 12928 800 13048
rect 121056 12928 121856 13048
rect 121056 12248 121856 12368
rect 0 11568 800 11688
rect 0 10888 800 11008
rect 121056 10888 121856 11008
rect 121056 10208 121856 10328
rect 0 9528 800 9648
rect 121056 9528 121856 9648
rect 0 8848 800 8968
rect 0 8168 800 8288
rect 121056 8168 121856 8288
rect 121056 7488 121856 7608
rect 0 6808 800 6928
rect 0 6128 800 6248
rect 121056 6128 121856 6248
rect 121056 5448 121856 5568
rect 0 4768 800 4888
rect 121056 4768 121856 4888
rect 0 4088 800 4208
rect 0 3408 800 3528
rect 121056 3408 121856 3528
rect 121056 2728 121856 2848
rect 0 2048 800 2168
rect 0 1368 800 1488
rect 121056 1368 121856 1488
rect 121056 688 121856 808
<< obsm3 >>
rect 800 123008 120976 123181
rect 800 122608 121056 123008
rect 880 122328 121056 122608
rect 800 121928 121056 122328
rect 880 121648 120976 121928
rect 800 121248 121056 121648
rect 880 120968 120976 121248
rect 800 120568 121056 120968
rect 800 120288 120976 120568
rect 800 119888 121056 120288
rect 880 119608 121056 119888
rect 800 119208 121056 119608
rect 880 118928 120976 119208
rect 800 118528 121056 118928
rect 800 118248 120976 118528
rect 800 117848 121056 118248
rect 880 117568 121056 117848
rect 800 117168 121056 117568
rect 880 116888 120976 117168
rect 800 116488 121056 116888
rect 880 116208 120976 116488
rect 800 115808 121056 116208
rect 800 115528 120976 115808
rect 800 115128 121056 115528
rect 880 114848 121056 115128
rect 800 114448 121056 114848
rect 880 114168 120976 114448
rect 800 113768 121056 114168
rect 800 113488 120976 113768
rect 800 113088 121056 113488
rect 880 112808 121056 113088
rect 800 112408 121056 112808
rect 880 112128 120976 112408
rect 800 111728 121056 112128
rect 880 111448 120976 111728
rect 800 111048 121056 111448
rect 800 110768 120976 111048
rect 800 110368 121056 110768
rect 880 110088 121056 110368
rect 800 109688 121056 110088
rect 880 109408 120976 109688
rect 800 109008 121056 109408
rect 800 108728 120976 109008
rect 800 108328 121056 108728
rect 880 108048 121056 108328
rect 800 107648 121056 108048
rect 880 107368 120976 107648
rect 800 106968 121056 107368
rect 880 106688 120976 106968
rect 800 106288 121056 106688
rect 800 106008 120976 106288
rect 800 105608 121056 106008
rect 880 105328 121056 105608
rect 800 104928 121056 105328
rect 880 104648 120976 104928
rect 800 104248 121056 104648
rect 800 103968 120976 104248
rect 800 103568 121056 103968
rect 880 103288 120976 103568
rect 800 102888 121056 103288
rect 880 102608 121056 102888
rect 800 102208 121056 102608
rect 880 101928 120976 102208
rect 800 101528 121056 101928
rect 800 101248 120976 101528
rect 800 100848 121056 101248
rect 880 100568 121056 100848
rect 800 100168 121056 100568
rect 880 99888 120976 100168
rect 800 99488 121056 99888
rect 800 99208 120976 99488
rect 800 98808 121056 99208
rect 880 98528 120976 98808
rect 800 98128 121056 98528
rect 880 97848 121056 98128
rect 800 97448 121056 97848
rect 880 97168 120976 97448
rect 800 96768 121056 97168
rect 800 96488 120976 96768
rect 800 96088 121056 96488
rect 880 95808 121056 96088
rect 800 95408 121056 95808
rect 880 95128 120976 95408
rect 800 94728 121056 95128
rect 880 94448 120976 94728
rect 800 94048 121056 94448
rect 800 93768 120976 94048
rect 800 93368 121056 93768
rect 880 93088 121056 93368
rect 800 92688 121056 93088
rect 880 92408 120976 92688
rect 800 92008 121056 92408
rect 800 91728 120976 92008
rect 800 91328 121056 91728
rect 880 91048 121056 91328
rect 800 90648 121056 91048
rect 880 90368 120976 90648
rect 800 89968 121056 90368
rect 880 89688 120976 89968
rect 800 89288 121056 89688
rect 800 89008 120976 89288
rect 800 88608 121056 89008
rect 880 88328 121056 88608
rect 800 87928 121056 88328
rect 880 87648 120976 87928
rect 800 87248 121056 87648
rect 800 86968 120976 87248
rect 800 86568 121056 86968
rect 880 86288 121056 86568
rect 800 85888 121056 86288
rect 880 85608 120976 85888
rect 800 85208 121056 85608
rect 880 84928 120976 85208
rect 800 84528 121056 84928
rect 800 84248 120976 84528
rect 800 83848 121056 84248
rect 880 83568 121056 83848
rect 800 83168 121056 83568
rect 880 82888 120976 83168
rect 800 82488 121056 82888
rect 800 82208 120976 82488
rect 800 81808 121056 82208
rect 880 81528 121056 81808
rect 800 81128 121056 81528
rect 880 80848 120976 81128
rect 800 80448 121056 80848
rect 880 80168 120976 80448
rect 800 79768 121056 80168
rect 800 79488 120976 79768
rect 800 79088 121056 79488
rect 880 78808 121056 79088
rect 800 78408 121056 78808
rect 880 78128 120976 78408
rect 800 77728 121056 78128
rect 800 77448 120976 77728
rect 800 77048 121056 77448
rect 880 76768 121056 77048
rect 800 76368 121056 76768
rect 880 76088 120976 76368
rect 800 75688 121056 76088
rect 880 75408 120976 75688
rect 800 75008 121056 75408
rect 800 74728 120976 75008
rect 800 74328 121056 74728
rect 880 74048 121056 74328
rect 800 73648 121056 74048
rect 880 73368 120976 73648
rect 800 72968 121056 73368
rect 800 72688 120976 72968
rect 800 72288 121056 72688
rect 880 72008 120976 72288
rect 800 71608 121056 72008
rect 880 71328 121056 71608
rect 800 70928 121056 71328
rect 880 70648 120976 70928
rect 800 70248 121056 70648
rect 800 69968 120976 70248
rect 800 69568 121056 69968
rect 880 69288 121056 69568
rect 800 68888 121056 69288
rect 880 68608 120976 68888
rect 800 68208 121056 68608
rect 800 67928 120976 68208
rect 800 67528 121056 67928
rect 880 67248 120976 67528
rect 800 66848 121056 67248
rect 880 66568 121056 66848
rect 800 66168 121056 66568
rect 880 65888 120976 66168
rect 800 65488 121056 65888
rect 800 65208 120976 65488
rect 800 64808 121056 65208
rect 880 64528 121056 64808
rect 800 64128 121056 64528
rect 880 63848 120976 64128
rect 800 63448 121056 63848
rect 880 63168 120976 63448
rect 800 62768 121056 63168
rect 800 62488 120976 62768
rect 800 62088 121056 62488
rect 880 61808 121056 62088
rect 800 61408 121056 61808
rect 880 61128 120976 61408
rect 800 60728 121056 61128
rect 800 60448 120976 60728
rect 800 60048 121056 60448
rect 880 59768 121056 60048
rect 800 59368 121056 59768
rect 880 59088 120976 59368
rect 800 58688 121056 59088
rect 880 58408 120976 58688
rect 800 58008 121056 58408
rect 800 57728 120976 58008
rect 800 57328 121056 57728
rect 880 57048 121056 57328
rect 800 56648 121056 57048
rect 880 56368 120976 56648
rect 800 55968 121056 56368
rect 800 55688 120976 55968
rect 800 55288 121056 55688
rect 880 55008 121056 55288
rect 800 54608 121056 55008
rect 880 54328 120976 54608
rect 800 53928 121056 54328
rect 880 53648 120976 53928
rect 800 53248 121056 53648
rect 800 52968 120976 53248
rect 800 52568 121056 52968
rect 880 52288 121056 52568
rect 800 51888 121056 52288
rect 880 51608 120976 51888
rect 800 51208 121056 51608
rect 800 50928 120976 51208
rect 800 50528 121056 50928
rect 880 50248 121056 50528
rect 800 49848 121056 50248
rect 880 49568 120976 49848
rect 800 49168 121056 49568
rect 880 48888 120976 49168
rect 800 48488 121056 48888
rect 800 48208 120976 48488
rect 800 47808 121056 48208
rect 880 47528 121056 47808
rect 800 47128 121056 47528
rect 880 46848 120976 47128
rect 800 46448 121056 46848
rect 800 46168 120976 46448
rect 800 45768 121056 46168
rect 880 45488 121056 45768
rect 800 45088 121056 45488
rect 880 44808 120976 45088
rect 800 44408 121056 44808
rect 880 44128 120976 44408
rect 800 43728 121056 44128
rect 800 43448 120976 43728
rect 800 43048 121056 43448
rect 880 42768 121056 43048
rect 800 42368 121056 42768
rect 880 42088 120976 42368
rect 800 41688 121056 42088
rect 800 41408 120976 41688
rect 800 41008 121056 41408
rect 880 40728 120976 41008
rect 800 40328 121056 40728
rect 880 40048 121056 40328
rect 800 39648 121056 40048
rect 880 39368 120976 39648
rect 800 38968 121056 39368
rect 800 38688 120976 38968
rect 800 38288 121056 38688
rect 880 38008 121056 38288
rect 800 37608 121056 38008
rect 880 37328 120976 37608
rect 800 36928 121056 37328
rect 800 36648 120976 36928
rect 800 36248 121056 36648
rect 880 35968 120976 36248
rect 800 35568 121056 35968
rect 880 35288 121056 35568
rect 800 34888 121056 35288
rect 880 34608 120976 34888
rect 800 34208 121056 34608
rect 800 33928 120976 34208
rect 800 33528 121056 33928
rect 880 33248 121056 33528
rect 800 32848 121056 33248
rect 880 32568 120976 32848
rect 800 32168 121056 32568
rect 880 31888 120976 32168
rect 800 31488 121056 31888
rect 800 31208 120976 31488
rect 800 30808 121056 31208
rect 880 30528 121056 30808
rect 800 30128 121056 30528
rect 880 29848 120976 30128
rect 800 29448 121056 29848
rect 800 29168 120976 29448
rect 800 28768 121056 29168
rect 880 28488 121056 28768
rect 800 28088 121056 28488
rect 880 27808 120976 28088
rect 800 27408 121056 27808
rect 880 27128 120976 27408
rect 800 26728 121056 27128
rect 800 26448 120976 26728
rect 800 26048 121056 26448
rect 880 25768 121056 26048
rect 800 25368 121056 25768
rect 880 25088 120976 25368
rect 800 24688 121056 25088
rect 800 24408 120976 24688
rect 800 24008 121056 24408
rect 880 23728 121056 24008
rect 800 23328 121056 23728
rect 880 23048 120976 23328
rect 800 22648 121056 23048
rect 880 22368 120976 22648
rect 800 21968 121056 22368
rect 800 21688 120976 21968
rect 800 21288 121056 21688
rect 880 21008 121056 21288
rect 800 20608 121056 21008
rect 880 20328 120976 20608
rect 800 19928 121056 20328
rect 800 19648 120976 19928
rect 800 19248 121056 19648
rect 880 18968 121056 19248
rect 800 18568 121056 18968
rect 880 18288 120976 18568
rect 800 17888 121056 18288
rect 880 17608 120976 17888
rect 800 17208 121056 17608
rect 800 16928 120976 17208
rect 800 16528 121056 16928
rect 880 16248 121056 16528
rect 800 15848 121056 16248
rect 880 15568 120976 15848
rect 800 15168 121056 15568
rect 800 14888 120976 15168
rect 800 14488 121056 14888
rect 880 14208 121056 14488
rect 800 13808 121056 14208
rect 880 13528 120976 13808
rect 800 13128 121056 13528
rect 880 12848 120976 13128
rect 800 12448 121056 12848
rect 800 12168 120976 12448
rect 800 11768 121056 12168
rect 880 11488 121056 11768
rect 800 11088 121056 11488
rect 880 10808 120976 11088
rect 800 10408 121056 10808
rect 800 10128 120976 10408
rect 800 9728 121056 10128
rect 880 9448 120976 9728
rect 800 9048 121056 9448
rect 880 8768 121056 9048
rect 800 8368 121056 8768
rect 880 8088 120976 8368
rect 800 7688 121056 8088
rect 800 7408 120976 7688
rect 800 7008 121056 7408
rect 880 6728 121056 7008
rect 800 6328 121056 6728
rect 880 6048 120976 6328
rect 800 5648 121056 6048
rect 800 5368 120976 5648
rect 800 4968 121056 5368
rect 880 4688 120976 4968
rect 800 4288 121056 4688
rect 880 4008 121056 4288
rect 800 3608 121056 4008
rect 880 3328 120976 3608
rect 800 2928 121056 3328
rect 800 2648 120976 2928
rect 800 2248 121056 2648
rect 880 1968 121056 2248
rect 800 1568 121056 1968
rect 880 1288 120976 1568
rect 800 888 121056 1288
rect 800 715 120976 888
<< metal4 >>
rect -8576 -7504 -7976 130992
rect -7636 -6564 -7036 130052
rect -6696 -5624 -6096 129112
rect -5756 -4684 -5156 128172
rect -4816 -3744 -4216 127232
rect -3876 -2804 -3276 126292
rect -2936 -1864 -2336 125352
rect -1996 -924 -1396 124412
rect 804 -1864 1404 125352
rect 4404 -3744 5004 127232
rect 8004 -5624 8604 129112
rect 11604 -7504 12204 130992
rect 18804 -1864 19404 125352
rect 22404 -3744 23004 127232
rect 26004 -5624 26604 129112
rect 29604 -7504 30204 130992
rect 36804 -1864 37404 125352
rect 40404 -3744 41004 127232
rect 44004 -5624 44604 129112
rect 47604 -7504 48204 130992
rect 54804 -1864 55404 125352
rect 58404 -3744 59004 127232
rect 62004 -5624 62604 129112
rect 65604 -7504 66204 130992
rect 72804 -1864 73404 125352
rect 76404 -3744 77004 127232
rect 80004 -5624 80604 129112
rect 83604 -7504 84204 130992
rect 90804 -1864 91404 125352
rect 94404 -3744 95004 127232
rect 98004 -5624 98604 129112
rect 101604 -7504 102204 130992
rect 108804 -1864 109404 125352
rect 112404 -3744 113004 127232
rect 116004 -5624 116604 129112
rect 119604 -7504 120204 130992
rect 123204 -924 123804 124412
rect 124144 -1864 124744 125352
rect 125084 -2804 125684 126292
rect 126024 -3744 126624 127232
rect 126964 -4684 127564 128172
rect 127904 -5624 128504 129112
rect 128844 -6564 129444 130052
rect 129784 -7504 130384 130992
<< obsm4 >>
rect 18091 3843 18724 120053
rect 19484 3843 22324 120053
rect 23084 3843 25924 120053
rect 26684 3843 29524 120053
rect 30284 3843 36724 120053
rect 37484 3843 40324 120053
rect 41084 3843 43924 120053
rect 44684 3843 47524 120053
rect 48284 3843 54724 120053
rect 55484 3843 58324 120053
rect 59084 3843 61924 120053
rect 62684 3843 65524 120053
rect 66284 3843 72724 120053
rect 73484 3843 76324 120053
rect 77084 3843 79924 120053
rect 80684 3843 83524 120053
rect 84284 3843 90724 120053
rect 91484 3843 94324 120053
rect 95084 3843 97924 120053
rect 98684 3843 101524 120053
rect 102284 3843 108724 120053
rect 109484 3843 112324 120053
rect 113084 3843 115924 120053
rect 116684 3843 118621 120053
<< metal5 >>
rect -8576 130392 130384 130992
rect -7636 129452 129444 130052
rect -6696 128512 128504 129112
rect -5756 127572 127564 128172
rect -4816 126632 126624 127232
rect -3876 125692 125684 126292
rect -2936 124752 124744 125352
rect -1996 123812 123804 124412
rect -6696 117076 128504 117676
rect -4816 113476 126624 114076
rect -2936 109828 124744 110428
rect -8576 102676 130384 103276
rect -6696 99076 128504 99676
rect -4816 95476 126624 96076
rect -2936 91828 124744 92428
rect -8576 84676 130384 85276
rect -6696 81076 128504 81676
rect -4816 77476 126624 78076
rect -2936 73828 124744 74428
rect -8576 66676 130384 67276
rect -6696 63076 128504 63676
rect -4816 59476 126624 60076
rect -2936 55828 124744 56428
rect -8576 48676 130384 49276
rect -6696 45076 128504 45676
rect -4816 41476 126624 42076
rect -2936 37828 124744 38428
rect -8576 30676 130384 31276
rect -6696 27076 128504 27676
rect -4816 23476 126624 24076
rect -2936 19828 124744 20428
rect -8576 12676 130384 13276
rect -6696 9076 128504 9676
rect -4816 5476 126624 6076
rect -2936 1828 124744 2428
rect -1996 -924 123804 -324
rect -2936 -1864 124744 -1264
rect -3876 -2804 125684 -2204
rect -4816 -3744 126624 -3144
rect -5756 -4684 127564 -4084
rect -6696 -5624 128504 -5024
rect -7636 -6564 129444 -5964
rect -8576 -7504 130384 -6904
<< obsm5 >>
rect -8576 130992 -7976 130994
rect 29604 130992 30204 130994
rect 65604 130992 66204 130994
rect 101604 130992 102204 130994
rect 129784 130992 130384 130994
rect -8576 130390 -7976 130392
rect 29604 130390 30204 130392
rect 65604 130390 66204 130392
rect 101604 130390 102204 130392
rect 129784 130390 130384 130392
rect -7636 130052 -7036 130054
rect 11604 130052 12204 130054
rect 47604 130052 48204 130054
rect 83604 130052 84204 130054
rect 119604 130052 120204 130054
rect 128844 130052 129444 130054
rect -7636 129450 -7036 129452
rect 11604 129450 12204 129452
rect 47604 129450 48204 129452
rect 83604 129450 84204 129452
rect 119604 129450 120204 129452
rect 128844 129450 129444 129452
rect -6696 129112 -6096 129114
rect 26004 129112 26604 129114
rect 62004 129112 62604 129114
rect 98004 129112 98604 129114
rect 127904 129112 128504 129114
rect -6696 128510 -6096 128512
rect 26004 128510 26604 128512
rect 62004 128510 62604 128512
rect 98004 128510 98604 128512
rect 127904 128510 128504 128512
rect -5756 128172 -5156 128174
rect 8004 128172 8604 128174
rect 44004 128172 44604 128174
rect 80004 128172 80604 128174
rect 116004 128172 116604 128174
rect 126964 128172 127564 128174
rect -5756 127570 -5156 127572
rect 8004 127570 8604 127572
rect 44004 127570 44604 127572
rect 80004 127570 80604 127572
rect 116004 127570 116604 127572
rect 126964 127570 127564 127572
rect -4816 127232 -4216 127234
rect 22404 127232 23004 127234
rect 58404 127232 59004 127234
rect 94404 127232 95004 127234
rect 126024 127232 126624 127234
rect -4816 126630 -4216 126632
rect 22404 126630 23004 126632
rect 58404 126630 59004 126632
rect 94404 126630 95004 126632
rect 126024 126630 126624 126632
rect -3876 126292 -3276 126294
rect 4404 126292 5004 126294
rect 40404 126292 41004 126294
rect 76404 126292 77004 126294
rect 112404 126292 113004 126294
rect 125084 126292 125684 126294
rect -3876 125690 -3276 125692
rect 4404 125690 5004 125692
rect 40404 125690 41004 125692
rect 76404 125690 77004 125692
rect 112404 125690 113004 125692
rect 125084 125690 125684 125692
rect -2936 125352 -2336 125354
rect 18804 125352 19404 125354
rect 54804 125352 55404 125354
rect 90804 125352 91404 125354
rect 124144 125352 124744 125354
rect -2936 124750 -2336 124752
rect 18804 124750 19404 124752
rect 54804 124750 55404 124752
rect 90804 124750 91404 124752
rect 124144 124750 124744 124752
rect -1996 124412 -1396 124414
rect 804 124412 1404 124414
rect 36804 124412 37404 124414
rect 72804 124412 73404 124414
rect 108804 124412 109404 124414
rect 123204 124412 123804 124414
rect -1996 123810 -1396 123812
rect 123204 123810 123804 123812
rect 0 117996 121856 123492
rect -5756 117676 -5156 117678
rect 126964 117676 127564 117678
rect -5756 117074 -5156 117076
rect 126964 117074 127564 117076
rect 0 114396 121856 116756
rect -3876 114076 -3276 114078
rect 125084 114076 125684 114078
rect -3876 113474 -3276 113476
rect 125084 113474 125684 113476
rect 0 110748 121856 113156
rect -1996 110428 -1396 110430
rect 123204 110428 123804 110430
rect -1996 109826 -1396 109828
rect 123204 109826 123804 109828
rect 0 103596 121856 109508
rect -8576 103276 -7976 103278
rect 129784 103276 130384 103278
rect -8576 102674 -7976 102676
rect 129784 102674 130384 102676
rect 0 99996 121856 102356
rect -6696 99676 -6096 99678
rect 127904 99676 128504 99678
rect -6696 99074 -6096 99076
rect 127904 99074 128504 99076
rect 0 96396 121856 98756
rect -4816 96076 -4216 96078
rect 126024 96076 126624 96078
rect -4816 95474 -4216 95476
rect 126024 95474 126624 95476
rect 0 92748 121856 95156
rect -2936 92428 -2336 92430
rect 124144 92428 124744 92430
rect -2936 91826 -2336 91828
rect 124144 91826 124744 91828
rect 0 85596 121856 91508
rect -7636 85276 -7036 85278
rect 128844 85276 129444 85278
rect -7636 84674 -7036 84676
rect 128844 84674 129444 84676
rect 0 81996 121856 84356
rect -5756 81676 -5156 81678
rect 126964 81676 127564 81678
rect -5756 81074 -5156 81076
rect 126964 81074 127564 81076
rect 0 78396 121856 80756
rect -3876 78076 -3276 78078
rect 125084 78076 125684 78078
rect -3876 77474 -3276 77476
rect 125084 77474 125684 77476
rect 0 74748 121856 77156
rect -1996 74428 -1396 74430
rect 123204 74428 123804 74430
rect -1996 73826 -1396 73828
rect 123204 73826 123804 73828
rect 0 67596 121856 73508
rect -8576 67276 -7976 67278
rect 129784 67276 130384 67278
rect -8576 66674 -7976 66676
rect 129784 66674 130384 66676
rect 0 63996 121856 66356
rect -6696 63676 -6096 63678
rect 127904 63676 128504 63678
rect -6696 63074 -6096 63076
rect 127904 63074 128504 63076
rect 0 60396 121856 62756
rect -4816 60076 -4216 60078
rect 126024 60076 126624 60078
rect -4816 59474 -4216 59476
rect 126024 59474 126624 59476
rect 0 56748 121856 59156
rect -2936 56428 -2336 56430
rect 124144 56428 124744 56430
rect -2936 55826 -2336 55828
rect 124144 55826 124744 55828
rect 0 49596 121856 55508
rect -7636 49276 -7036 49278
rect 128844 49276 129444 49278
rect -7636 48674 -7036 48676
rect 128844 48674 129444 48676
rect 0 45996 121856 48356
rect -5756 45676 -5156 45678
rect 126964 45676 127564 45678
rect -5756 45074 -5156 45076
rect 126964 45074 127564 45076
rect 0 42396 121856 44756
rect -3876 42076 -3276 42078
rect 125084 42076 125684 42078
rect -3876 41474 -3276 41476
rect 125084 41474 125684 41476
rect 0 38748 121856 41156
rect -1996 38428 -1396 38430
rect 123204 38428 123804 38430
rect -1996 37826 -1396 37828
rect 123204 37826 123804 37828
rect 0 31596 121856 37508
rect -8576 31276 -7976 31278
rect 129784 31276 130384 31278
rect -8576 30674 -7976 30676
rect 129784 30674 130384 30676
rect 0 27996 121856 30356
rect -6696 27676 -6096 27678
rect 127904 27676 128504 27678
rect -6696 27074 -6096 27076
rect 127904 27074 128504 27076
rect 0 24396 121856 26756
rect -4816 24076 -4216 24078
rect 126024 24076 126624 24078
rect -4816 23474 -4216 23476
rect 126024 23474 126624 23476
rect 0 20748 121856 23156
rect -2936 20428 -2336 20430
rect 124144 20428 124744 20430
rect -2936 19826 -2336 19828
rect 124144 19826 124744 19828
rect 0 13596 121856 19508
rect -7636 13276 -7036 13278
rect 128844 13276 129444 13278
rect -7636 12674 -7036 12676
rect 128844 12674 129444 12676
rect 0 9996 121856 12356
rect -5756 9676 -5156 9678
rect 126964 9676 127564 9678
rect -5756 9074 -5156 9076
rect 126964 9074 127564 9076
rect 0 6396 121856 8756
rect -3876 6076 -3276 6078
rect 125084 6076 125684 6078
rect -3876 5474 -3276 5476
rect 125084 5474 125684 5476
rect 0 2748 121856 5156
rect -1996 2428 -1396 2430
rect 123204 2428 123804 2430
rect -1996 1826 -1396 1828
rect 123204 1826 123804 1828
rect 0 0 121856 1508
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 123204 -324 123804 -322
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 123204 -926 123804 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 124144 -1264 124744 -1262
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 124144 -1866 124744 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 125084 -2204 125684 -2202
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 125084 -2806 125684 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 126024 -3144 126624 -3142
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 126024 -3746 126624 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 126964 -4084 127564 -4082
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 126964 -4686 127564 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 127904 -5024 128504 -5022
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 127904 -5626 128504 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 128844 -5964 129444 -5962
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 128844 -6566 129444 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 129784 -6904 130384 -6902
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 129784 -7506 130384 -7504
<< labels >>
rlabel metal2 s 2778 123200 2834 124000 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 121056 95208 121856 95328 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 94318 0 94374 800 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal3 s 0 117648 800 117768 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal3 s 121056 97248 121856 97368 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 108578 0 108634 800 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal3 s 0 88408 800 88528 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 5998 0 6054 800 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 82818 0 82874 800 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal2 s 65798 0 65854 800 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 73618 123200 73674 124000 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal2 s 114558 0 114614 800 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 0 1368 800 1488 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal2 s 72238 0 72294 800 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 121056 51008 121856 51128 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 80058 123200 80114 124000 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal2 s 74538 0 74594 800 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal2 s 90638 123200 90694 124000 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal2 s 7378 0 7434 800 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 0 40128 800 40248 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 121056 80248 121856 80368 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 0 53728 800 53848 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 121056 114248 121856 114368 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal2 s 77298 0 77354 800 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 0 119008 800 119128 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal2 s 34978 0 35034 800 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal2 s 57978 0 58034 800 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 98458 123200 98514 124000 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal3 s 121056 63928 121856 64048 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal2 s 109958 0 110014 800 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 io_in[10]
port 31 nsew signal input
rlabel metal2 s 113178 123200 113234 124000 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 io_in[12]
port 33 nsew signal input
rlabel metal2 s 41878 123200 41934 124000 6 io_in[13]
port 34 nsew signal input
rlabel metal2 s 21638 123200 21694 124000 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 io_in[15]
port 36 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 io_in[16]
port 37 nsew signal input
rlabel metal3 s 121056 72768 121856 72888 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 108578 123200 108634 124000 6 io_in[18]
port 39 nsew signal input
rlabel metal3 s 121056 2728 121856 2848 6 io_in[19]
port 40 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 70858 123200 70914 124000 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 74538 123200 74594 124000 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 46018 123200 46074 124000 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 io_in[24]
port 46 nsew signal input
rlabel metal3 s 121056 58488 121856 58608 6 io_in[25]
port 47 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 io_in[26]
port 48 nsew signal input
rlabel metal2 s 31298 123200 31354 124000 6 io_in[27]
port 49 nsew signal input
rlabel metal2 s 31758 123200 31814 124000 6 io_in[28]
port 50 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 io_in[29]
port 51 nsew signal input
rlabel metal2 s 101218 123200 101274 124000 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s 121056 10888 121856 11008 6 io_in[30]
port 53 nsew signal input
rlabel metal3 s 121056 7488 121856 7608 6 io_in[31]
port 54 nsew signal input
rlabel metal2 s 9218 123200 9274 124000 6 io_in[32]
port 55 nsew signal input
rlabel metal3 s 0 122408 800 122528 6 io_in[33]
port 56 nsew signal input
rlabel metal3 s 121056 91808 121856 91928 6 io_in[34]
port 57 nsew signal input
rlabel metal2 s 118698 0 118754 800 6 io_in[35]
port 58 nsew signal input
rlabel metal2 s 56598 123200 56654 124000 6 io_in[36]
port 59 nsew signal input
rlabel metal2 s 15658 123200 15714 124000 6 io_in[37]
port 60 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 io_in[3]
port 61 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 121056 20408 121856 20528 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 0 102688 800 102808 6 io_in[6]
port 64 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 io_in[7]
port 65 nsew signal input
rlabel metal2 s 113638 123200 113694 124000 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 121056 109488 121856 109608 6 io_in[9]
port 67 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 io_oeb[0]
port 68 nsew signal output
rlabel metal2 s 112258 0 112314 800 6 io_oeb[10]
port 69 nsew signal output
rlabel metal2 s 100758 0 100814 800 6 io_oeb[11]
port 70 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 io_oeb[12]
port 71 nsew signal output
rlabel metal2 s 40038 123200 40094 124000 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 121056 70728 121856 70848 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 106278 123200 106334 124000 6 io_oeb[15]
port 74 nsew signal output
rlabel metal3 s 121056 27888 121856 28008 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 111338 123200 111394 124000 6 io_oeb[18]
port 77 nsew signal output
rlabel metal3 s 121056 46248 121856 46368 6 io_oeb[19]
port 78 nsew signal output
rlabel metal2 s 89258 0 89314 800 6 io_oeb[1]
port 79 nsew signal output
rlabel metal3 s 121056 74808 121856 74928 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 10138 123200 10194 124000 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 2318 0 2374 800 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s 121056 21768 121856 21888 6 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s 0 116288 800 116408 6 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 io_oeb[26]
port 86 nsew signal output
rlabel metal2 s 54758 123200 54814 124000 6 io_oeb[27]
port 87 nsew signal output
rlabel metal2 s 24858 123200 24914 124000 6 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 io_oeb[29]
port 89 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 io_oeb[30]
port 91 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 io_oeb[31]
port 92 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s 121056 17688 121856 17808 6 io_oeb[33]
port 94 nsew signal output
rlabel metal2 s 35438 123200 35494 124000 6 io_oeb[34]
port 95 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 io_oeb[36]
port 97 nsew signal output
rlabel metal2 s 16578 123200 16634 124000 6 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 121056 688 121856 808 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 io_oeb[4]
port 100 nsew signal output
rlabel metal2 s 104898 0 104954 800 6 io_oeb[5]
port 101 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 io_oeb[6]
port 102 nsew signal output
rlabel metal2 s 25778 123200 25834 124000 6 io_oeb[7]
port 103 nsew signal output
rlabel metal2 s 76378 0 76434 800 6 io_oeb[8]
port 104 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 io_oeb[9]
port 105 nsew signal output
rlabel metal2 s 55678 123200 55734 124000 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 io_out[10]
port 107 nsew signal output
rlabel metal2 s 60738 0 60794 800 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 121056 75488 121856 75608 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 0 73448 800 73568 6 io_out[13]
port 110 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 106738 123200 106794 124000 6 io_out[15]
port 112 nsew signal output
rlabel metal3 s 121056 118328 121856 118448 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 6918 123200 6974 124000 6 io_out[17]
port 114 nsew signal output
rlabel metal3 s 121056 18368 121856 18488 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 0 106768 800 106888 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 81898 123200 81954 124000 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 53378 123200 53434 124000 6 io_out[21]
port 119 nsew signal output
rlabel metal3 s 0 89768 800 89888 6 io_out[22]
port 120 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s 121056 106088 121856 106208 6 io_out[24]
port 122 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 io_out[25]
port 123 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 io_out[26]
port 124 nsew signal output
rlabel metal2 s 110418 123200 110474 124000 6 io_out[27]
port 125 nsew signal output
rlabel metal2 s 103978 0 104034 800 6 io_out[28]
port 126 nsew signal output
rlabel metal2 s 73158 0 73214 800 6 io_out[29]
port 127 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 io_out[2]
port 128 nsew signal output
rlabel metal2 s 42798 123200 42854 124000 6 io_out[30]
port 129 nsew signal output
rlabel metal3 s 121056 73448 121856 73568 6 io_out[31]
port 130 nsew signal output
rlabel metal3 s 0 97248 800 97368 6 io_out[32]
port 131 nsew signal output
rlabel metal2 s 46938 123200 46994 124000 6 io_out[33]
port 132 nsew signal output
rlabel metal2 s 2318 123200 2374 124000 6 io_out[34]
port 133 nsew signal output
rlabel metal3 s 121056 55768 121856 55888 6 io_out[35]
port 134 nsew signal output
rlabel metal2 s 7838 123200 7894 124000 6 io_out[36]
port 135 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 io_out[37]
port 136 nsew signal output
rlabel metal2 s 117778 123200 117834 124000 6 io_out[3]
port 137 nsew signal output
rlabel metal2 s 95238 123200 95294 124000 6 io_out[4]
port 138 nsew signal output
rlabel metal2 s 115018 123200 115074 124000 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 0 70728 800 70848 6 io_out[6]
port 140 nsew signal output
rlabel metal2 s 107658 123200 107714 124000 6 io_out[7]
port 141 nsew signal output
rlabel metal2 s 110418 0 110474 800 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 0 68688 800 68808 6 io_out[9]
port 143 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 la_data_in[100]
port 145 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 la_data_in[101]
port 146 nsew signal input
rlabel metal3 s 121056 31968 121856 32088 6 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 89258 123200 89314 124000 6 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_data_in[104]
port 149 nsew signal input
rlabel metal3 s 0 86368 800 86488 6 la_data_in[105]
port 150 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 la_data_in[106]
port 151 nsew signal input
rlabel metal3 s 121056 94528 121856 94648 6 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 la_data_in[109]
port 154 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 la_data_in[10]
port 155 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 la_data_in[110]
port 156 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 la_data_in[111]
port 157 nsew signal input
rlabel metal3 s 0 97928 800 98048 6 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 65338 123200 65394 124000 6 la_data_in[114]
port 160 nsew signal input
rlabel metal3 s 121056 29248 121856 29368 6 la_data_in[115]
port 161 nsew signal input
rlabel metal3 s 121056 77528 121856 77648 6 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 938 0 994 800 6 la_data_in[118]
port 164 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 la_data_in[119]
port 165 nsew signal input
rlabel metal3 s 121056 48968 121856 49088 6 la_data_in[11]
port 166 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 96618 123200 96674 124000 6 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 36818 123200 36874 124000 6 la_data_in[124]
port 171 nsew signal input
rlabel metal3 s 121056 13608 121856 13728 6 la_data_in[125]
port 172 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 13358 123200 13414 124000 6 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 52918 123200 52974 124000 6 la_data_in[12]
port 175 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 la_data_in[13]
port 176 nsew signal input
rlabel metal3 s 121056 119008 121856 119128 6 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 la_data_in[15]
port 178 nsew signal input
rlabel metal3 s 0 99968 800 100088 6 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 478 123200 534 124000 6 la_data_in[17]
port 180 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 8758 123200 8814 124000 6 la_data_in[19]
port 182 nsew signal input
rlabel metal3 s 121056 51688 121856 51808 6 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 88338 123200 88394 124000 6 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 74078 123200 74134 124000 6 la_data_in[21]
port 185 nsew signal input
rlabel metal3 s 121056 54408 121856 54528 6 la_data_in[22]
port 186 nsew signal input
rlabel metal3 s 121056 112208 121856 112328 6 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 80978 123200 81034 124000 6 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_data_in[27]
port 191 nsew signal input
rlabel metal3 s 121056 23128 121856 23248 6 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 64418 123200 64474 124000 6 la_data_in[2]
port 194 nsew signal input
rlabel metal3 s 121056 41488 121856 41608 6 la_data_in[30]
port 195 nsew signal input
rlabel metal3 s 121056 12248 121856 12368 6 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 23478 123200 23534 124000 6 la_data_in[32]
port 197 nsew signal input
rlabel metal3 s 121056 113568 121856 113688 6 la_data_in[33]
port 198 nsew signal input
rlabel metal3 s 121056 44888 121856 45008 6 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 97998 123200 98054 124000 6 la_data_in[35]
port 200 nsew signal input
rlabel metal3 s 121056 25168 121856 25288 6 la_data_in[36]
port 201 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 la_data_in[37]
port 202 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 116858 123200 116914 124000 6 la_data_in[39]
port 204 nsew signal input
rlabel metal3 s 121056 31288 121856 31408 6 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 103058 123200 103114 124000 6 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 la_data_in[41]
port 207 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 38198 123200 38254 124000 6 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 86498 123200 86554 124000 6 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 60738 123200 60794 124000 6 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 28538 123200 28594 124000 6 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 20258 123200 20314 124000 6 la_data_in[47]
port 213 nsew signal input
rlabel metal3 s 121056 104728 121856 104848 6 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 4158 123200 4214 124000 6 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_data_in[4]
port 216 nsew signal input
rlabel metal3 s 121056 76168 121856 76288 6 la_data_in[50]
port 217 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 56138 123200 56194 124000 6 la_data_in[52]
port 219 nsew signal input
rlabel metal3 s 121056 89088 121856 89208 6 la_data_in[53]
port 220 nsew signal input
rlabel metal3 s 121056 106768 121856 106888 6 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 40958 123200 41014 124000 6 la_data_in[55]
port 222 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 43258 123200 43314 124000 6 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 112718 123200 112774 124000 6 la_data_in[59]
port 226 nsew signal input
rlabel metal3 s 121056 44208 121856 44328 6 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 108118 123200 108174 124000 6 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 59818 123200 59874 124000 6 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 105358 123200 105414 124000 6 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 51538 123200 51594 124000 6 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 62118 123200 62174 124000 6 la_data_in[65]
port 233 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[67]
port 235 nsew signal input
rlabel metal3 s 121056 36048 121856 36168 6 la_data_in[68]
port 236 nsew signal input
rlabel metal3 s 121056 121048 121856 121168 6 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 la_data_in[6]
port 238 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 la_data_in[70]
port 239 nsew signal input
rlabel metal3 s 121056 99288 121856 99408 6 la_data_in[71]
port 240 nsew signal input
rlabel metal3 s 121056 108808 121856 108928 6 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 80518 123200 80574 124000 6 la_data_in[73]
port 242 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 la_data_in[74]
port 243 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 26698 123200 26754 124000 6 la_data_in[78]
port 247 nsew signal input
rlabel metal3 s 121056 63248 121856 63368 6 la_data_in[79]
port 248 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 13818 123200 13874 124000 6 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 104438 123200 104494 124000 6 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 120078 123200 120134 124000 6 la_data_in[84]
port 254 nsew signal input
rlabel metal3 s 0 108128 800 108248 6 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 67638 123200 67694 124000 6 la_data_in[86]
port 256 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 19798 123200 19854 124000 6 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 65798 123200 65854 124000 6 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_data_in[8]
port 260 nsew signal input
rlabel metal3 s 121056 79568 121856 79688 6 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 91558 123200 91614 124000 6 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 44178 123200 44234 124000 6 la_data_in[93]
port 264 nsew signal input
rlabel metal3 s 0 114248 800 114368 6 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 87418 123200 87474 124000 6 la_data_in[98]
port 269 nsew signal input
rlabel metal3 s 121056 68008 121856 68128 6 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 102138 123200 102194 124000 6 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 la_data_out[100]
port 273 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 la_data_out[101]
port 274 nsew signal output
rlabel metal3 s 121056 84328 121856 84448 6 la_data_out[102]
port 275 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 69018 123200 69074 124000 6 la_data_out[104]
port 277 nsew signal output
rlabel metal3 s 0 112208 800 112328 6 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 85118 0 85174 800 6 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 la_data_out[107]
port 280 nsew signal output
rlabel metal3 s 121056 1368 121856 1488 6 la_data_out[108]
port 281 nsew signal output
rlabel metal3 s 0 102008 800 102128 6 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 36358 123200 36414 124000 6 la_data_out[10]
port 283 nsew signal output
rlabel metal3 s 0 64608 800 64728 6 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 23018 123200 23074 124000 6 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 97078 123200 97134 124000 6 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 76838 123200 76894 124000 6 la_data_out[114]
port 288 nsew signal output
rlabel metal3 s 0 65968 800 66088 6 la_data_out[115]
port 289 nsew signal output
rlabel metal3 s 0 67328 800 67448 6 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 32218 123200 32274 124000 6 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 28998 123200 29054 124000 6 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 120998 123200 121054 124000 6 la_data_out[119]
port 293 nsew signal output
rlabel metal3 s 121056 92488 121856 92608 6 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 la_data_out[120]
port 295 nsew signal output
rlabel metal3 s 0 116968 800 117088 6 la_data_out[121]
port 296 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 119158 123200 119214 124000 6 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 116858 0 116914 800 6 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 la_data_out[125]
port 300 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 la_data_out[126]
port 301 nsew signal output
rlabel metal3 s 0 112888 800 113008 6 la_data_out[127]
port 302 nsew signal output
rlabel metal3 s 121056 70048 121856 70168 6 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 108118 0 108174 800 6 la_data_out[13]
port 304 nsew signal output
rlabel metal3 s 121056 53728 121856 53848 6 la_data_out[14]
port 305 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 118238 0 118294 800 6 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 41418 123200 41474 124000 6 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 84198 0 84254 800 6 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 90178 123200 90234 124000 6 la_data_out[21]
port 313 nsew signal output
rlabel metal3 s 121056 89768 121856 89888 6 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 48318 123200 48374 124000 6 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 44638 123200 44694 124000 6 la_data_out[24]
port 316 nsew signal output
rlabel metal3 s 121056 110848 121856 110968 6 la_data_out[25]
port 317 nsew signal output
rlabel metal3 s 121056 8168 121856 8288 6 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 la_data_out[27]
port 319 nsew signal output
rlabel metal3 s 121056 34008 121856 34128 6 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 la_data_out[2]
port 322 nsew signal output
rlabel metal3 s 121056 56448 121856 56568 6 la_data_out[30]
port 323 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 la_data_out[31]
port 324 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 23938 123200 23994 124000 6 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 la_data_out[34]
port 327 nsew signal output
rlabel metal3 s 121056 59168 121856 59288 6 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 117778 0 117834 800 6 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 102138 0 102194 800 6 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 116398 123200 116454 124000 6 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 la_data_out[39]
port 332 nsew signal output
rlabel metal3 s 0 103368 800 103488 6 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 la_data_out[41]
port 335 nsew signal output
rlabel metal3 s 121056 65968 121856 66088 6 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 98458 0 98514 800 6 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 111798 0 111854 800 6 la_data_out[45]
port 339 nsew signal output
rlabel metal3 s 121056 27208 121856 27328 6 la_data_out[46]
port 340 nsew signal output
rlabel metal3 s 121056 17008 121856 17128 6 la_data_out[47]
port 341 nsew signal output
rlabel metal3 s 121056 6128 121856 6248 6 la_data_out[48]
port 342 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 la_data_out[49]
port 343 nsew signal output
rlabel metal3 s 121056 72088 121856 72208 6 la_data_out[4]
port 344 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 85578 123200 85634 124000 6 la_data_out[51]
port 346 nsew signal output
rlabel metal3 s 121056 62568 121856 62688 6 la_data_out[52]
port 347 nsew signal output
rlabel metal3 s 121056 120368 121856 120488 6 la_data_out[53]
port 348 nsew signal output
rlabel metal3 s 121056 123088 121856 123208 6 la_data_out[54]
port 349 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 103058 0 103114 800 6 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 52458 123200 52514 124000 6 la_data_out[58]
port 353 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 104898 123200 104954 124000 6 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 105358 0 105414 800 6 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 la_data_out[61]
port 357 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 la_data_out[62]
port 358 nsew signal output
rlabel metal3 s 121056 34688 121856 34808 6 la_data_out[63]
port 359 nsew signal output
rlabel metal3 s 121056 43528 121856 43648 6 la_data_out[64]
port 360 nsew signal output
rlabel metal3 s 121056 19728 121856 19848 6 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 67178 123200 67234 124000 6 la_data_out[66]
port 362 nsew signal output
rlabel metal3 s 121056 24488 121856 24608 6 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 66258 123200 66314 124000 6 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 la_data_out[69]
port 365 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 34978 123200 35034 124000 6 la_data_out[70]
port 367 nsew signal output
rlabel metal3 s 121056 111528 121856 111648 6 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 115938 123200 115994 124000 6 la_data_out[72]
port 369 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 la_data_out[73]
port 370 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 61658 0 61714 800 6 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 40038 0 40094 800 6 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 la_data_out[77]
port 374 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 70398 123200 70454 124000 6 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 118238 123200 118294 124000 6 la_data_out[7]
port 377 nsew signal output
rlabel metal3 s 121056 82288 121856 82408 6 la_data_out[80]
port 378 nsew signal output
rlabel metal3 s 121056 22448 121856 22568 6 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 57978 123200 58034 124000 6 la_data_out[82]
port 380 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 100298 0 100354 800 6 la_data_out[85]
port 383 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 la_data_out[86]
port 384 nsew signal output
rlabel metal3 s 121056 48288 121856 48408 6 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 109958 123200 110014 124000 6 la_data_out[88]
port 386 nsew signal output
rlabel metal3 s 0 83648 800 83768 6 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 84198 123200 84254 124000 6 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 18878 123200 18934 124000 6 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 17038 123200 17094 124000 6 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 83738 123200 83794 124000 6 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 93858 123200 93914 124000 6 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 1398 0 1454 800 6 la_data_out[94]
port 393 nsew signal output
rlabel metal3 s 121056 42168 121856 42288 6 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 38658 123200 38714 124000 6 la_data_out[96]
port 395 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 la_data_out[98]
port 397 nsew signal output
rlabel metal3 s 121056 90448 121856 90568 6 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 64878 0 64934 800 6 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 la_oenb[100]
port 401 nsew signal input
rlabel metal3 s 121056 5448 121856 5568 6 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 29918 123200 29974 124000 6 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 la_oenb[104]
port 405 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 la_oenb[105]
port 406 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 la_oenb[106]
port 407 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 71318 123200 71374 124000 6 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 34518 123200 34574 124000 6 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 46478 123200 46534 124000 6 la_oenb[110]
port 412 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 la_oenb[111]
port 413 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_oenb[113]
port 415 nsew signal input
rlabel metal3 s 121056 116288 121856 116408 6 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 la_oenb[115]
port 417 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 37738 123200 37794 124000 6 la_oenb[117]
port 419 nsew signal input
rlabel metal3 s 121056 101328 121856 101448 6 la_oenb[118]
port 420 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 109498 123200 109554 124000 6 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_oenb[120]
port 423 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 la_oenb[121]
port 424 nsew signal input
rlabel metal3 s 121056 85688 121856 85808 6 la_oenb[122]
port 425 nsew signal input
rlabel metal3 s 121056 12928 121856 13048 6 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 4618 123200 4674 124000 6 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 la_oenb[127]
port 430 nsew signal input
rlabel metal3 s 121056 99968 121856 100088 6 la_oenb[12]
port 431 nsew signal input
rlabel metal3 s 121056 82968 121856 83088 6 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 98918 123200 98974 124000 6 la_oenb[14]
port 433 nsew signal input
rlabel metal3 s 121056 85008 121856 85128 6 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 14278 123200 14334 124000 6 la_oenb[17]
port 436 nsew signal input
rlabel metal3 s 121056 78208 121856 78328 6 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 la_oenb[19]
port 438 nsew signal input
rlabel metal3 s 0 121728 800 121848 6 la_oenb[1]
port 439 nsew signal input
rlabel metal3 s 121056 65288 121856 65408 6 la_oenb[20]
port 440 nsew signal input
rlabel metal3 s 0 105408 800 105528 6 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 63038 123200 63094 124000 6 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 45098 123200 45154 124000 6 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 94778 123200 94834 124000 6 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 10598 123200 10654 124000 6 la_oenb[27]
port 447 nsew signal input
rlabel metal3 s 121056 10208 121856 10328 6 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_oenb[29]
port 449 nsew signal input
rlabel metal3 s 121056 67328 121856 67448 6 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 la_oenb[31]
port 452 nsew signal input
rlabel metal3 s 121056 49648 121856 49768 6 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 62578 123200 62634 124000 6 la_oenb[33]
port 454 nsew signal input
rlabel metal3 s 121056 39448 121856 39568 6 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 120998 0 121054 800 6 la_oenb[37]
port 458 nsew signal input
rlabel metal3 s 121056 107448 121856 107568 6 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 la_oenb[39]
port 460 nsew signal input
rlabel metal3 s 0 95888 800 96008 6 la_oenb[3]
port 461 nsew signal input
rlabel metal3 s 0 85008 800 85128 6 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 75458 123200 75514 124000 6 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_oenb[42]
port 464 nsew signal input
rlabel metal3 s 121056 53048 121856 53168 6 la_oenb[43]
port 465 nsew signal input
rlabel metal3 s 0 109488 800 109608 6 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 la_oenb[45]
port 467 nsew signal input
rlabel metal3 s 121056 46928 121856 47048 6 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 114558 123200 114614 124000 6 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 49238 123200 49294 124000 6 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 478 0 534 800 6 la_oenb[4]
port 472 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 938 123200 994 124000 6 la_oenb[51]
port 474 nsew signal input
rlabel metal3 s 121056 26528 121856 26648 6 la_oenb[52]
port 475 nsew signal input
rlabel metal3 s 121056 60528 121856 60648 6 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_oenb[54]
port 477 nsew signal input
rlabel metal3 s 0 92488 800 92608 6 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 28078 123200 28134 124000 6 la_oenb[56]
port 479 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 63958 123200 64014 124000 6 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 82358 123200 82414 124000 6 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_oenb[60]
port 484 nsew signal input
rlabel metal3 s 121056 38768 121856 38888 6 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 la_oenb[62]
port 486 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 la_oenb[63]
port 487 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 la_oenb[64]
port 488 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 7378 123200 7434 124000 6 la_oenb[66]
port 490 nsew signal input
rlabel metal3 s 121056 15648 121856 15768 6 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 69478 123200 69534 124000 6 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 86958 123200 87014 124000 6 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 33598 123200 33654 124000 6 la_oenb[71]
port 496 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 54298 123200 54354 124000 6 la_oenb[74]
port 499 nsew signal input
rlabel metal3 s 0 114928 800 115048 6 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 12438 123200 12494 124000 6 la_oenb[76]
port 501 nsew signal input
rlabel metal3 s 121056 4768 121856 4888 6 la_oenb[77]
port 502 nsew signal input
rlabel metal3 s 0 121048 800 121168 6 la_oenb[78]
port 503 nsew signal input
rlabel metal3 s 121056 29928 121856 30048 6 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 la_oenb[7]
port 505 nsew signal input
rlabel metal3 s 121056 103368 121856 103488 6 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 92018 123200 92074 124000 6 la_oenb[81]
port 507 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_oenb[83]
port 509 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 la_oenb[84]
port 510 nsew signal input
rlabel metal3 s 121056 57808 121856 57928 6 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 103518 123200 103574 124000 6 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 51078 123200 51134 124000 6 la_oenb[87]
port 513 nsew signal input
rlabel metal3 s 121056 116968 121856 117088 6 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 la_oenb[89]
port 515 nsew signal input
rlabel metal3 s 121056 93848 121856 93968 6 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 77758 123200 77814 124000 6 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 119618 123200 119674 124000 6 la_oenb[93]
port 520 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 la_oenb[94]
port 521 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 la_oenb[96]
port 523 nsew signal input
rlabel metal3 s 121056 102008 121856 102128 6 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 61198 123200 61254 124000 6 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 101678 123200 101734 124000 6 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 user_clock2
port 528 nsew signal input
rlabel metal2 s 17498 123200 17554 124000 6 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 88798 123200 88854 124000 6 user_irq[2]
port 531 nsew signal output
rlabel metal2 s 58898 123200 58954 124000 6 wb_clk_i
port 532 nsew signal input
rlabel metal3 s 121056 3408 121856 3528 6 wb_rst_i
port 533 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 wbs_ack_o
port 534 nsew signal output
rlabel metal2 s 57518 123200 57574 124000 6 wbs_adr_i[0]
port 535 nsew signal input
rlabel metal3 s 121056 36728 121856 36848 6 wbs_adr_i[10]
port 536 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 wbs_adr_i[11]
port 537 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 wbs_adr_i[12]
port 538 nsew signal input
rlabel metal3 s 0 119688 800 119808 6 wbs_adr_i[13]
port 539 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 wbs_adr_i[14]
port 540 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 wbs_adr_i[15]
port 541 nsew signal input
rlabel metal3 s 121056 96568 121856 96688 6 wbs_adr_i[16]
port 542 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 wbs_adr_i[17]
port 543 nsew signal input
rlabel metal3 s 121056 9528 121856 9648 6 wbs_adr_i[18]
port 544 nsew signal input
rlabel metal2 s 72698 123200 72754 124000 6 wbs_adr_i[19]
port 545 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_adr_i[1]
port 546 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 wbs_adr_i[20]
port 547 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[21]
port 548 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 wbs_adr_i[22]
port 549 nsew signal input
rlabel metal2 s 49698 123200 49754 124000 6 wbs_adr_i[23]
port 550 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_adr_i[24]
port 551 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 wbs_adr_i[25]
port 552 nsew signal input
rlabel metal3 s 0 95208 800 95328 6 wbs_adr_i[26]
port 553 nsew signal input
rlabel metal2 s 78678 123200 78734 124000 6 wbs_adr_i[27]
port 554 nsew signal input
rlabel metal2 s 5998 123200 6054 124000 6 wbs_adr_i[28]
port 555 nsew signal input
rlabel metal3 s 121056 121728 121856 121848 6 wbs_adr_i[29]
port 556 nsew signal input
rlabel metal2 s 15198 123200 15254 124000 6 wbs_adr_i[2]
port 557 nsew signal input
rlabel metal2 s 47858 123200 47914 124000 6 wbs_adr_i[30]
port 558 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_adr_i[31]
port 559 nsew signal input
rlabel metal3 s 121056 68688 121856 68808 6 wbs_adr_i[3]
port 560 nsew signal input
rlabel metal2 s 25318 123200 25374 124000 6 wbs_adr_i[4]
port 561 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 wbs_adr_i[5]
port 562 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 wbs_adr_i[6]
port 563 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 wbs_adr_i[7]
port 564 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 wbs_adr_i[8]
port 565 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 wbs_adr_i[9]
port 566 nsew signal input
rlabel metal2 s 59358 123200 59414 124000 6 wbs_cyc_i
port 567 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 wbs_dat_i[0]
port 568 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 wbs_dat_i[10]
port 569 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 wbs_dat_i[11]
port 570 nsew signal input
rlabel metal2 s 99838 123200 99894 124000 6 wbs_dat_i[12]
port 571 nsew signal input
rlabel metal3 s 121056 104048 121856 104168 6 wbs_dat_i[13]
port 572 nsew signal input
rlabel metal3 s 121056 37408 121856 37528 6 wbs_dat_i[14]
port 573 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 wbs_dat_i[15]
port 574 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 wbs_dat_i[16]
port 575 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 wbs_dat_i[17]
port 576 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 wbs_dat_i[18]
port 577 nsew signal input
rlabel metal2 s 83278 123200 83334 124000 6 wbs_dat_i[19]
port 578 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 wbs_dat_i[1]
port 579 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 wbs_dat_i[20]
port 580 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_i[21]
port 581 nsew signal input
rlabel metal2 s 111798 123200 111854 124000 6 wbs_dat_i[22]
port 582 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 wbs_dat_i[23]
port 583 nsew signal input
rlabel metal2 s 11978 123200 12034 124000 6 wbs_dat_i[24]
port 584 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_i[25]
port 585 nsew signal input
rlabel metal3 s 121056 14968 121856 15088 6 wbs_dat_i[26]
port 586 nsew signal input
rlabel metal3 s 121056 40808 121856 40928 6 wbs_dat_i[27]
port 587 nsew signal input
rlabel metal2 s 39578 123200 39634 124000 6 wbs_dat_i[28]
port 588 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 wbs_dat_i[29]
port 589 nsew signal input
rlabel metal3 s 121056 115608 121856 115728 6 wbs_dat_i[2]
port 590 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_i[30]
port 591 nsew signal input
rlabel metal2 s 30378 123200 30434 124000 6 wbs_dat_i[31]
port 592 nsew signal input
rlabel metal2 s 79138 123200 79194 124000 6 wbs_dat_i[3]
port 593 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 wbs_dat_i[4]
port 594 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_i[5]
port 595 nsew signal input
rlabel metal2 s 95698 123200 95754 124000 6 wbs_dat_i[6]
port 596 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wbs_dat_i[7]
port 597 nsew signal input
rlabel metal2 s 75918 123200 75974 124000 6 wbs_dat_i[8]
port 598 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 wbs_dat_i[9]
port 599 nsew signal input
rlabel metal2 s 3698 123200 3754 124000 6 wbs_dat_o[0]
port 600 nsew signal output
rlabel metal3 s 121056 98608 121856 98728 6 wbs_dat_o[10]
port 601 nsew signal output
rlabel metal2 s 78678 0 78734 800 6 wbs_dat_o[11]
port 602 nsew signal output
rlabel metal2 s 113638 0 113694 800 6 wbs_dat_o[12]
port 603 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_o[13]
port 604 nsew signal output
rlabel metal3 s 0 90448 800 90568 6 wbs_dat_o[14]
port 605 nsew signal output
rlabel metal2 s 115478 0 115534 800 6 wbs_dat_o[15]
port 606 nsew signal output
rlabel metal2 s 93398 123200 93454 124000 6 wbs_dat_o[16]
port 607 nsew signal output
rlabel metal2 s 1858 123200 1914 124000 6 wbs_dat_o[17]
port 608 nsew signal output
rlabel metal3 s 121056 61208 121856 61328 6 wbs_dat_o[18]
port 609 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 wbs_dat_o[19]
port 610 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 wbs_dat_o[1]
port 611 nsew signal output
rlabel metal2 s 50158 123200 50214 124000 6 wbs_dat_o[20]
port 612 nsew signal output
rlabel metal2 s 27158 123200 27214 124000 6 wbs_dat_o[21]
port 613 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 wbs_dat_o[22]
port 614 nsew signal output
rlabel metal2 s 5538 123200 5594 124000 6 wbs_dat_o[23]
port 615 nsew signal output
rlabel metal2 s 77298 123200 77354 124000 6 wbs_dat_o[24]
port 616 nsew signal output
rlabel metal3 s 121056 80928 121856 81048 6 wbs_dat_o[25]
port 617 nsew signal output
rlabel metal2 s 85118 123200 85174 124000 6 wbs_dat_o[26]
port 618 nsew signal output
rlabel metal2 s 100298 123200 100354 124000 6 wbs_dat_o[27]
port 619 nsew signal output
rlabel metal3 s 121056 32648 121856 32768 6 wbs_dat_o[28]
port 620 nsew signal output
rlabel metal2 s 18418 123200 18474 124000 6 wbs_dat_o[29]
port 621 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 wbs_dat_o[2]
port 622 nsew signal output
rlabel metal2 s 92478 123200 92534 124000 6 wbs_dat_o[30]
port 623 nsew signal output
rlabel metal2 s 33138 123200 33194 124000 6 wbs_dat_o[31]
port 624 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 wbs_dat_o[3]
port 625 nsew signal output
rlabel metal2 s 20718 123200 20774 124000 6 wbs_dat_o[4]
port 626 nsew signal output
rlabel metal2 s 72238 123200 72294 124000 6 wbs_dat_o[5]
port 627 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 wbs_dat_o[6]
port 628 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_o[7]
port 629 nsew signal output
rlabel metal3 s 121056 87048 121856 87168 6 wbs_dat_o[8]
port 630 nsew signal output
rlabel metal3 s 121056 87728 121856 87848 6 wbs_dat_o[9]
port 631 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 wbs_sel_i[0]
port 632 nsew signal input
rlabel metal2 s 11058 123200 11114 124000 6 wbs_sel_i[1]
port 633 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 wbs_sel_i[2]
port 634 nsew signal input
rlabel metal2 s 22098 123200 22154 124000 6 wbs_sel_i[3]
port 635 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 wbs_stb_i
port 636 nsew signal input
rlabel metal2 s 68098 123200 68154 124000 6 wbs_we_i
port 637 nsew signal input
rlabel metal4 s 108804 -1864 109404 125352 6 vccd1
port 638 nsew power bidirectional
rlabel metal4 s 72804 -1864 73404 125352 6 vccd1
port 639 nsew power bidirectional
rlabel metal4 s 36804 -1864 37404 125352 6 vccd1
port 640 nsew power bidirectional
rlabel metal4 s 804 -1864 1404 125352 6 vccd1
port 641 nsew power bidirectional
rlabel metal4 s 123204 -924 123804 124412 6 vccd1
port 642 nsew power bidirectional
rlabel metal4 s -1996 -924 -1396 124412 4 vccd1
port 643 nsew power bidirectional
rlabel metal5 s -1996 123812 123804 124412 6 vccd1
port 644 nsew power bidirectional
rlabel metal5 s -2936 109828 124744 110428 6 vccd1
port 645 nsew power bidirectional
rlabel metal5 s -2936 73828 124744 74428 6 vccd1
port 646 nsew power bidirectional
rlabel metal5 s -2936 37828 124744 38428 6 vccd1
port 647 nsew power bidirectional
rlabel metal5 s -2936 1828 124744 2428 6 vccd1
port 648 nsew power bidirectional
rlabel metal5 s -1996 -924 123804 -324 8 vccd1
port 649 nsew power bidirectional
rlabel metal4 s 124144 -1864 124744 125352 6 vssd1
port 650 nsew ground bidirectional
rlabel metal4 s 90804 -1864 91404 125352 6 vssd1
port 651 nsew ground bidirectional
rlabel metal4 s 54804 -1864 55404 125352 6 vssd1
port 652 nsew ground bidirectional
rlabel metal4 s 18804 -1864 19404 125352 6 vssd1
port 653 nsew ground bidirectional
rlabel metal4 s -2936 -1864 -2336 125352 4 vssd1
port 654 nsew ground bidirectional
rlabel metal5 s -2936 124752 124744 125352 6 vssd1
port 655 nsew ground bidirectional
rlabel metal5 s -2936 91828 124744 92428 6 vssd1
port 656 nsew ground bidirectional
rlabel metal5 s -2936 55828 124744 56428 6 vssd1
port 657 nsew ground bidirectional
rlabel metal5 s -2936 19828 124744 20428 6 vssd1
port 658 nsew ground bidirectional
rlabel metal5 s -2936 -1864 124744 -1264 8 vssd1
port 659 nsew ground bidirectional
rlabel metal4 s 112404 -3744 113004 127232 6 vccd2
port 660 nsew power bidirectional
rlabel metal4 s 76404 -3744 77004 127232 6 vccd2
port 661 nsew power bidirectional
rlabel metal4 s 40404 -3744 41004 127232 6 vccd2
port 662 nsew power bidirectional
rlabel metal4 s 4404 -3744 5004 127232 6 vccd2
port 663 nsew power bidirectional
rlabel metal4 s 125084 -2804 125684 126292 6 vccd2
port 664 nsew power bidirectional
rlabel metal4 s -3876 -2804 -3276 126292 4 vccd2
port 665 nsew power bidirectional
rlabel metal5 s -3876 125692 125684 126292 6 vccd2
port 666 nsew power bidirectional
rlabel metal5 s -4816 113476 126624 114076 6 vccd2
port 667 nsew power bidirectional
rlabel metal5 s -4816 77476 126624 78076 6 vccd2
port 668 nsew power bidirectional
rlabel metal5 s -4816 41476 126624 42076 6 vccd2
port 669 nsew power bidirectional
rlabel metal5 s -4816 5476 126624 6076 6 vccd2
port 670 nsew power bidirectional
rlabel metal5 s -3876 -2804 125684 -2204 8 vccd2
port 671 nsew power bidirectional
rlabel metal4 s 126024 -3744 126624 127232 6 vssd2
port 672 nsew ground bidirectional
rlabel metal4 s 94404 -3744 95004 127232 6 vssd2
port 673 nsew ground bidirectional
rlabel metal4 s 58404 -3744 59004 127232 6 vssd2
port 674 nsew ground bidirectional
rlabel metal4 s 22404 -3744 23004 127232 6 vssd2
port 675 nsew ground bidirectional
rlabel metal4 s -4816 -3744 -4216 127232 4 vssd2
port 676 nsew ground bidirectional
rlabel metal5 s -4816 126632 126624 127232 6 vssd2
port 677 nsew ground bidirectional
rlabel metal5 s -4816 95476 126624 96076 6 vssd2
port 678 nsew ground bidirectional
rlabel metal5 s -4816 59476 126624 60076 6 vssd2
port 679 nsew ground bidirectional
rlabel metal5 s -4816 23476 126624 24076 6 vssd2
port 680 nsew ground bidirectional
rlabel metal5 s -4816 -3744 126624 -3144 8 vssd2
port 681 nsew ground bidirectional
rlabel metal4 s 116004 -5624 116604 129112 6 vdda1
port 682 nsew power bidirectional
rlabel metal4 s 80004 -5624 80604 129112 6 vdda1
port 683 nsew power bidirectional
rlabel metal4 s 44004 -5624 44604 129112 6 vdda1
port 684 nsew power bidirectional
rlabel metal4 s 8004 -5624 8604 129112 6 vdda1
port 685 nsew power bidirectional
rlabel metal4 s 126964 -4684 127564 128172 6 vdda1
port 686 nsew power bidirectional
rlabel metal4 s -5756 -4684 -5156 128172 4 vdda1
port 687 nsew power bidirectional
rlabel metal5 s -5756 127572 127564 128172 6 vdda1
port 688 nsew power bidirectional
rlabel metal5 s -6696 117076 128504 117676 6 vdda1
port 689 nsew power bidirectional
rlabel metal5 s -6696 81076 128504 81676 6 vdda1
port 690 nsew power bidirectional
rlabel metal5 s -6696 45076 128504 45676 6 vdda1
port 691 nsew power bidirectional
rlabel metal5 s -6696 9076 128504 9676 6 vdda1
port 692 nsew power bidirectional
rlabel metal5 s -5756 -4684 127564 -4084 8 vdda1
port 693 nsew power bidirectional
rlabel metal4 s 127904 -5624 128504 129112 6 vssa1
port 694 nsew ground bidirectional
rlabel metal4 s 98004 -5624 98604 129112 6 vssa1
port 695 nsew ground bidirectional
rlabel metal4 s 62004 -5624 62604 129112 6 vssa1
port 696 nsew ground bidirectional
rlabel metal4 s 26004 -5624 26604 129112 6 vssa1
port 697 nsew ground bidirectional
rlabel metal4 s -6696 -5624 -6096 129112 4 vssa1
port 698 nsew ground bidirectional
rlabel metal5 s -6696 128512 128504 129112 6 vssa1
port 699 nsew ground bidirectional
rlabel metal5 s -6696 99076 128504 99676 6 vssa1
port 700 nsew ground bidirectional
rlabel metal5 s -6696 63076 128504 63676 6 vssa1
port 701 nsew ground bidirectional
rlabel metal5 s -6696 27076 128504 27676 6 vssa1
port 702 nsew ground bidirectional
rlabel metal5 s -6696 -5624 128504 -5024 8 vssa1
port 703 nsew ground bidirectional
rlabel metal4 s 119604 -7504 120204 130992 6 vdda2
port 704 nsew power bidirectional
rlabel metal4 s 83604 -7504 84204 130992 6 vdda2
port 705 nsew power bidirectional
rlabel metal4 s 47604 -7504 48204 130992 6 vdda2
port 706 nsew power bidirectional
rlabel metal4 s 11604 -7504 12204 130992 6 vdda2
port 707 nsew power bidirectional
rlabel metal4 s 128844 -6564 129444 130052 6 vdda2
port 708 nsew power bidirectional
rlabel metal4 s -7636 -6564 -7036 130052 4 vdda2
port 709 nsew power bidirectional
rlabel metal5 s -7636 129452 129444 130052 6 vdda2
port 710 nsew power bidirectional
rlabel metal5 s -8576 84676 130384 85276 6 vdda2
port 711 nsew power bidirectional
rlabel metal5 s -8576 48676 130384 49276 6 vdda2
port 712 nsew power bidirectional
rlabel metal5 s -8576 12676 130384 13276 6 vdda2
port 713 nsew power bidirectional
rlabel metal5 s -7636 -6564 129444 -5964 8 vdda2
port 714 nsew power bidirectional
rlabel metal4 s 129784 -7504 130384 130992 6 vssa2
port 715 nsew ground bidirectional
rlabel metal4 s 101604 -7504 102204 130992 6 vssa2
port 716 nsew ground bidirectional
rlabel metal4 s 65604 -7504 66204 130992 6 vssa2
port 717 nsew ground bidirectional
rlabel metal4 s 29604 -7504 30204 130992 6 vssa2
port 718 nsew ground bidirectional
rlabel metal4 s -8576 -7504 -7976 130992 4 vssa2
port 719 nsew ground bidirectional
rlabel metal5 s -8576 130392 130384 130992 6 vssa2
port 720 nsew ground bidirectional
rlabel metal5 s -8576 102676 130384 103276 6 vssa2
port 721 nsew ground bidirectional
rlabel metal5 s -8576 66676 130384 67276 6 vssa2
port 722 nsew ground bidirectional
rlabel metal5 s -8576 30676 130384 31276 6 vssa2
port 723 nsew ground bidirectional
rlabel metal5 s -8576 -7504 130384 -6904 8 vssa2
port 724 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 121856 124000
string LEFview TRUE
string GDS_FILE /project/openlane/user_project_wrapper/runs/user_project_wrapper/results/magic/user_project_wrapper.gds
string GDS_END 32522604
string GDS_START 130
<< end >>

