magic
tech sky130A
magscale 1 2
timestamp 1622197323
<< obsli1 >>
rect 949 1377 142847 143531
<< obsm1 >>
rect 937 1368 143598 143664
<< metal2 >>
rect 938 145428 994 146228
rect 1398 145428 1454 146228
rect 2318 145428 2374 146228
rect 3238 145428 3294 146228
rect 3698 145428 3754 146228
rect 4618 145428 4674 146228
rect 5538 145428 5594 146228
rect 5998 145428 6054 146228
rect 6918 145428 6974 146228
rect 7838 145428 7894 146228
rect 8298 145428 8354 146228
rect 9218 145428 9274 146228
rect 10138 145428 10194 146228
rect 10598 145428 10654 146228
rect 11518 145428 11574 146228
rect 12438 145428 12494 146228
rect 12898 145428 12954 146228
rect 13818 145428 13874 146228
rect 14278 145428 14334 146228
rect 15198 145428 15254 146228
rect 16118 145428 16174 146228
rect 16578 145428 16634 146228
rect 17498 145428 17554 146228
rect 18418 145428 18474 146228
rect 18878 145428 18934 146228
rect 19798 145428 19854 146228
rect 20718 145428 20774 146228
rect 21178 145428 21234 146228
rect 22098 145428 22154 146228
rect 23018 145428 23074 146228
rect 23478 145428 23534 146228
rect 24398 145428 24454 146228
rect 25318 145428 25374 146228
rect 25778 145428 25834 146228
rect 26698 145428 26754 146228
rect 27158 145428 27214 146228
rect 28078 145428 28134 146228
rect 28998 145428 29054 146228
rect 29458 145428 29514 146228
rect 30378 145428 30434 146228
rect 31298 145428 31354 146228
rect 31758 145428 31814 146228
rect 32678 145428 32734 146228
rect 33598 145428 33654 146228
rect 34058 145428 34114 146228
rect 34978 145428 35034 146228
rect 35898 145428 35954 146228
rect 36358 145428 36414 146228
rect 37278 145428 37334 146228
rect 38198 145428 38254 146228
rect 38658 145428 38714 146228
rect 39578 145428 39634 146228
rect 40038 145428 40094 146228
rect 40958 145428 41014 146228
rect 41878 145428 41934 146228
rect 42338 145428 42394 146228
rect 43258 145428 43314 146228
rect 44178 145428 44234 146228
rect 44638 145428 44694 146228
rect 45558 145428 45614 146228
rect 46478 145428 46534 146228
rect 46938 145428 46994 146228
rect 47858 145428 47914 146228
rect 48778 145428 48834 146228
rect 49238 145428 49294 146228
rect 50158 145428 50214 146228
rect 51078 145428 51134 146228
rect 51538 145428 51594 146228
rect 52458 145428 52514 146228
rect 53378 145428 53434 146228
rect 53838 145428 53894 146228
rect 54758 145428 54814 146228
rect 55218 145428 55274 146228
rect 56138 145428 56194 146228
rect 57058 145428 57114 146228
rect 57518 145428 57574 146228
rect 58438 145428 58494 146228
rect 59358 145428 59414 146228
rect 59818 145428 59874 146228
rect 60738 145428 60794 146228
rect 61658 145428 61714 146228
rect 62118 145428 62174 146228
rect 63038 145428 63094 146228
rect 63958 145428 64014 146228
rect 64418 145428 64474 146228
rect 65338 145428 65394 146228
rect 66258 145428 66314 146228
rect 66718 145428 66774 146228
rect 67638 145428 67694 146228
rect 68098 145428 68154 146228
rect 69018 145428 69074 146228
rect 69938 145428 69994 146228
rect 70398 145428 70454 146228
rect 71318 145428 71374 146228
rect 72238 145428 72294 146228
rect 72698 145428 72754 146228
rect 73618 145428 73674 146228
rect 74538 145428 74594 146228
rect 74998 145428 75054 146228
rect 75918 145428 75974 146228
rect 76838 145428 76894 146228
rect 77298 145428 77354 146228
rect 78218 145428 78274 146228
rect 79138 145428 79194 146228
rect 79598 145428 79654 146228
rect 80518 145428 80574 146228
rect 81438 145428 81494 146228
rect 81898 145428 81954 146228
rect 82818 145428 82874 146228
rect 83278 145428 83334 146228
rect 84198 145428 84254 146228
rect 85118 145428 85174 146228
rect 85578 145428 85634 146228
rect 86498 145428 86554 146228
rect 87418 145428 87474 146228
rect 87878 145428 87934 146228
rect 88798 145428 88854 146228
rect 89718 145428 89774 146228
rect 90178 145428 90234 146228
rect 91098 145428 91154 146228
rect 92018 145428 92074 146228
rect 92478 145428 92534 146228
rect 93398 145428 93454 146228
rect 94318 145428 94374 146228
rect 94778 145428 94834 146228
rect 95698 145428 95754 146228
rect 96158 145428 96214 146228
rect 97078 145428 97134 146228
rect 97998 145428 98054 146228
rect 98458 145428 98514 146228
rect 99378 145428 99434 146228
rect 100298 145428 100354 146228
rect 100758 145428 100814 146228
rect 101678 145428 101734 146228
rect 102598 145428 102654 146228
rect 103058 145428 103114 146228
rect 103978 145428 104034 146228
rect 104898 145428 104954 146228
rect 105358 145428 105414 146228
rect 106278 145428 106334 146228
rect 107198 145428 107254 146228
rect 107658 145428 107714 146228
rect 108578 145428 108634 146228
rect 109038 145428 109094 146228
rect 109958 145428 110014 146228
rect 110878 145428 110934 146228
rect 111338 145428 111394 146228
rect 112258 145428 112314 146228
rect 113178 145428 113234 146228
rect 113638 145428 113694 146228
rect 114558 145428 114614 146228
rect 115478 145428 115534 146228
rect 115938 145428 115994 146228
rect 116858 145428 116914 146228
rect 117778 145428 117834 146228
rect 118238 145428 118294 146228
rect 119158 145428 119214 146228
rect 120078 145428 120134 146228
rect 120538 145428 120594 146228
rect 121458 145428 121514 146228
rect 122378 145428 122434 146228
rect 122838 145428 122894 146228
rect 123758 145428 123814 146228
rect 124218 145428 124274 146228
rect 125138 145428 125194 146228
rect 126058 145428 126114 146228
rect 126518 145428 126574 146228
rect 127438 145428 127494 146228
rect 128358 145428 128414 146228
rect 128818 145428 128874 146228
rect 129738 145428 129794 146228
rect 130658 145428 130714 146228
rect 131118 145428 131174 146228
rect 132038 145428 132094 146228
rect 132958 145428 133014 146228
rect 133418 145428 133474 146228
rect 134338 145428 134394 146228
rect 135258 145428 135314 146228
rect 135718 145428 135774 146228
rect 136638 145428 136694 146228
rect 137098 145428 137154 146228
rect 138018 145428 138074 146228
rect 138938 145428 138994 146228
rect 139398 145428 139454 146228
rect 140318 145428 140374 146228
rect 141238 145428 141294 146228
rect 141698 145428 141754 146228
rect 142618 145428 142674 146228
rect 143538 145428 143594 146228
rect 478 0 534 800
rect 938 0 994 800
rect 1858 0 1914 800
rect 2318 0 2374 800
rect 3238 0 3294 800
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 5538 0 5594 800
rect 6458 0 6514 800
rect 6918 0 6974 800
rect 7838 0 7894 800
rect 8758 0 8814 800
rect 9218 0 9274 800
rect 10138 0 10194 800
rect 11058 0 11114 800
rect 11518 0 11574 800
rect 12438 0 12494 800
rect 13358 0 13414 800
rect 13818 0 13874 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 16118 0 16174 800
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 18418 0 18474 800
rect 19338 0 19394 800
rect 19798 0 19854 800
rect 20718 0 20774 800
rect 21638 0 21694 800
rect 22098 0 22154 800
rect 23018 0 23074 800
rect 23938 0 23994 800
rect 24398 0 24454 800
rect 25318 0 25374 800
rect 26238 0 26294 800
rect 26698 0 26754 800
rect 27618 0 27674 800
rect 28078 0 28134 800
rect 28998 0 29054 800
rect 29918 0 29974 800
rect 30378 0 30434 800
rect 31298 0 31354 800
rect 32218 0 32274 800
rect 32678 0 32734 800
rect 33598 0 33654 800
rect 34518 0 34574 800
rect 34978 0 35034 800
rect 35898 0 35954 800
rect 36818 0 36874 800
rect 37278 0 37334 800
rect 38198 0 38254 800
rect 39118 0 39174 800
rect 39578 0 39634 800
rect 40498 0 40554 800
rect 41418 0 41474 800
rect 41878 0 41934 800
rect 42798 0 42854 800
rect 43258 0 43314 800
rect 44178 0 44234 800
rect 45098 0 45154 800
rect 45558 0 45614 800
rect 46478 0 46534 800
rect 47398 0 47454 800
rect 47858 0 47914 800
rect 48778 0 48834 800
rect 49698 0 49754 800
rect 50158 0 50214 800
rect 51078 0 51134 800
rect 51998 0 52054 800
rect 52458 0 52514 800
rect 53378 0 53434 800
rect 54298 0 54354 800
rect 54758 0 54814 800
rect 55678 0 55734 800
rect 56138 0 56194 800
rect 57058 0 57114 800
rect 57978 0 58034 800
rect 58438 0 58494 800
rect 59358 0 59414 800
rect 60278 0 60334 800
rect 60738 0 60794 800
rect 61658 0 61714 800
rect 62578 0 62634 800
rect 63038 0 63094 800
rect 63958 0 64014 800
rect 64878 0 64934 800
rect 65338 0 65394 800
rect 66258 0 66314 800
rect 67178 0 67234 800
rect 67638 0 67694 800
rect 68558 0 68614 800
rect 69478 0 69534 800
rect 69938 0 69994 800
rect 70858 0 70914 800
rect 71318 0 71374 800
rect 72238 0 72294 800
rect 73158 0 73214 800
rect 73618 0 73674 800
rect 74538 0 74594 800
rect 75458 0 75514 800
rect 75918 0 75974 800
rect 76838 0 76894 800
rect 77758 0 77814 800
rect 78218 0 78274 800
rect 79138 0 79194 800
rect 80058 0 80114 800
rect 80518 0 80574 800
rect 81438 0 81494 800
rect 82358 0 82414 800
rect 82818 0 82874 800
rect 83738 0 83794 800
rect 84198 0 84254 800
rect 85118 0 85174 800
rect 86038 0 86094 800
rect 86498 0 86554 800
rect 87418 0 87474 800
rect 88338 0 88394 800
rect 88798 0 88854 800
rect 89718 0 89774 800
rect 90638 0 90694 800
rect 91098 0 91154 800
rect 92018 0 92074 800
rect 92938 0 92994 800
rect 93398 0 93454 800
rect 94318 0 94374 800
rect 95238 0 95294 800
rect 95698 0 95754 800
rect 96618 0 96674 800
rect 97078 0 97134 800
rect 97998 0 98054 800
rect 98918 0 98974 800
rect 99378 0 99434 800
rect 100298 0 100354 800
rect 101218 0 101274 800
rect 101678 0 101734 800
rect 102598 0 102654 800
rect 103518 0 103574 800
rect 103978 0 104034 800
rect 104898 0 104954 800
rect 105818 0 105874 800
rect 106278 0 106334 800
rect 107198 0 107254 800
rect 108118 0 108174 800
rect 108578 0 108634 800
rect 109498 0 109554 800
rect 110418 0 110474 800
rect 110878 0 110934 800
rect 111798 0 111854 800
rect 112258 0 112314 800
rect 113178 0 113234 800
rect 114098 0 114154 800
rect 114558 0 114614 800
rect 115478 0 115534 800
rect 116398 0 116454 800
rect 116858 0 116914 800
rect 117778 0 117834 800
rect 118698 0 118754 800
rect 119158 0 119214 800
rect 120078 0 120134 800
rect 120998 0 121054 800
rect 121458 0 121514 800
rect 122378 0 122434 800
rect 123298 0 123354 800
rect 123758 0 123814 800
rect 124678 0 124734 800
rect 125138 0 125194 800
rect 126058 0 126114 800
rect 126978 0 127034 800
rect 127438 0 127494 800
rect 128358 0 128414 800
rect 129278 0 129334 800
rect 129738 0 129794 800
rect 130658 0 130714 800
rect 131578 0 131634 800
rect 132038 0 132094 800
rect 132958 0 133014 800
rect 133878 0 133934 800
rect 134338 0 134394 800
rect 135258 0 135314 800
rect 136178 0 136234 800
rect 136638 0 136694 800
rect 137558 0 137614 800
rect 138478 0 138534 800
rect 138938 0 138994 800
rect 139858 0 139914 800
rect 140318 0 140374 800
rect 141238 0 141294 800
rect 142158 0 142214 800
rect 142618 0 142674 800
rect 143538 0 143594 800
<< obsm2 >>
rect 1124 145372 1342 145428
rect 1510 145372 2262 145428
rect 2430 145372 3182 145428
rect 3350 145372 3642 145428
rect 3810 145372 4562 145428
rect 4730 145372 5482 145428
rect 5650 145372 5942 145428
rect 6110 145372 6862 145428
rect 7030 145372 7782 145428
rect 7950 145372 8242 145428
rect 8410 145372 9162 145428
rect 9330 145372 10082 145428
rect 10250 145372 10542 145428
rect 10710 145372 11462 145428
rect 11630 145372 12382 145428
rect 12550 145372 12842 145428
rect 13010 145372 13762 145428
rect 13930 145372 14222 145428
rect 14390 145372 15142 145428
rect 15310 145372 16062 145428
rect 16230 145372 16522 145428
rect 16690 145372 17442 145428
rect 17610 145372 18362 145428
rect 18530 145372 18822 145428
rect 18990 145372 19742 145428
rect 19910 145372 20662 145428
rect 20830 145372 21122 145428
rect 21290 145372 22042 145428
rect 22210 145372 22962 145428
rect 23130 145372 23422 145428
rect 23590 145372 24342 145428
rect 24510 145372 25262 145428
rect 25430 145372 25722 145428
rect 25890 145372 26642 145428
rect 26810 145372 27102 145428
rect 27270 145372 28022 145428
rect 28190 145372 28942 145428
rect 29110 145372 29402 145428
rect 29570 145372 30322 145428
rect 30490 145372 31242 145428
rect 31410 145372 31702 145428
rect 31870 145372 32622 145428
rect 32790 145372 33542 145428
rect 33710 145372 34002 145428
rect 34170 145372 34922 145428
rect 35090 145372 35842 145428
rect 36010 145372 36302 145428
rect 36470 145372 37222 145428
rect 37390 145372 38142 145428
rect 38310 145372 38602 145428
rect 38770 145372 39522 145428
rect 39690 145372 39982 145428
rect 40150 145372 40902 145428
rect 41070 145372 41822 145428
rect 41990 145372 42282 145428
rect 42450 145372 43202 145428
rect 43370 145372 44122 145428
rect 44290 145372 44582 145428
rect 44750 145372 45502 145428
rect 45670 145372 46422 145428
rect 46590 145372 46882 145428
rect 47050 145372 47802 145428
rect 47970 145372 48722 145428
rect 48890 145372 49182 145428
rect 49350 145372 50102 145428
rect 50270 145372 51022 145428
rect 51190 145372 51482 145428
rect 51650 145372 52402 145428
rect 52570 145372 53322 145428
rect 53490 145372 53782 145428
rect 53950 145372 54702 145428
rect 54870 145372 55162 145428
rect 55330 145372 56082 145428
rect 56250 145372 57002 145428
rect 57170 145372 57462 145428
rect 57630 145372 58382 145428
rect 58550 145372 59302 145428
rect 59470 145372 59762 145428
rect 59930 145372 60682 145428
rect 60850 145372 61602 145428
rect 61770 145372 62062 145428
rect 62230 145372 62982 145428
rect 63150 145372 63902 145428
rect 64070 145372 64362 145428
rect 64530 145372 65282 145428
rect 65450 145372 66202 145428
rect 66370 145372 66662 145428
rect 66830 145372 67582 145428
rect 67750 145372 68042 145428
rect 68210 145372 68962 145428
rect 69130 145372 69882 145428
rect 70050 145372 70342 145428
rect 70510 145372 71262 145428
rect 71430 145372 72182 145428
rect 72350 145372 72642 145428
rect 72810 145372 73562 145428
rect 73730 145372 74482 145428
rect 74650 145372 74942 145428
rect 75110 145372 75862 145428
rect 76030 145372 76782 145428
rect 76950 145372 77242 145428
rect 77410 145372 78162 145428
rect 78330 145372 79082 145428
rect 79250 145372 79542 145428
rect 79710 145372 80462 145428
rect 80630 145372 81382 145428
rect 81550 145372 81842 145428
rect 82010 145372 82762 145428
rect 82930 145372 83222 145428
rect 83390 145372 84142 145428
rect 84310 145372 85062 145428
rect 85230 145372 85522 145428
rect 85690 145372 86442 145428
rect 86610 145372 87362 145428
rect 87530 145372 87822 145428
rect 87990 145372 88742 145428
rect 88910 145372 89662 145428
rect 89830 145372 90122 145428
rect 90290 145372 91042 145428
rect 91210 145372 91962 145428
rect 92130 145372 92422 145428
rect 92590 145372 93342 145428
rect 93510 145372 94262 145428
rect 94430 145372 94722 145428
rect 94890 145372 95642 145428
rect 95810 145372 96102 145428
rect 96270 145372 97022 145428
rect 97190 145372 97942 145428
rect 98110 145372 98402 145428
rect 98570 145372 99322 145428
rect 99490 145372 100242 145428
rect 100410 145372 100702 145428
rect 100870 145372 101622 145428
rect 101790 145372 102542 145428
rect 102710 145372 103002 145428
rect 103170 145372 103922 145428
rect 104090 145372 104842 145428
rect 105010 145372 105302 145428
rect 105470 145372 106222 145428
rect 106390 145372 107142 145428
rect 107310 145372 107602 145428
rect 107770 145372 108522 145428
rect 108690 145372 108982 145428
rect 109150 145372 109902 145428
rect 110070 145372 110822 145428
rect 110990 145372 111282 145428
rect 111450 145372 112202 145428
rect 112370 145372 113122 145428
rect 113290 145372 113582 145428
rect 113750 145372 114502 145428
rect 114670 145372 115422 145428
rect 115590 145372 115882 145428
rect 116050 145372 116802 145428
rect 116970 145372 117722 145428
rect 117890 145372 118182 145428
rect 118350 145372 119102 145428
rect 119270 145372 120022 145428
rect 120190 145372 120482 145428
rect 120650 145372 121402 145428
rect 121570 145372 122322 145428
rect 122490 145372 122782 145428
rect 122950 145372 123702 145428
rect 123870 145372 124162 145428
rect 124330 145372 125082 145428
rect 125250 145372 126002 145428
rect 126170 145372 126462 145428
rect 126630 145372 127382 145428
rect 127550 145372 128302 145428
rect 128470 145372 128762 145428
rect 128930 145372 129682 145428
rect 129850 145372 130602 145428
rect 130770 145372 131062 145428
rect 131230 145372 131982 145428
rect 132150 145372 132902 145428
rect 133070 145372 133362 145428
rect 133530 145372 134282 145428
rect 134450 145372 135202 145428
rect 135370 145372 135662 145428
rect 135830 145372 136582 145428
rect 136750 145372 137042 145428
rect 137210 145372 137962 145428
rect 138130 145372 138882 145428
rect 139050 145372 139342 145428
rect 139510 145372 140262 145428
rect 140430 145372 141182 145428
rect 141350 145372 141642 145428
rect 141810 145372 142562 145428
rect 142730 145372 143482 145428
rect 1124 856 143592 145372
rect 1124 800 1802 856
rect 1970 800 2262 856
rect 2430 800 3182 856
rect 3350 800 4102 856
rect 4270 800 4562 856
rect 4730 800 5482 856
rect 5650 800 6402 856
rect 6570 800 6862 856
rect 7030 800 7782 856
rect 7950 800 8702 856
rect 8870 800 9162 856
rect 9330 800 10082 856
rect 10250 800 11002 856
rect 11170 800 11462 856
rect 11630 800 12382 856
rect 12550 800 13302 856
rect 13470 800 13762 856
rect 13930 800 14682 856
rect 14850 800 15142 856
rect 15310 800 16062 856
rect 16230 800 16982 856
rect 17150 800 17442 856
rect 17610 800 18362 856
rect 18530 800 19282 856
rect 19450 800 19742 856
rect 19910 800 20662 856
rect 20830 800 21582 856
rect 21750 800 22042 856
rect 22210 800 22962 856
rect 23130 800 23882 856
rect 24050 800 24342 856
rect 24510 800 25262 856
rect 25430 800 26182 856
rect 26350 800 26642 856
rect 26810 800 27562 856
rect 27730 800 28022 856
rect 28190 800 28942 856
rect 29110 800 29862 856
rect 30030 800 30322 856
rect 30490 800 31242 856
rect 31410 800 32162 856
rect 32330 800 32622 856
rect 32790 800 33542 856
rect 33710 800 34462 856
rect 34630 800 34922 856
rect 35090 800 35842 856
rect 36010 800 36762 856
rect 36930 800 37222 856
rect 37390 800 38142 856
rect 38310 800 39062 856
rect 39230 800 39522 856
rect 39690 800 40442 856
rect 40610 800 41362 856
rect 41530 800 41822 856
rect 41990 800 42742 856
rect 42910 800 43202 856
rect 43370 800 44122 856
rect 44290 800 45042 856
rect 45210 800 45502 856
rect 45670 800 46422 856
rect 46590 800 47342 856
rect 47510 800 47802 856
rect 47970 800 48722 856
rect 48890 800 49642 856
rect 49810 800 50102 856
rect 50270 800 51022 856
rect 51190 800 51942 856
rect 52110 800 52402 856
rect 52570 800 53322 856
rect 53490 800 54242 856
rect 54410 800 54702 856
rect 54870 800 55622 856
rect 55790 800 56082 856
rect 56250 800 57002 856
rect 57170 800 57922 856
rect 58090 800 58382 856
rect 58550 800 59302 856
rect 59470 800 60222 856
rect 60390 800 60682 856
rect 60850 800 61602 856
rect 61770 800 62522 856
rect 62690 800 62982 856
rect 63150 800 63902 856
rect 64070 800 64822 856
rect 64990 800 65282 856
rect 65450 800 66202 856
rect 66370 800 67122 856
rect 67290 800 67582 856
rect 67750 800 68502 856
rect 68670 800 69422 856
rect 69590 800 69882 856
rect 70050 800 70802 856
rect 70970 800 71262 856
rect 71430 800 72182 856
rect 72350 800 73102 856
rect 73270 800 73562 856
rect 73730 800 74482 856
rect 74650 800 75402 856
rect 75570 800 75862 856
rect 76030 800 76782 856
rect 76950 800 77702 856
rect 77870 800 78162 856
rect 78330 800 79082 856
rect 79250 800 80002 856
rect 80170 800 80462 856
rect 80630 800 81382 856
rect 81550 800 82302 856
rect 82470 800 82762 856
rect 82930 800 83682 856
rect 83850 800 84142 856
rect 84310 800 85062 856
rect 85230 800 85982 856
rect 86150 800 86442 856
rect 86610 800 87362 856
rect 87530 800 88282 856
rect 88450 800 88742 856
rect 88910 800 89662 856
rect 89830 800 90582 856
rect 90750 800 91042 856
rect 91210 800 91962 856
rect 92130 800 92882 856
rect 93050 800 93342 856
rect 93510 800 94262 856
rect 94430 800 95182 856
rect 95350 800 95642 856
rect 95810 800 96562 856
rect 96730 800 97022 856
rect 97190 800 97942 856
rect 98110 800 98862 856
rect 99030 800 99322 856
rect 99490 800 100242 856
rect 100410 800 101162 856
rect 101330 800 101622 856
rect 101790 800 102542 856
rect 102710 800 103462 856
rect 103630 800 103922 856
rect 104090 800 104842 856
rect 105010 800 105762 856
rect 105930 800 106222 856
rect 106390 800 107142 856
rect 107310 800 108062 856
rect 108230 800 108522 856
rect 108690 800 109442 856
rect 109610 800 110362 856
rect 110530 800 110822 856
rect 110990 800 111742 856
rect 111910 800 112202 856
rect 112370 800 113122 856
rect 113290 800 114042 856
rect 114210 800 114502 856
rect 114670 800 115422 856
rect 115590 800 116342 856
rect 116510 800 116802 856
rect 116970 800 117722 856
rect 117890 800 118642 856
rect 118810 800 119102 856
rect 119270 800 120022 856
rect 120190 800 120942 856
rect 121110 800 121402 856
rect 121570 800 122322 856
rect 122490 800 123242 856
rect 123410 800 123702 856
rect 123870 800 124622 856
rect 124790 800 125082 856
rect 125250 800 126002 856
rect 126170 800 126922 856
rect 127090 800 127382 856
rect 127550 800 128302 856
rect 128470 800 129222 856
rect 129390 800 129682 856
rect 129850 800 130602 856
rect 130770 800 131522 856
rect 131690 800 131982 856
rect 132150 800 132902 856
rect 133070 800 133822 856
rect 133990 800 134282 856
rect 134450 800 135202 856
rect 135370 800 136122 856
rect 136290 800 136582 856
rect 136750 800 137502 856
rect 137670 800 138422 856
rect 138590 800 138882 856
rect 139050 800 139802 856
rect 139970 800 140262 856
rect 140430 800 141182 856
rect 141350 800 142102 856
rect 142270 800 142562 856
rect 142730 800 143482 856
<< metal3 >>
rect 0 144848 800 144968
rect 143284 144848 144084 144968
rect 0 143488 800 143608
rect 143284 143488 144084 143608
rect 0 142808 800 142928
rect 143284 142128 144084 142248
rect 0 141448 800 141568
rect 143284 141448 144084 141568
rect 0 140768 800 140888
rect 143284 140088 144084 140208
rect 0 139408 800 139528
rect 143284 138728 144084 138848
rect 0 138048 800 138168
rect 143284 138048 144084 138168
rect 0 137368 800 137488
rect 143284 136688 144084 136808
rect 0 136008 800 136128
rect 143284 135328 144084 135448
rect 0 134648 800 134768
rect 143284 134648 144084 134768
rect 0 133968 800 134088
rect 143284 133288 144084 133408
rect 0 132608 800 132728
rect 143284 132608 144084 132728
rect 0 131248 800 131368
rect 143284 131248 144084 131368
rect 0 130568 800 130688
rect 143284 129888 144084 130008
rect 0 129208 800 129328
rect 143284 129208 144084 129328
rect 0 127848 800 127968
rect 143284 127848 144084 127968
rect 0 127168 800 127288
rect 143284 126488 144084 126608
rect 0 125808 800 125928
rect 143284 125808 144084 125928
rect 0 124448 800 124568
rect 143284 124448 144084 124568
rect 0 123768 800 123888
rect 143284 123088 144084 123208
rect 0 122408 800 122528
rect 143284 122408 144084 122528
rect 0 121728 800 121848
rect 143284 121048 144084 121168
rect 0 120368 800 120488
rect 143284 119688 144084 119808
rect 0 119008 800 119128
rect 143284 119008 144084 119128
rect 0 118328 800 118448
rect 143284 117648 144084 117768
rect 0 116968 800 117088
rect 143284 116288 144084 116408
rect 0 115608 800 115728
rect 143284 115608 144084 115728
rect 0 114928 800 115048
rect 143284 114248 144084 114368
rect 0 113568 800 113688
rect 143284 113568 144084 113688
rect 0 112208 800 112328
rect 143284 112208 144084 112328
rect 0 111528 800 111648
rect 143284 110848 144084 110968
rect 0 110168 800 110288
rect 143284 110168 144084 110288
rect 0 108808 800 108928
rect 143284 108808 144084 108928
rect 0 108128 800 108248
rect 143284 107448 144084 107568
rect 0 106768 800 106888
rect 143284 106768 144084 106888
rect 0 105408 800 105528
rect 143284 105408 144084 105528
rect 0 104728 800 104848
rect 143284 104048 144084 104168
rect 0 103368 800 103488
rect 143284 103368 144084 103488
rect 0 102008 800 102128
rect 143284 102008 144084 102128
rect 0 101328 800 101448
rect 143284 100648 144084 100768
rect 0 99968 800 100088
rect 143284 99968 144084 100088
rect 0 99288 800 99408
rect 143284 98608 144084 98728
rect 0 97928 800 98048
rect 143284 97248 144084 97368
rect 0 96568 800 96688
rect 143284 96568 144084 96688
rect 0 95888 800 96008
rect 143284 95208 144084 95328
rect 0 94528 800 94648
rect 143284 94528 144084 94648
rect 0 93168 800 93288
rect 143284 93168 144084 93288
rect 0 92488 800 92608
rect 143284 91808 144084 91928
rect 0 91128 800 91248
rect 143284 91128 144084 91248
rect 0 89768 800 89888
rect 143284 89768 144084 89888
rect 0 89088 800 89208
rect 143284 88408 144084 88528
rect 0 87728 800 87848
rect 143284 87728 144084 87848
rect 0 86368 800 86488
rect 143284 86368 144084 86488
rect 0 85688 800 85808
rect 143284 85008 144084 85128
rect 0 84328 800 84448
rect 143284 84328 144084 84448
rect 0 82968 800 83088
rect 143284 82968 144084 83088
rect 0 82288 800 82408
rect 143284 81608 144084 81728
rect 0 80928 800 81048
rect 143284 80928 144084 81048
rect 0 80248 800 80368
rect 143284 79568 144084 79688
rect 0 78888 800 79008
rect 143284 78208 144084 78328
rect 0 77528 800 77648
rect 143284 77528 144084 77648
rect 0 76848 800 76968
rect 143284 76168 144084 76288
rect 0 75488 800 75608
rect 143284 74808 144084 74928
rect 0 74128 800 74248
rect 143284 74128 144084 74248
rect 0 73448 800 73568
rect 143284 72768 144084 72888
rect 0 72088 800 72208
rect 143284 72088 144084 72208
rect 0 70728 800 70848
rect 143284 70728 144084 70848
rect 0 70048 800 70168
rect 143284 69368 144084 69488
rect 0 68688 800 68808
rect 143284 68688 144084 68808
rect 0 67328 800 67448
rect 143284 67328 144084 67448
rect 0 66648 800 66768
rect 143284 65968 144084 66088
rect 0 65288 800 65408
rect 143284 65288 144084 65408
rect 0 63928 800 64048
rect 143284 63928 144084 64048
rect 0 63248 800 63368
rect 143284 62568 144084 62688
rect 0 61888 800 62008
rect 143284 61888 144084 62008
rect 0 61208 800 61328
rect 143284 60528 144084 60648
rect 0 59848 800 59968
rect 143284 59168 144084 59288
rect 0 58488 800 58608
rect 143284 58488 144084 58608
rect 0 57808 800 57928
rect 143284 57128 144084 57248
rect 0 56448 800 56568
rect 143284 55768 144084 55888
rect 0 55088 800 55208
rect 143284 55088 144084 55208
rect 0 54408 800 54528
rect 143284 53728 144084 53848
rect 0 53048 800 53168
rect 143284 53048 144084 53168
rect 0 51688 800 51808
rect 143284 51688 144084 51808
rect 0 51008 800 51128
rect 143284 50328 144084 50448
rect 0 49648 800 49768
rect 143284 49648 144084 49768
rect 0 48288 800 48408
rect 143284 48288 144084 48408
rect 0 47608 800 47728
rect 143284 46928 144084 47048
rect 0 46248 800 46368
rect 143284 46248 144084 46368
rect 0 44888 800 45008
rect 143284 44888 144084 45008
rect 0 44208 800 44328
rect 143284 43528 144084 43648
rect 0 42848 800 42968
rect 143284 42848 144084 42968
rect 0 41488 800 41608
rect 143284 41488 144084 41608
rect 0 40808 800 40928
rect 143284 40128 144084 40248
rect 0 39448 800 39568
rect 143284 39448 144084 39568
rect 0 38768 800 38888
rect 143284 38088 144084 38208
rect 0 37408 800 37528
rect 143284 36728 144084 36848
rect 0 36048 800 36168
rect 143284 36048 144084 36168
rect 0 35368 800 35488
rect 143284 34688 144084 34808
rect 0 34008 800 34128
rect 143284 33328 144084 33448
rect 0 32648 800 32768
rect 143284 32648 144084 32768
rect 0 31968 800 32088
rect 143284 31288 144084 31408
rect 0 30608 800 30728
rect 143284 30608 144084 30728
rect 0 29248 800 29368
rect 143284 29248 144084 29368
rect 0 28568 800 28688
rect 143284 27888 144084 28008
rect 0 27208 800 27328
rect 143284 27208 144084 27328
rect 0 25848 800 25968
rect 143284 25848 144084 25968
rect 0 25168 800 25288
rect 143284 24488 144084 24608
rect 0 23808 800 23928
rect 143284 23808 144084 23928
rect 0 22448 800 22568
rect 143284 22448 144084 22568
rect 0 21768 800 21888
rect 143284 21088 144084 21208
rect 0 20408 800 20528
rect 143284 20408 144084 20528
rect 0 19728 800 19848
rect 143284 19048 144084 19168
rect 0 18368 800 18488
rect 143284 17688 144084 17808
rect 0 17008 800 17128
rect 143284 17008 144084 17128
rect 0 16328 800 16448
rect 143284 15648 144084 15768
rect 0 14968 800 15088
rect 143284 14288 144084 14408
rect 0 13608 800 13728
rect 143284 13608 144084 13728
rect 0 12928 800 13048
rect 143284 12248 144084 12368
rect 0 11568 800 11688
rect 143284 11568 144084 11688
rect 0 10208 800 10328
rect 143284 10208 144084 10328
rect 0 9528 800 9648
rect 143284 8848 144084 8968
rect 0 8168 800 8288
rect 143284 8168 144084 8288
rect 0 6808 800 6928
rect 143284 6808 144084 6928
rect 0 6128 800 6248
rect 143284 5448 144084 5568
rect 0 4768 800 4888
rect 143284 4768 144084 4888
rect 0 3408 800 3528
rect 143284 3408 144084 3528
rect 0 2728 800 2848
rect 143284 2048 144084 2168
rect 0 1368 800 1488
rect 143284 1368 144084 1488
<< obsm3 >>
rect 880 144768 143204 144941
rect 800 143688 143284 144768
rect 880 143408 143204 143688
rect 800 143008 143284 143408
rect 880 142728 143284 143008
rect 800 142328 143284 142728
rect 800 142048 143204 142328
rect 800 141648 143284 142048
rect 880 141368 143204 141648
rect 800 140968 143284 141368
rect 880 140688 143284 140968
rect 800 140288 143284 140688
rect 800 140008 143204 140288
rect 800 139608 143284 140008
rect 880 139328 143284 139608
rect 800 138928 143284 139328
rect 800 138648 143204 138928
rect 800 138248 143284 138648
rect 880 137968 143204 138248
rect 800 137568 143284 137968
rect 880 137288 143284 137568
rect 800 136888 143284 137288
rect 800 136608 143204 136888
rect 800 136208 143284 136608
rect 880 135928 143284 136208
rect 800 135528 143284 135928
rect 800 135248 143204 135528
rect 800 134848 143284 135248
rect 880 134568 143204 134848
rect 800 134168 143284 134568
rect 880 133888 143284 134168
rect 800 133488 143284 133888
rect 800 133208 143204 133488
rect 800 132808 143284 133208
rect 880 132528 143204 132808
rect 800 131448 143284 132528
rect 880 131168 143204 131448
rect 800 130768 143284 131168
rect 880 130488 143284 130768
rect 800 130088 143284 130488
rect 800 129808 143204 130088
rect 800 129408 143284 129808
rect 880 129128 143204 129408
rect 800 128048 143284 129128
rect 880 127768 143204 128048
rect 800 127368 143284 127768
rect 880 127088 143284 127368
rect 800 126688 143284 127088
rect 800 126408 143204 126688
rect 800 126008 143284 126408
rect 880 125728 143204 126008
rect 800 124648 143284 125728
rect 880 124368 143204 124648
rect 800 123968 143284 124368
rect 880 123688 143284 123968
rect 800 123288 143284 123688
rect 800 123008 143204 123288
rect 800 122608 143284 123008
rect 880 122328 143204 122608
rect 800 121928 143284 122328
rect 880 121648 143284 121928
rect 800 121248 143284 121648
rect 800 120968 143204 121248
rect 800 120568 143284 120968
rect 880 120288 143284 120568
rect 800 119888 143284 120288
rect 800 119608 143204 119888
rect 800 119208 143284 119608
rect 880 118928 143204 119208
rect 800 118528 143284 118928
rect 880 118248 143284 118528
rect 800 117848 143284 118248
rect 800 117568 143204 117848
rect 800 117168 143284 117568
rect 880 116888 143284 117168
rect 800 116488 143284 116888
rect 800 116208 143204 116488
rect 800 115808 143284 116208
rect 880 115528 143204 115808
rect 800 115128 143284 115528
rect 880 114848 143284 115128
rect 800 114448 143284 114848
rect 800 114168 143204 114448
rect 800 113768 143284 114168
rect 880 113488 143204 113768
rect 800 112408 143284 113488
rect 880 112128 143204 112408
rect 800 111728 143284 112128
rect 880 111448 143284 111728
rect 800 111048 143284 111448
rect 800 110768 143204 111048
rect 800 110368 143284 110768
rect 880 110088 143204 110368
rect 800 109008 143284 110088
rect 880 108728 143204 109008
rect 800 108328 143284 108728
rect 880 108048 143284 108328
rect 800 107648 143284 108048
rect 800 107368 143204 107648
rect 800 106968 143284 107368
rect 880 106688 143204 106968
rect 800 105608 143284 106688
rect 880 105328 143204 105608
rect 800 104928 143284 105328
rect 880 104648 143284 104928
rect 800 104248 143284 104648
rect 800 103968 143204 104248
rect 800 103568 143284 103968
rect 880 103288 143204 103568
rect 800 102208 143284 103288
rect 880 101928 143204 102208
rect 800 101528 143284 101928
rect 880 101248 143284 101528
rect 800 100848 143284 101248
rect 800 100568 143204 100848
rect 800 100168 143284 100568
rect 880 99888 143204 100168
rect 800 99488 143284 99888
rect 880 99208 143284 99488
rect 800 98808 143284 99208
rect 800 98528 143204 98808
rect 800 98128 143284 98528
rect 880 97848 143284 98128
rect 800 97448 143284 97848
rect 800 97168 143204 97448
rect 800 96768 143284 97168
rect 880 96488 143204 96768
rect 800 96088 143284 96488
rect 880 95808 143284 96088
rect 800 95408 143284 95808
rect 800 95128 143204 95408
rect 800 94728 143284 95128
rect 880 94448 143204 94728
rect 800 93368 143284 94448
rect 880 93088 143204 93368
rect 800 92688 143284 93088
rect 880 92408 143284 92688
rect 800 92008 143284 92408
rect 800 91728 143204 92008
rect 800 91328 143284 91728
rect 880 91048 143204 91328
rect 800 89968 143284 91048
rect 880 89688 143204 89968
rect 800 89288 143284 89688
rect 880 89008 143284 89288
rect 800 88608 143284 89008
rect 800 88328 143204 88608
rect 800 87928 143284 88328
rect 880 87648 143204 87928
rect 800 86568 143284 87648
rect 880 86288 143204 86568
rect 800 85888 143284 86288
rect 880 85608 143284 85888
rect 800 85208 143284 85608
rect 800 84928 143204 85208
rect 800 84528 143284 84928
rect 880 84248 143204 84528
rect 800 83168 143284 84248
rect 880 82888 143204 83168
rect 800 82488 143284 82888
rect 880 82208 143284 82488
rect 800 81808 143284 82208
rect 800 81528 143204 81808
rect 800 81128 143284 81528
rect 880 80848 143204 81128
rect 800 80448 143284 80848
rect 880 80168 143284 80448
rect 800 79768 143284 80168
rect 800 79488 143204 79768
rect 800 79088 143284 79488
rect 880 78808 143284 79088
rect 800 78408 143284 78808
rect 800 78128 143204 78408
rect 800 77728 143284 78128
rect 880 77448 143204 77728
rect 800 77048 143284 77448
rect 880 76768 143284 77048
rect 800 76368 143284 76768
rect 800 76088 143204 76368
rect 800 75688 143284 76088
rect 880 75408 143284 75688
rect 800 75008 143284 75408
rect 800 74728 143204 75008
rect 800 74328 143284 74728
rect 880 74048 143204 74328
rect 800 73648 143284 74048
rect 880 73368 143284 73648
rect 800 72968 143284 73368
rect 800 72688 143204 72968
rect 800 72288 143284 72688
rect 880 72008 143204 72288
rect 800 70928 143284 72008
rect 880 70648 143204 70928
rect 800 70248 143284 70648
rect 880 69968 143284 70248
rect 800 69568 143284 69968
rect 800 69288 143204 69568
rect 800 68888 143284 69288
rect 880 68608 143204 68888
rect 800 67528 143284 68608
rect 880 67248 143204 67528
rect 800 66848 143284 67248
rect 880 66568 143284 66848
rect 800 66168 143284 66568
rect 800 65888 143204 66168
rect 800 65488 143284 65888
rect 880 65208 143204 65488
rect 800 64128 143284 65208
rect 880 63848 143204 64128
rect 800 63448 143284 63848
rect 880 63168 143284 63448
rect 800 62768 143284 63168
rect 800 62488 143204 62768
rect 800 62088 143284 62488
rect 880 61808 143204 62088
rect 800 61408 143284 61808
rect 880 61128 143284 61408
rect 800 60728 143284 61128
rect 800 60448 143204 60728
rect 800 60048 143284 60448
rect 880 59768 143284 60048
rect 800 59368 143284 59768
rect 800 59088 143204 59368
rect 800 58688 143284 59088
rect 880 58408 143204 58688
rect 800 58008 143284 58408
rect 880 57728 143284 58008
rect 800 57328 143284 57728
rect 800 57048 143204 57328
rect 800 56648 143284 57048
rect 880 56368 143284 56648
rect 800 55968 143284 56368
rect 800 55688 143204 55968
rect 800 55288 143284 55688
rect 880 55008 143204 55288
rect 800 54608 143284 55008
rect 880 54328 143284 54608
rect 800 53928 143284 54328
rect 800 53648 143204 53928
rect 800 53248 143284 53648
rect 880 52968 143204 53248
rect 800 51888 143284 52968
rect 880 51608 143204 51888
rect 800 51208 143284 51608
rect 880 50928 143284 51208
rect 800 50528 143284 50928
rect 800 50248 143204 50528
rect 800 49848 143284 50248
rect 880 49568 143204 49848
rect 800 48488 143284 49568
rect 880 48208 143204 48488
rect 800 47808 143284 48208
rect 880 47528 143284 47808
rect 800 47128 143284 47528
rect 800 46848 143204 47128
rect 800 46448 143284 46848
rect 880 46168 143204 46448
rect 800 45088 143284 46168
rect 880 44808 143204 45088
rect 800 44408 143284 44808
rect 880 44128 143284 44408
rect 800 43728 143284 44128
rect 800 43448 143204 43728
rect 800 43048 143284 43448
rect 880 42768 143204 43048
rect 800 41688 143284 42768
rect 880 41408 143204 41688
rect 800 41008 143284 41408
rect 880 40728 143284 41008
rect 800 40328 143284 40728
rect 800 40048 143204 40328
rect 800 39648 143284 40048
rect 880 39368 143204 39648
rect 800 38968 143284 39368
rect 880 38688 143284 38968
rect 800 38288 143284 38688
rect 800 38008 143204 38288
rect 800 37608 143284 38008
rect 880 37328 143284 37608
rect 800 36928 143284 37328
rect 800 36648 143204 36928
rect 800 36248 143284 36648
rect 880 35968 143204 36248
rect 800 35568 143284 35968
rect 880 35288 143284 35568
rect 800 34888 143284 35288
rect 800 34608 143204 34888
rect 800 34208 143284 34608
rect 880 33928 143284 34208
rect 800 33528 143284 33928
rect 800 33248 143204 33528
rect 800 32848 143284 33248
rect 880 32568 143204 32848
rect 800 32168 143284 32568
rect 880 31888 143284 32168
rect 800 31488 143284 31888
rect 800 31208 143204 31488
rect 800 30808 143284 31208
rect 880 30528 143204 30808
rect 800 29448 143284 30528
rect 880 29168 143204 29448
rect 800 28768 143284 29168
rect 880 28488 143284 28768
rect 800 28088 143284 28488
rect 800 27808 143204 28088
rect 800 27408 143284 27808
rect 880 27128 143204 27408
rect 800 26048 143284 27128
rect 880 25768 143204 26048
rect 800 25368 143284 25768
rect 880 25088 143284 25368
rect 800 24688 143284 25088
rect 800 24408 143204 24688
rect 800 24008 143284 24408
rect 880 23728 143204 24008
rect 800 22648 143284 23728
rect 880 22368 143204 22648
rect 800 21968 143284 22368
rect 880 21688 143284 21968
rect 800 21288 143284 21688
rect 800 21008 143204 21288
rect 800 20608 143284 21008
rect 880 20328 143204 20608
rect 800 19928 143284 20328
rect 880 19648 143284 19928
rect 800 19248 143284 19648
rect 800 18968 143204 19248
rect 800 18568 143284 18968
rect 880 18288 143284 18568
rect 800 17888 143284 18288
rect 800 17608 143204 17888
rect 800 17208 143284 17608
rect 880 16928 143204 17208
rect 800 16528 143284 16928
rect 880 16248 143284 16528
rect 800 15848 143284 16248
rect 800 15568 143204 15848
rect 800 15168 143284 15568
rect 880 14888 143284 15168
rect 800 14488 143284 14888
rect 800 14208 143204 14488
rect 800 13808 143284 14208
rect 880 13528 143204 13808
rect 800 13128 143284 13528
rect 880 12848 143284 13128
rect 800 12448 143284 12848
rect 800 12168 143204 12448
rect 800 11768 143284 12168
rect 880 11488 143204 11768
rect 800 10408 143284 11488
rect 880 10128 143204 10408
rect 800 9728 143284 10128
rect 880 9448 143284 9728
rect 800 9048 143284 9448
rect 800 8768 143204 9048
rect 800 8368 143284 8768
rect 880 8088 143204 8368
rect 800 7008 143284 8088
rect 880 6728 143204 7008
rect 800 6328 143284 6728
rect 880 6048 143284 6328
rect 800 5648 143284 6048
rect 800 5368 143204 5648
rect 800 4968 143284 5368
rect 880 4688 143204 4968
rect 800 3608 143284 4688
rect 880 3328 143204 3608
rect 800 2928 143284 3328
rect 880 2648 143284 2928
rect 800 2248 143284 2648
rect 800 1968 143204 2248
rect 800 1568 143284 1968
rect 880 1395 143204 1568
<< metal4 >>
rect -8576 -7504 -7976 153296
rect -7636 -6564 -7036 152356
rect -6696 -5624 -6096 151416
rect -5756 -4684 -5156 150476
rect -4816 -3744 -4216 149536
rect -3876 -2804 -3276 148596
rect -2936 -1864 -2336 147656
rect -1996 -924 -1396 146716
rect 804 -1864 1404 147656
rect 4404 -3744 5004 149536
rect 8004 -5624 8604 151416
rect 11604 -7504 12204 153296
rect 18804 -1864 19404 147656
rect 22404 -3744 23004 149536
rect 26004 -5624 26604 151416
rect 29604 -7504 30204 153296
rect 36804 -1864 37404 147656
rect 40404 -3744 41004 149536
rect 44004 -5624 44604 151416
rect 47604 -7504 48204 153296
rect 54804 -1864 55404 147656
rect 58404 -3744 59004 149536
rect 62004 -5624 62604 151416
rect 65604 -7504 66204 153296
rect 72804 -1864 73404 147656
rect 76404 -3744 77004 149536
rect 80004 -5624 80604 151416
rect 83604 -7504 84204 153296
rect 90804 -1864 91404 147656
rect 94404 -3744 95004 149536
rect 98004 -5624 98604 151416
rect 101604 -7504 102204 153296
rect 108804 -1864 109404 147656
rect 112404 -3744 113004 149536
rect 116004 -5624 116604 151416
rect 119604 -7504 120204 153296
rect 126804 -1864 127404 147656
rect 130404 -3744 131004 149536
rect 134004 -5624 134604 151416
rect 137604 -7504 138204 153296
rect 145468 -924 146068 146716
rect 146408 -1864 147008 147656
rect 147348 -2804 147948 148596
rect 148288 -3744 148888 149536
rect 149228 -4684 149828 150476
rect 150168 -5624 150768 151416
rect 151108 -6564 151708 152356
rect 152048 -7504 152648 153296
<< obsm4 >>
rect 5947 3435 7924 141813
rect 8684 3435 11524 141813
rect 12284 3435 18724 141813
rect 19484 3435 22324 141813
rect 23084 3435 25924 141813
rect 26684 3435 29524 141813
rect 30284 3435 36724 141813
rect 37484 3435 40324 141813
rect 41084 3435 43924 141813
rect 44684 3435 47524 141813
rect 48284 3435 54724 141813
rect 55484 3435 58324 141813
rect 59084 3435 61924 141813
rect 62684 3435 65524 141813
rect 66284 3435 72724 141813
rect 73484 3435 76324 141813
rect 77084 3435 79924 141813
rect 80684 3435 83524 141813
rect 84284 3435 90724 141813
rect 91484 3435 94324 141813
rect 95084 3435 97924 141813
rect 98684 3435 101524 141813
rect 102284 3435 106661 141813
<< metal5 >>
rect -8576 152696 152648 153296
rect -7636 151756 151708 152356
rect -6696 150816 150768 151416
rect -5756 149876 149828 150476
rect -4816 148936 148888 149536
rect -3876 147996 147948 148596
rect -2936 147056 147008 147656
rect -1996 146116 146068 146716
rect -8576 138676 152648 139276
rect -6696 135076 150768 135676
rect -4816 131476 148888 132076
rect -2936 127828 147008 128428
rect -8576 120676 152648 121276
rect -6696 117076 150768 117676
rect -4816 113476 148888 114076
rect -2936 109828 147008 110428
rect -8576 102676 152648 103276
rect -6696 99076 150768 99676
rect -4816 95476 148888 96076
rect -2936 91828 147008 92428
rect -8576 84676 152648 85276
rect -6696 81076 150768 81676
rect -4816 77476 148888 78076
rect -2936 73828 147008 74428
rect -8576 66676 152648 67276
rect -6696 63076 150768 63676
rect -4816 59476 148888 60076
rect -2936 55828 147008 56428
rect -8576 48676 152648 49276
rect -6696 45076 150768 45676
rect -4816 41476 148888 42076
rect -2936 37828 147008 38428
rect -8576 30676 152648 31276
rect -6696 27076 150768 27676
rect -4816 23476 148888 24076
rect -2936 19828 147008 20428
rect -8576 12676 152648 13276
rect -6696 9076 150768 9676
rect -4816 5476 148888 6076
rect -2936 1828 147008 2428
rect -1996 -924 146068 -324
rect -2936 -1864 147008 -1264
rect -3876 -2804 147948 -2204
rect -4816 -3744 148888 -3144
rect -5756 -4684 149828 -4084
rect -6696 -5624 150768 -5024
rect -7636 -6564 151708 -5964
rect -8576 -7504 152648 -6904
<< obsm5 >>
rect -8576 153296 -7976 153298
rect 29604 153296 30204 153298
rect 65604 153296 66204 153298
rect 101604 153296 102204 153298
rect 137604 153296 138204 153298
rect 152048 153296 152648 153298
rect -8576 152694 -7976 152696
rect 29604 152694 30204 152696
rect 65604 152694 66204 152696
rect 101604 152694 102204 152696
rect 137604 152694 138204 152696
rect 152048 152694 152648 152696
rect -7636 152356 -7036 152358
rect 11604 152356 12204 152358
rect 47604 152356 48204 152358
rect 83604 152356 84204 152358
rect 119604 152356 120204 152358
rect 151108 152356 151708 152358
rect -7636 151754 -7036 151756
rect 11604 151754 12204 151756
rect 47604 151754 48204 151756
rect 83604 151754 84204 151756
rect 119604 151754 120204 151756
rect 151108 151754 151708 151756
rect -6696 151416 -6096 151418
rect 26004 151416 26604 151418
rect 62004 151416 62604 151418
rect 98004 151416 98604 151418
rect 134004 151416 134604 151418
rect 150168 151416 150768 151418
rect -6696 150814 -6096 150816
rect 26004 150814 26604 150816
rect 62004 150814 62604 150816
rect 98004 150814 98604 150816
rect 134004 150814 134604 150816
rect 150168 150814 150768 150816
rect -5756 150476 -5156 150478
rect 8004 150476 8604 150478
rect 44004 150476 44604 150478
rect 80004 150476 80604 150478
rect 116004 150476 116604 150478
rect 149228 150476 149828 150478
rect -5756 149874 -5156 149876
rect 8004 149874 8604 149876
rect 44004 149874 44604 149876
rect 80004 149874 80604 149876
rect 116004 149874 116604 149876
rect 149228 149874 149828 149876
rect -4816 149536 -4216 149538
rect 22404 149536 23004 149538
rect 58404 149536 59004 149538
rect 94404 149536 95004 149538
rect 130404 149536 131004 149538
rect 148288 149536 148888 149538
rect -4816 148934 -4216 148936
rect 22404 148934 23004 148936
rect 58404 148934 59004 148936
rect 94404 148934 95004 148936
rect 130404 148934 131004 148936
rect 148288 148934 148888 148936
rect -3876 148596 -3276 148598
rect 4404 148596 5004 148598
rect 40404 148596 41004 148598
rect 76404 148596 77004 148598
rect 112404 148596 113004 148598
rect 147348 148596 147948 148598
rect -3876 147994 -3276 147996
rect 4404 147994 5004 147996
rect 40404 147994 41004 147996
rect 76404 147994 77004 147996
rect 112404 147994 113004 147996
rect 147348 147994 147948 147996
rect -2936 147656 -2336 147658
rect 18804 147656 19404 147658
rect 54804 147656 55404 147658
rect 90804 147656 91404 147658
rect 126804 147656 127404 147658
rect 146408 147656 147008 147658
rect -2936 147054 -2336 147056
rect 18804 147054 19404 147056
rect 54804 147054 55404 147056
rect 90804 147054 91404 147056
rect 126804 147054 127404 147056
rect 146408 147054 147008 147056
rect -1996 146716 -1396 146718
rect 804 146716 1404 146718
rect 36804 146716 37404 146718
rect 72804 146716 73404 146718
rect 108804 146716 109404 146718
rect 145468 146716 146068 146718
rect -1996 146114 -1396 146116
rect 145468 146114 146068 146116
rect 0 139596 144084 145796
rect -8576 139276 -7976 139278
rect 152048 139276 152648 139278
rect -8576 138674 -7976 138676
rect 152048 138674 152648 138676
rect 0 135996 144084 138356
rect -6696 135676 -6096 135678
rect 150168 135676 150768 135678
rect -6696 135074 -6096 135076
rect 150168 135074 150768 135076
rect 0 132396 144084 134756
rect -4816 132076 -4216 132078
rect 148288 132076 148888 132078
rect -4816 131474 -4216 131476
rect 148288 131474 148888 131476
rect 0 128748 144084 131156
rect -2936 128428 -2336 128430
rect 146408 128428 147008 128430
rect -2936 127826 -2336 127828
rect 146408 127826 147008 127828
rect 0 121596 144084 127508
rect -7636 121276 -7036 121278
rect 151108 121276 151708 121278
rect -7636 120674 -7036 120676
rect 151108 120674 151708 120676
rect 0 117996 144084 120356
rect -5756 117676 -5156 117678
rect 149228 117676 149828 117678
rect -5756 117074 -5156 117076
rect 149228 117074 149828 117076
rect 0 114396 144084 116756
rect -3876 114076 -3276 114078
rect 147348 114076 147948 114078
rect -3876 113474 -3276 113476
rect 147348 113474 147948 113476
rect 0 110748 144084 113156
rect -1996 110428 -1396 110430
rect 145468 110428 146068 110430
rect -1996 109826 -1396 109828
rect 145468 109826 146068 109828
rect 0 103596 144084 109508
rect -8576 103276 -7976 103278
rect 152048 103276 152648 103278
rect -8576 102674 -7976 102676
rect 152048 102674 152648 102676
rect 0 99996 144084 102356
rect -6696 99676 -6096 99678
rect 150168 99676 150768 99678
rect -6696 99074 -6096 99076
rect 150168 99074 150768 99076
rect 0 96396 144084 98756
rect -4816 96076 -4216 96078
rect 148288 96076 148888 96078
rect -4816 95474 -4216 95476
rect 148288 95474 148888 95476
rect 0 92748 144084 95156
rect -2936 92428 -2336 92430
rect 146408 92428 147008 92430
rect -2936 91826 -2336 91828
rect 146408 91826 147008 91828
rect 0 85596 144084 91508
rect -7636 85276 -7036 85278
rect 151108 85276 151708 85278
rect -7636 84674 -7036 84676
rect 151108 84674 151708 84676
rect 0 81996 144084 84356
rect -5756 81676 -5156 81678
rect 149228 81676 149828 81678
rect -5756 81074 -5156 81076
rect 149228 81074 149828 81076
rect 0 78396 144084 80756
rect -3876 78076 -3276 78078
rect 147348 78076 147948 78078
rect -3876 77474 -3276 77476
rect 147348 77474 147948 77476
rect 0 74748 144084 77156
rect -1996 74428 -1396 74430
rect 145468 74428 146068 74430
rect -1996 73826 -1396 73828
rect 145468 73826 146068 73828
rect 0 67596 144084 73508
rect -8576 67276 -7976 67278
rect 152048 67276 152648 67278
rect -8576 66674 -7976 66676
rect 152048 66674 152648 66676
rect 0 63996 144084 66356
rect -6696 63676 -6096 63678
rect 150168 63676 150768 63678
rect -6696 63074 -6096 63076
rect 150168 63074 150768 63076
rect 0 60396 144084 62756
rect -4816 60076 -4216 60078
rect 148288 60076 148888 60078
rect -4816 59474 -4216 59476
rect 148288 59474 148888 59476
rect 0 56748 144084 59156
rect -2936 56428 -2336 56430
rect 146408 56428 147008 56430
rect -2936 55826 -2336 55828
rect 146408 55826 147008 55828
rect 0 49596 144084 55508
rect -7636 49276 -7036 49278
rect 151108 49276 151708 49278
rect -7636 48674 -7036 48676
rect 151108 48674 151708 48676
rect 0 45996 144084 48356
rect -5756 45676 -5156 45678
rect 149228 45676 149828 45678
rect -5756 45074 -5156 45076
rect 149228 45074 149828 45076
rect 0 42396 144084 44756
rect -3876 42076 -3276 42078
rect 147348 42076 147948 42078
rect -3876 41474 -3276 41476
rect 147348 41474 147948 41476
rect 0 38748 144084 41156
rect -1996 38428 -1396 38430
rect 145468 38428 146068 38430
rect -1996 37826 -1396 37828
rect 145468 37826 146068 37828
rect 0 31596 144084 37508
rect -8576 31276 -7976 31278
rect 152048 31276 152648 31278
rect -8576 30674 -7976 30676
rect 152048 30674 152648 30676
rect 0 27996 144084 30356
rect -6696 27676 -6096 27678
rect 150168 27676 150768 27678
rect -6696 27074 -6096 27076
rect 150168 27074 150768 27076
rect 0 24396 144084 26756
rect -4816 24076 -4216 24078
rect 148288 24076 148888 24078
rect -4816 23474 -4216 23476
rect 148288 23474 148888 23476
rect 0 20748 144084 23156
rect -2936 20428 -2336 20430
rect 146408 20428 147008 20430
rect -2936 19826 -2336 19828
rect 146408 19826 147008 19828
rect 0 13596 144084 19508
rect -7636 13276 -7036 13278
rect 151108 13276 151708 13278
rect -7636 12674 -7036 12676
rect 151108 12674 151708 12676
rect 0 9996 144084 12356
rect -5756 9676 -5156 9678
rect 149228 9676 149828 9678
rect -5756 9074 -5156 9076
rect 149228 9074 149828 9076
rect 0 6396 144084 8756
rect -3876 6076 -3276 6078
rect 147348 6076 147948 6078
rect -3876 5474 -3276 5476
rect 147348 5474 147948 5476
rect 0 2748 144084 5156
rect -1996 2428 -1396 2430
rect 145468 2428 146068 2430
rect -1996 1826 -1396 1828
rect 145468 1826 146068 1828
rect 0 0 144084 1508
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 145468 -324 146068 -322
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 145468 -926 146068 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 146408 -1264 147008 -1262
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 146408 -1866 147008 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 147348 -2204 147948 -2202
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 147348 -2806 147948 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 148288 -3144 148888 -3142
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 148288 -3746 148888 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 149228 -4084 149828 -4082
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 149228 -4686 149828 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 150168 -5024 150768 -5022
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 150168 -5626 150768 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 151108 -5964 151708 -5962
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 151108 -6566 151708 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 152048 -6904 152648 -6902
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 152048 -7506 152648 -7504
<< labels >>
rlabel metal2 s 3698 145428 3754 146228 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 143284 112208 144084 112328 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 111798 0 111854 800 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal3 s 0 139408 800 139528 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal3 s 143284 114248 144084 114368 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 128358 0 128414 800 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal3 s 0 104728 800 104848 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 6918 0 6974 800 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 97998 0 98054 800 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal2 s 77758 0 77814 800 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 87418 145428 87474 146228 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal2 s 135258 0 135314 800 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 0 1368 800 1488 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal2 s 85118 0 85174 800 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 143284 59168 144084 59288 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 94778 145428 94834 146228 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal2 s 88338 0 88394 800 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal2 s 107658 145428 107714 146228 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal2 s 8758 0 8814 800 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 0 47608 800 47728 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 143284 94528 144084 94648 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 0 63248 800 63368 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 143284 134648 144084 134768 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal2 s 91098 0 91154 800 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 0 140768 800 140888 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal2 s 41418 0 41474 800 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal2 s 68558 0 68614 800 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 116858 145428 116914 146228 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal3 s 143284 74808 144084 74928 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal2 s 129738 0 129794 800 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 io_in[10]
port 31 nsew signal input
rlabel metal2 s 134338 145428 134394 146228 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 io_in[12]
port 33 nsew signal input
rlabel metal2 s 50158 145428 50214 146228 6 io_in[13]
port 34 nsew signal input
rlabel metal2 s 25778 145428 25834 146228 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 io_in[15]
port 36 nsew signal input
rlabel metal3 s 0 92488 800 92608 6 io_in[16]
port 37 nsew signal input
rlabel metal3 s 143284 85008 144084 85128 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 128818 145428 128874 146228 6 io_in[18]
port 39 nsew signal input
rlabel metal3 s 143284 2048 144084 2168 6 io_in[19]
port 40 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 84198 145428 84254 146228 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 88798 145428 88854 146228 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 54758 145428 54814 146228 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 io_in[24]
port 46 nsew signal input
rlabel metal3 s 143284 68688 144084 68808 6 io_in[25]
port 47 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 io_in[26]
port 48 nsew signal input
rlabel metal2 s 37278 145428 37334 146228 6 io_in[27]
port 49 nsew signal input
rlabel metal2 s 38198 145428 38254 146228 6 io_in[28]
port 50 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 io_in[29]
port 51 nsew signal input
rlabel metal2 s 120078 145428 120134 146228 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s 143284 12248 144084 12368 6 io_in[30]
port 53 nsew signal input
rlabel metal3 s 143284 8168 144084 8288 6 io_in[31]
port 54 nsew signal input
rlabel metal2 s 11518 145428 11574 146228 6 io_in[32]
port 55 nsew signal input
rlabel metal3 s 0 144848 800 144968 6 io_in[33]
port 56 nsew signal input
rlabel metal3 s 143284 107448 144084 107568 6 io_in[34]
port 57 nsew signal input
rlabel metal2 s 140318 0 140374 800 6 io_in[35]
port 58 nsew signal input
rlabel metal2 s 67638 145428 67694 146228 6 io_in[36]
port 59 nsew signal input
rlabel metal2 s 18878 145428 18934 146228 6 io_in[37]
port 60 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 io_in[3]
port 61 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 143284 23808 144084 23928 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 0 121728 800 121848 6 io_in[6]
port 64 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 io_in[7]
port 65 nsew signal input
rlabel metal2 s 135258 145428 135314 146228 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 143284 129208 144084 129328 6 io_in[9]
port 67 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 io_oeb[0]
port 68 nsew signal output
rlabel metal2 s 132958 0 133014 800 6 io_oeb[10]
port 69 nsew signal output
rlabel metal2 s 119158 0 119214 800 6 io_oeb[11]
port 70 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 io_oeb[12]
port 71 nsew signal output
rlabel metal2 s 47858 145428 47914 146228 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 143284 82968 144084 83088 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 126058 145428 126114 146228 6 io_oeb[15]
port 74 nsew signal output
rlabel metal3 s 143284 32648 144084 32768 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 132038 145428 132094 146228 6 io_oeb[18]
port 77 nsew signal output
rlabel metal3 s 143284 53728 144084 53848 6 io_oeb[19]
port 78 nsew signal output
rlabel metal2 s 105818 0 105874 800 6 io_oeb[1]
port 79 nsew signal output
rlabel metal3 s 143284 87728 144084 87848 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 12438 145428 12494 146228 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 2318 0 2374 800 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 125138 0 125194 800 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s 143284 24488 144084 24608 6 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s 0 137368 800 137488 6 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 io_oeb[26]
port 86 nsew signal output
rlabel metal2 s 65338 145428 65394 146228 6 io_oeb[27]
port 87 nsew signal output
rlabel metal2 s 29458 145428 29514 146228 6 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 io_oeb[29]
port 89 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s 0 110168 800 110288 6 io_oeb[30]
port 91 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 io_oeb[31]
port 92 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s 143284 20408 144084 20528 6 io_oeb[33]
port 94 nsew signal output
rlabel metal2 s 42338 145428 42394 146228 6 io_oeb[34]
port 95 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 io_oeb[36]
port 97 nsew signal output
rlabel metal2 s 19798 145428 19854 146228 6 io_oeb[37]
port 98 nsew signal output
rlabel metal2 s 143538 0 143594 800 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 io_oeb[4]
port 100 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 io_oeb[5]
port 101 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 io_oeb[6]
port 102 nsew signal output
rlabel metal2 s 31298 145428 31354 146228 6 io_oeb[7]
port 103 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 io_oeb[8]
port 104 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 io_oeb[9]
port 105 nsew signal output
rlabel metal2 s 66258 145428 66314 146228 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 io_out[10]
port 107 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 143284 88408 144084 88528 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 0 86368 800 86488 6 io_out[13]
port 110 nsew signal output
rlabel metal2 s 84198 0 84254 800 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 126518 145428 126574 146228 6 io_out[15]
port 112 nsew signal output
rlabel metal3 s 143284 138728 144084 138848 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 8298 145428 8354 146228 6 io_out[17]
port 114 nsew signal output
rlabel metal3 s 143284 21088 144084 21208 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 0 125808 800 125928 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 97078 145428 97134 146228 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 63958 145428 64014 146228 6 io_out[21]
port 119 nsew signal output
rlabel metal3 s 0 105408 800 105528 6 io_out[22]
port 120 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s 143284 124448 144084 124568 6 io_out[24]
port 122 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 io_out[25]
port 123 nsew signal output
rlabel metal2 s 61658 0 61714 800 6 io_out[26]
port 124 nsew signal output
rlabel metal2 s 131118 145428 131174 146228 6 io_out[27]
port 125 nsew signal output
rlabel metal2 s 123298 0 123354 800 6 io_out[28]
port 126 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 io_out[29]
port 127 nsew signal output
rlabel metal2 s 101218 0 101274 800 6 io_out[2]
port 128 nsew signal output
rlabel metal2 s 51078 145428 51134 146228 6 io_out[30]
port 129 nsew signal output
rlabel metal3 s 143284 86368 144084 86488 6 io_out[31]
port 130 nsew signal output
rlabel metal3 s 0 114928 800 115048 6 io_out[32]
port 131 nsew signal output
rlabel metal2 s 56138 145428 56194 146228 6 io_out[33]
port 132 nsew signal output
rlabel metal2 s 3238 145428 3294 146228 6 io_out[34]
port 133 nsew signal output
rlabel metal3 s 143284 65288 144084 65408 6 io_out[35]
port 134 nsew signal output
rlabel metal2 s 10138 145428 10194 146228 6 io_out[36]
port 135 nsew signal output
rlabel metal3 s 0 82288 800 82408 6 io_out[37]
port 136 nsew signal output
rlabel metal2 s 139398 145428 139454 146228 6 io_out[3]
port 137 nsew signal output
rlabel metal2 s 113178 145428 113234 146228 6 io_out[4]
port 138 nsew signal output
rlabel metal2 s 136638 145428 136694 146228 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 io_out[6]
port 140 nsew signal output
rlabel metal2 s 127438 145428 127494 146228 6 io_out[7]
port 141 nsew signal output
rlabel metal2 s 130658 0 130714 800 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 io_out[9]
port 143 nsew signal output
rlabel metal3 s 0 119008 800 119128 6 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 la_data_in[100]
port 145 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 la_data_in[101]
port 146 nsew signal input
rlabel metal3 s 143284 36728 144084 36848 6 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 106278 145428 106334 146228 6 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_data_in[104]
port 149 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 la_data_in[105]
port 150 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 la_data_in[106]
port 151 nsew signal input
rlabel metal3 s 143284 110848 144084 110968 6 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_data_in[109]
port 154 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 la_data_in[10]
port 155 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 la_data_in[110]
port 156 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 la_data_in[111]
port 157 nsew signal input
rlabel metal3 s 0 115608 800 115728 6 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 77298 145428 77354 146228 6 la_data_in[114]
port 160 nsew signal input
rlabel metal3 s 143284 33328 144084 33448 6 la_data_in[115]
port 161 nsew signal input
rlabel metal3 s 143284 91128 144084 91248 6 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 938 0 994 800 6 la_data_in[118]
port 164 nsew signal input
rlabel metal3 s 0 67328 800 67448 6 la_data_in[119]
port 165 nsew signal input
rlabel metal3 s 143284 57128 144084 57248 6 la_data_in[11]
port 166 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 114558 145428 114614 146228 6 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 44178 145428 44234 146228 6 la_data_in[124]
port 171 nsew signal input
rlabel metal3 s 143284 15648 144084 15768 6 la_data_in[125]
port 172 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 16118 145428 16174 146228 6 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 63038 145428 63094 146228 6 la_data_in[12]
port 175 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 la_data_in[13]
port 176 nsew signal input
rlabel metal3 s 143284 140088 144084 140208 6 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 la_data_in[15]
port 178 nsew signal input
rlabel metal3 s 0 118328 800 118448 6 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 938 145428 994 146228 6 la_data_in[17]
port 180 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 10598 145428 10654 146228 6 la_data_in[19]
port 182 nsew signal input
rlabel metal3 s 143284 60528 144084 60648 6 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 104898 145428 104954 146228 6 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 87878 145428 87934 146228 6 la_data_in[21]
port 185 nsew signal input
rlabel metal3 s 143284 63928 144084 64048 6 la_data_in[22]
port 186 nsew signal input
rlabel metal3 s 143284 132608 144084 132728 6 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 96158 145428 96214 146228 6 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 114098 0 114154 800 6 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 la_data_in[27]
port 191 nsew signal input
rlabel metal3 s 143284 27208 144084 27328 6 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 76838 145428 76894 146228 6 la_data_in[2]
port 194 nsew signal input
rlabel metal3 s 143284 48288 144084 48408 6 la_data_in[30]
port 195 nsew signal input
rlabel metal3 s 143284 13608 144084 13728 6 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 28078 145428 28134 146228 6 la_data_in[32]
port 197 nsew signal input
rlabel metal3 s 143284 133288 144084 133408 6 la_data_in[33]
port 198 nsew signal input
rlabel metal3 s 143284 53048 144084 53168 6 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 115938 145428 115994 146228 6 la_data_in[35]
port 200 nsew signal input
rlabel metal3 s 143284 29248 144084 29368 6 la_data_in[36]
port 201 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 la_data_in[37]
port 202 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 138938 145428 138994 146228 6 la_data_in[39]
port 204 nsew signal input
rlabel metal3 s 143284 36048 144084 36168 6 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 122378 145428 122434 146228 6 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 la_data_in[41]
port 207 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 45558 145428 45614 146228 6 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 102598 145428 102654 146228 6 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 72238 145428 72294 146228 6 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 34058 145428 34114 146228 6 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 24398 145428 24454 146228 6 la_data_in[47]
port 213 nsew signal input
rlabel metal3 s 143284 123088 144084 123208 6 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 5538 145428 5594 146228 6 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 la_data_in[4]
port 216 nsew signal input
rlabel metal3 s 143284 89768 144084 89888 6 la_data_in[50]
port 217 nsew signal input
rlabel metal3 s 0 130568 800 130688 6 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 66718 145428 66774 146228 6 la_data_in[52]
port 219 nsew signal input
rlabel metal3 s 143284 104048 144084 104168 6 la_data_in[53]
port 220 nsew signal input
rlabel metal3 s 143284 125808 144084 125928 6 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 48778 145428 48834 146228 6 la_data_in[55]
port 222 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 51538 145428 51594 146228 6 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 136178 0 136234 800 6 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 133418 145428 133474 146228 6 la_data_in[59]
port 226 nsew signal input
rlabel metal3 s 143284 51688 144084 51808 6 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 128358 145428 128414 146228 6 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 71318 145428 71374 146228 6 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 125138 145428 125194 146228 6 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 61658 145428 61714 146228 6 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 73618 145428 73674 146228 6 la_data_in[65]
port 233 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_data_in[67]
port 235 nsew signal input
rlabel metal3 s 143284 41488 144084 41608 6 la_data_in[68]
port 236 nsew signal input
rlabel metal3 s 143284 142128 144084 142248 6 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 la_data_in[6]
port 238 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 la_data_in[70]
port 239 nsew signal input
rlabel metal3 s 143284 116288 144084 116408 6 la_data_in[71]
port 240 nsew signal input
rlabel metal3 s 143284 127848 144084 127968 6 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 95698 145428 95754 146228 6 la_data_in[73]
port 242 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 la_data_in[74]
port 243 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 31758 145428 31814 146228 6 la_data_in[78]
port 247 nsew signal input
rlabel metal3 s 143284 74128 144084 74248 6 la_data_in[79]
port 248 nsew signal input
rlabel metal3 s 0 75488 800 75608 6 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 16578 145428 16634 146228 6 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 123758 145428 123814 146228 6 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 142618 145428 142674 146228 6 la_data_in[84]
port 254 nsew signal input
rlabel metal3 s 0 127848 800 127968 6 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 80518 145428 80574 146228 6 la_data_in[86]
port 256 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 23478 145428 23534 146228 6 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 78218 145428 78274 146228 6 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_data_in[8]
port 260 nsew signal input
rlabel metal3 s 143284 93168 144084 93288 6 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 108578 145428 108634 146228 6 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 52458 145428 52514 146228 6 la_data_in[93]
port 264 nsew signal input
rlabel metal3 s 0 134648 800 134768 6 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 103978 145428 104034 146228 6 la_data_in[98]
port 269 nsew signal input
rlabel metal3 s 143284 79568 144084 79688 6 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 121458 145428 121514 146228 6 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 la_data_out[100]
port 273 nsew signal output
rlabel metal3 s 0 61888 800 62008 6 la_data_out[101]
port 274 nsew signal output
rlabel metal3 s 143284 98608 144084 98728 6 la_data_out[102]
port 275 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 81898 145428 81954 146228 6 la_data_out[104]
port 277 nsew signal output
rlabel metal3 s 0 132608 800 132728 6 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 100298 0 100354 800 6 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 la_data_out[107]
port 280 nsew signal output
rlabel metal3 s 143284 1368 144084 1488 6 la_data_out[108]
port 281 nsew signal output
rlabel metal3 s 0 120368 800 120488 6 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 43258 145428 43314 146228 6 la_data_out[10]
port 283 nsew signal output
rlabel metal3 s 0 76848 800 76968 6 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 27158 145428 27214 146228 6 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 82818 0 82874 800 6 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 115478 145428 115534 146228 6 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 91098 145428 91154 146228 6 la_data_out[114]
port 288 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 la_data_out[115]
port 289 nsew signal output
rlabel metal3 s 0 80248 800 80368 6 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 38658 145428 38714 146228 6 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 34978 145428 35034 146228 6 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 143538 145428 143594 146228 6 la_data_out[119]
port 293 nsew signal output
rlabel metal3 s 143284 108808 144084 108928 6 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 la_data_out[120]
port 295 nsew signal output
rlabel metal3 s 0 138048 800 138168 6 la_data_out[121]
port 296 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 141238 145428 141294 146228 6 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 138478 0 138534 800 6 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 47858 0 47914 800 6 la_data_out[125]
port 300 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 la_data_out[126]
port 301 nsew signal output
rlabel metal3 s 0 133968 800 134088 6 la_data_out[127]
port 302 nsew signal output
rlabel metal3 s 143284 81608 144084 81728 6 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 127438 0 127494 800 6 la_data_out[13]
port 304 nsew signal output
rlabel metal3 s 143284 62568 144084 62688 6 la_data_out[14]
port 305 nsew signal output
rlabel metal3 s 0 101328 800 101448 6 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 139858 0 139914 800 6 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 49238 145428 49294 146228 6 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 72238 0 72294 800 6 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 60278 0 60334 800 6 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 107198 145428 107254 146228 6 la_data_out[21]
port 313 nsew signal output
rlabel metal3 s 143284 105408 144084 105528 6 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 57518 145428 57574 146228 6 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 53378 145428 53434 146228 6 la_data_out[24]
port 316 nsew signal output
rlabel metal3 s 143284 129888 144084 130008 6 la_data_out[25]
port 317 nsew signal output
rlabel metal3 s 143284 8848 144084 8968 6 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 103518 0 103574 800 6 la_data_out[27]
port 319 nsew signal output
rlabel metal3 s 143284 39448 144084 39568 6 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 la_data_out[2]
port 322 nsew signal output
rlabel metal3 s 143284 65968 144084 66088 6 la_data_out[30]
port 323 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 la_data_out[31]
port 324 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 28998 145428 29054 146228 6 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 la_data_out[34]
port 327 nsew signal output
rlabel metal3 s 143284 69368 144084 69488 6 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 138938 0 138994 800 6 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 120998 0 121054 800 6 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 138018 145428 138074 146228 6 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 55678 0 55734 800 6 la_data_out[39]
port 332 nsew signal output
rlabel metal3 s 0 122408 800 122528 6 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 95238 0 95294 800 6 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 la_data_out[41]
port 335 nsew signal output
rlabel metal3 s 143284 77528 144084 77648 6 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 116398 0 116454 800 6 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 la_data_out[45]
port 339 nsew signal output
rlabel metal3 s 143284 31288 144084 31408 6 la_data_out[46]
port 340 nsew signal output
rlabel metal3 s 143284 19048 144084 19168 6 la_data_out[47]
port 341 nsew signal output
rlabel metal3 s 143284 6808 144084 6928 6 la_data_out[48]
port 342 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 la_data_out[49]
port 343 nsew signal output
rlabel metal3 s 143284 84328 144084 84448 6 la_data_out[4]
port 344 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 101678 145428 101734 146228 6 la_data_out[51]
port 346 nsew signal output
rlabel metal3 s 143284 72768 144084 72888 6 la_data_out[52]
port 347 nsew signal output
rlabel metal3 s 143284 141448 144084 141568 6 la_data_out[53]
port 348 nsew signal output
rlabel metal3 s 143284 144848 144084 144968 6 la_data_out[54]
port 349 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 121458 0 121514 800 6 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 62118 145428 62174 146228 6 la_data_out[58]
port 353 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 124218 145428 124274 146228 6 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 124678 0 124734 800 6 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 la_data_out[61]
port 357 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 la_data_out[62]
port 358 nsew signal output
rlabel metal3 s 143284 40128 144084 40248 6 la_data_out[63]
port 359 nsew signal output
rlabel metal3 s 143284 50328 144084 50448 6 la_data_out[64]
port 360 nsew signal output
rlabel metal3 s 143284 22448 144084 22568 6 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 79598 145428 79654 146228 6 la_data_out[66]
port 362 nsew signal output
rlabel metal3 s 143284 27888 144084 28008 6 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 79138 145428 79194 146228 6 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 la_data_out[69]
port 365 nsew signal output
rlabel metal3 s 0 123768 800 123888 6 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 41878 145428 41934 146228 6 la_data_out[70]
port 367 nsew signal output
rlabel metal3 s 143284 131248 144084 131368 6 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 137098 145428 137154 146228 6 la_data_out[72]
port 369 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 la_data_out[73]
port 370 nsew signal output
rlabel metal3 s 0 97928 800 98048 6 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 73158 0 73214 800 6 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 la_data_out[77]
port 374 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 83278 145428 83334 146228 6 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 140318 145428 140374 146228 6 la_data_out[7]
port 377 nsew signal output
rlabel metal3 s 143284 96568 144084 96688 6 la_data_out[80]
port 378 nsew signal output
rlabel metal3 s 143284 25848 144084 25968 6 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 69018 145428 69074 146228 6 la_data_out[82]
port 380 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 118698 0 118754 800 6 la_data_out[85]
port 383 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 la_data_out[86]
port 384 nsew signal output
rlabel metal3 s 143284 55768 144084 55888 6 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 130658 145428 130714 146228 6 la_data_out[88]
port 386 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 100298 145428 100354 146228 6 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 23018 145428 23074 146228 6 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 20718 145428 20774 146228 6 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 99378 145428 99434 146228 6 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 111338 145428 111394 146228 6 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 la_data_out[94]
port 393 nsew signal output
rlabel metal3 s 143284 49648 144084 49768 6 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 46478 145428 46534 146228 6 la_data_out[96]
port 395 nsew signal output
rlabel metal3 s 0 78888 800 79008 6 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 la_data_out[98]
port 397 nsew signal output
rlabel metal3 s 143284 106768 144084 106888 6 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 76838 0 76894 800 6 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 la_oenb[100]
port 401 nsew signal input
rlabel metal3 s 143284 5448 144084 5568 6 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 35898 145428 35954 146228 6 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 la_oenb[104]
port 405 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 la_oenb[105]
port 406 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 la_oenb[106]
port 407 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 85118 145428 85174 146228 6 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 40958 145428 41014 146228 6 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 55218 145428 55274 146228 6 la_oenb[110]
port 412 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 la_oenb[111]
port 413 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 115478 0 115534 800 6 la_oenb[113]
port 415 nsew signal input
rlabel metal3 s 143284 136688 144084 136808 6 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 la_oenb[115]
port 417 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 44638 145428 44694 146228 6 la_oenb[117]
port 419 nsew signal input
rlabel metal3 s 143284 119008 144084 119128 6 la_oenb[118]
port 420 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 129738 145428 129794 146228 6 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 la_oenb[120]
port 423 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 la_oenb[121]
port 424 nsew signal input
rlabel metal3 s 143284 100648 144084 100768 6 la_oenb[122]
port 425 nsew signal input
rlabel metal3 s 143284 14288 144084 14408 6 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 5998 145428 6054 146228 6 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 la_oenb[127]
port 430 nsew signal input
rlabel metal3 s 143284 117648 144084 117768 6 la_oenb[12]
port 431 nsew signal input
rlabel metal3 s 143284 97248 144084 97368 6 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 117778 145428 117834 146228 6 la_oenb[14]
port 433 nsew signal input
rlabel metal3 s 143284 99968 144084 100088 6 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 17498 145428 17554 146228 6 la_oenb[17]
port 436 nsew signal input
rlabel metal3 s 143284 91808 144084 91928 6 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 126058 0 126114 800 6 la_oenb[19]
port 438 nsew signal input
rlabel metal3 s 0 143488 800 143608 6 la_oenb[1]
port 439 nsew signal input
rlabel metal3 s 143284 76168 144084 76288 6 la_oenb[20]
port 440 nsew signal input
rlabel metal3 s 0 124448 800 124568 6 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 74998 145428 75054 146228 6 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 53838 145428 53894 146228 6 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 112258 145428 112314 146228 6 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 12898 145428 12954 146228 6 la_oenb[27]
port 447 nsew signal input
rlabel metal3 s 143284 11568 144084 11688 6 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 la_oenb[29]
port 449 nsew signal input
rlabel metal3 s 143284 78208 144084 78328 6 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 la_oenb[31]
port 452 nsew signal input
rlabel metal3 s 143284 58488 144084 58608 6 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 74538 145428 74594 146228 6 la_oenb[33]
port 454 nsew signal input
rlabel metal3 s 143284 46248 144084 46368 6 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 142618 0 142674 800 6 la_oenb[37]
port 458 nsew signal input
rlabel metal3 s 143284 126488 144084 126608 6 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_oenb[39]
port 460 nsew signal input
rlabel metal3 s 0 113568 800 113688 6 la_oenb[3]
port 461 nsew signal input
rlabel metal3 s 0 99968 800 100088 6 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 89718 145428 89774 146228 6 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 la_oenb[42]
port 464 nsew signal input
rlabel metal3 s 143284 61888 144084 62008 6 la_oenb[43]
port 465 nsew signal input
rlabel metal3 s 0 129208 800 129328 6 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_oenb[45]
port 467 nsew signal input
rlabel metal3 s 143284 55088 144084 55208 6 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 135718 145428 135774 146228 6 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 58438 145428 58494 146228 6 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 478 0 534 800 6 la_oenb[4]
port 472 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 1398 145428 1454 146228 6 la_oenb[51]
port 474 nsew signal input
rlabel metal3 s 143284 30608 144084 30728 6 la_oenb[52]
port 475 nsew signal input
rlabel metal3 s 143284 70728 144084 70848 6 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_oenb[54]
port 477 nsew signal input
rlabel metal3 s 0 108808 800 108928 6 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 33598 145428 33654 146228 6 la_oenb[56]
port 479 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 75918 145428 75974 146228 6 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 97998 145428 98054 146228 6 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 la_oenb[60]
port 484 nsew signal input
rlabel metal3 s 143284 44888 144084 45008 6 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 la_oenb[62]
port 486 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 la_oenb[63]
port 487 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 la_oenb[64]
port 488 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 9218 145428 9274 146228 6 la_oenb[66]
port 490 nsew signal input
rlabel metal3 s 143284 17688 144084 17808 6 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 82818 145428 82874 146228 6 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 112258 0 112314 800 6 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 103058 145428 103114 146228 6 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 40038 145428 40094 146228 6 la_oenb[71]
port 496 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 64418 145428 64474 146228 6 la_oenb[74]
port 499 nsew signal input
rlabel metal3 s 0 136008 800 136128 6 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 15198 145428 15254 146228 6 la_oenb[76]
port 501 nsew signal input
rlabel metal3 s 143284 4768 144084 4888 6 la_oenb[77]
port 502 nsew signal input
rlabel metal3 s 0 142808 800 142928 6 la_oenb[78]
port 503 nsew signal input
rlabel metal3 s 143284 34688 144084 34808 6 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_oenb[7]
port 505 nsew signal input
rlabel metal3 s 143284 121048 144084 121168 6 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 109038 145428 109094 146228 6 la_oenb[81]
port 507 nsew signal input
rlabel metal3 s 0 95888 800 96008 6 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 la_oenb[83]
port 509 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 la_oenb[84]
port 510 nsew signal input
rlabel metal3 s 143284 67328 144084 67448 6 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 122838 145428 122894 146228 6 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 60738 145428 60794 146228 6 la_oenb[87]
port 513 nsew signal input
rlabel metal3 s 143284 138048 144084 138168 6 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_oenb[89]
port 515 nsew signal input
rlabel metal3 s 143284 110168 144084 110288 6 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 92478 145428 92534 146228 6 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 141698 145428 141754 146228 6 la_oenb[93]
port 520 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 la_oenb[94]
port 521 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_oenb[96]
port 523 nsew signal input
rlabel metal3 s 143284 119688 144084 119808 6 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 72698 145428 72754 146228 6 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 120538 145428 120594 146228 6 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 user_clock2
port 528 nsew signal input
rlabel metal2 s 21178 145428 21234 146228 6 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 105358 145428 105414 146228 6 user_irq[2]
port 531 nsew signal output
rlabel metal2 s 69938 145428 69994 146228 6 wb_clk_i
port 532 nsew signal input
rlabel metal3 s 143284 3408 144084 3528 6 wb_rst_i
port 533 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 wbs_ack_o
port 534 nsew signal output
rlabel metal2 s 68098 145428 68154 146228 6 wbs_adr_i[0]
port 535 nsew signal input
rlabel metal3 s 143284 42848 144084 42968 6 wbs_adr_i[10]
port 536 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 wbs_adr_i[11]
port 537 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 wbs_adr_i[12]
port 538 nsew signal input
rlabel metal3 s 0 141448 800 141568 6 wbs_adr_i[13]
port 539 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 wbs_adr_i[14]
port 540 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 wbs_adr_i[15]
port 541 nsew signal input
rlabel metal3 s 143284 113568 144084 113688 6 wbs_adr_i[16]
port 542 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 wbs_adr_i[17]
port 543 nsew signal input
rlabel metal3 s 143284 10208 144084 10328 6 wbs_adr_i[18]
port 544 nsew signal input
rlabel metal2 s 86498 145428 86554 146228 6 wbs_adr_i[19]
port 545 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_adr_i[1]
port 546 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 wbs_adr_i[20]
port 547 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_adr_i[21]
port 548 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 wbs_adr_i[22]
port 549 nsew signal input
rlabel metal2 s 59358 145428 59414 146228 6 wbs_adr_i[23]
port 550 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wbs_adr_i[24]
port 551 nsew signal input
rlabel metal2 s 133878 0 133934 800 6 wbs_adr_i[25]
port 552 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 wbs_adr_i[26]
port 553 nsew signal input
rlabel metal2 s 93398 145428 93454 146228 6 wbs_adr_i[27]
port 554 nsew signal input
rlabel metal2 s 7838 145428 7894 146228 6 wbs_adr_i[28]
port 555 nsew signal input
rlabel metal3 s 143284 143488 144084 143608 6 wbs_adr_i[29]
port 556 nsew signal input
rlabel metal2 s 18418 145428 18474 146228 6 wbs_adr_i[2]
port 557 nsew signal input
rlabel metal2 s 57058 145428 57114 146228 6 wbs_adr_i[30]
port 558 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_adr_i[31]
port 559 nsew signal input
rlabel metal3 s 143284 80928 144084 81048 6 wbs_adr_i[3]
port 560 nsew signal input
rlabel metal2 s 30378 145428 30434 146228 6 wbs_adr_i[4]
port 561 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 wbs_adr_i[5]
port 562 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 wbs_adr_i[6]
port 563 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 wbs_adr_i[7]
port 564 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 wbs_adr_i[8]
port 565 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 wbs_adr_i[9]
port 566 nsew signal input
rlabel metal2 s 70398 145428 70454 146228 6 wbs_cyc_i
port 567 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 wbs_dat_i[0]
port 568 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 wbs_dat_i[10]
port 569 nsew signal input
rlabel metal3 s 0 103368 800 103488 6 wbs_dat_i[11]
port 570 nsew signal input
rlabel metal2 s 118238 145428 118294 146228 6 wbs_dat_i[12]
port 571 nsew signal input
rlabel metal3 s 143284 122408 144084 122528 6 wbs_dat_i[13]
port 572 nsew signal input
rlabel metal3 s 143284 43528 144084 43648 6 wbs_dat_i[14]
port 573 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wbs_dat_i[15]
port 574 nsew signal input
rlabel metal3 s 0 56448 800 56568 6 wbs_dat_i[16]
port 575 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 wbs_dat_i[17]
port 576 nsew signal input
rlabel metal3 s 0 108128 800 108248 6 wbs_dat_i[18]
port 577 nsew signal input
rlabel metal2 s 98458 145428 98514 146228 6 wbs_dat_i[19]
port 578 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 wbs_dat_i[1]
port 579 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 wbs_dat_i[20]
port 580 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_i[21]
port 581 nsew signal input
rlabel metal2 s 132958 145428 133014 146228 6 wbs_dat_i[22]
port 582 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 wbs_dat_i[23]
port 583 nsew signal input
rlabel metal2 s 14278 145428 14334 146228 6 wbs_dat_i[24]
port 584 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 wbs_dat_i[25]
port 585 nsew signal input
rlabel metal3 s 143284 17008 144084 17128 6 wbs_dat_i[26]
port 586 nsew signal input
rlabel metal3 s 143284 46928 144084 47048 6 wbs_dat_i[27]
port 587 nsew signal input
rlabel metal2 s 46938 145428 46994 146228 6 wbs_dat_i[28]
port 588 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 wbs_dat_i[29]
port 589 nsew signal input
rlabel metal3 s 143284 135328 144084 135448 6 wbs_dat_i[2]
port 590 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wbs_dat_i[30]
port 591 nsew signal input
rlabel metal2 s 36358 145428 36414 146228 6 wbs_dat_i[31]
port 592 nsew signal input
rlabel metal2 s 94318 145428 94374 146228 6 wbs_dat_i[3]
port 593 nsew signal input
rlabel metal3 s 0 127168 800 127288 6 wbs_dat_i[4]
port 594 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_dat_i[5]
port 595 nsew signal input
rlabel metal2 s 113638 145428 113694 146228 6 wbs_dat_i[6]
port 596 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 wbs_dat_i[7]
port 597 nsew signal input
rlabel metal2 s 90178 145428 90234 146228 6 wbs_dat_i[8]
port 598 nsew signal input
rlabel metal3 s 0 131248 800 131368 6 wbs_dat_i[9]
port 599 nsew signal input
rlabel metal2 s 4618 145428 4674 146228 6 wbs_dat_o[0]
port 600 nsew signal output
rlabel metal3 s 143284 115608 144084 115728 6 wbs_dat_o[10]
port 601 nsew signal output
rlabel metal2 s 92938 0 92994 800 6 wbs_dat_o[11]
port 602 nsew signal output
rlabel metal2 s 134338 0 134394 800 6 wbs_dat_o[12]
port 603 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_o[13]
port 604 nsew signal output
rlabel metal3 s 0 106768 800 106888 6 wbs_dat_o[14]
port 605 nsew signal output
rlabel metal2 s 136638 0 136694 800 6 wbs_dat_o[15]
port 606 nsew signal output
rlabel metal2 s 110878 145428 110934 146228 6 wbs_dat_o[16]
port 607 nsew signal output
rlabel metal2 s 2318 145428 2374 146228 6 wbs_dat_o[17]
port 608 nsew signal output
rlabel metal3 s 143284 72088 144084 72208 6 wbs_dat_o[18]
port 609 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 wbs_dat_o[19]
port 610 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 wbs_dat_o[1]
port 611 nsew signal output
rlabel metal2 s 59818 145428 59874 146228 6 wbs_dat_o[20]
port 612 nsew signal output
rlabel metal2 s 32678 145428 32734 146228 6 wbs_dat_o[21]
port 613 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 wbs_dat_o[22]
port 614 nsew signal output
rlabel metal2 s 6918 145428 6974 146228 6 wbs_dat_o[23]
port 615 nsew signal output
rlabel metal2 s 92018 145428 92074 146228 6 wbs_dat_o[24]
port 616 nsew signal output
rlabel metal3 s 143284 95208 144084 95328 6 wbs_dat_o[25]
port 617 nsew signal output
rlabel metal2 s 100758 145428 100814 146228 6 wbs_dat_o[26]
port 618 nsew signal output
rlabel metal2 s 119158 145428 119214 146228 6 wbs_dat_o[27]
port 619 nsew signal output
rlabel metal3 s 143284 38088 144084 38208 6 wbs_dat_o[28]
port 620 nsew signal output
rlabel metal2 s 22098 145428 22154 146228 6 wbs_dat_o[29]
port 621 nsew signal output
rlabel metal3 s 0 89088 800 89208 6 wbs_dat_o[2]
port 622 nsew signal output
rlabel metal2 s 109958 145428 110014 146228 6 wbs_dat_o[30]
port 623 nsew signal output
rlabel metal2 s 39578 145428 39634 146228 6 wbs_dat_o[31]
port 624 nsew signal output
rlabel metal3 s 0 89768 800 89888 6 wbs_dat_o[3]
port 625 nsew signal output
rlabel metal2 s 25318 145428 25374 146228 6 wbs_dat_o[4]
port 626 nsew signal output
rlabel metal2 s 85578 145428 85634 146228 6 wbs_dat_o[5]
port 627 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 wbs_dat_o[6]
port 628 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_o[7]
port 629 nsew signal output
rlabel metal3 s 143284 102008 144084 102128 6 wbs_dat_o[8]
port 630 nsew signal output
rlabel metal3 s 143284 103368 144084 103488 6 wbs_dat_o[9]
port 631 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 wbs_sel_i[0]
port 632 nsew signal input
rlabel metal2 s 13818 145428 13874 146228 6 wbs_sel_i[1]
port 633 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 wbs_sel_i[2]
port 634 nsew signal input
rlabel metal2 s 26698 145428 26754 146228 6 wbs_sel_i[3]
port 635 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 wbs_stb_i
port 636 nsew signal input
rlabel metal2 s 81438 145428 81494 146228 6 wbs_we_i
port 637 nsew signal input
rlabel metal4 s 108804 -1864 109404 147656 6 vccd1
port 638 nsew power bidirectional
rlabel metal4 s 72804 -1864 73404 147656 6 vccd1
port 639 nsew power bidirectional
rlabel metal4 s 36804 -1864 37404 147656 6 vccd1
port 640 nsew power bidirectional
rlabel metal4 s 804 -1864 1404 147656 6 vccd1
port 641 nsew power bidirectional
rlabel metal4 s 145468 -924 146068 146716 6 vccd1
port 642 nsew power bidirectional
rlabel metal4 s -1996 -924 -1396 146716 4 vccd1
port 643 nsew power bidirectional
rlabel metal5 s -1996 146116 146068 146716 6 vccd1
port 644 nsew power bidirectional
rlabel metal5 s -2936 109828 147008 110428 6 vccd1
port 645 nsew power bidirectional
rlabel metal5 s -2936 73828 147008 74428 6 vccd1
port 646 nsew power bidirectional
rlabel metal5 s -2936 37828 147008 38428 6 vccd1
port 647 nsew power bidirectional
rlabel metal5 s -2936 1828 147008 2428 6 vccd1
port 648 nsew power bidirectional
rlabel metal5 s -1996 -924 146068 -324 8 vccd1
port 649 nsew power bidirectional
rlabel metal4 s 146408 -1864 147008 147656 6 vssd1
port 650 nsew ground bidirectional
rlabel metal4 s 126804 -1864 127404 147656 6 vssd1
port 651 nsew ground bidirectional
rlabel metal4 s 90804 -1864 91404 147656 6 vssd1
port 652 nsew ground bidirectional
rlabel metal4 s 54804 -1864 55404 147656 6 vssd1
port 653 nsew ground bidirectional
rlabel metal4 s 18804 -1864 19404 147656 6 vssd1
port 654 nsew ground bidirectional
rlabel metal4 s -2936 -1864 -2336 147656 4 vssd1
port 655 nsew ground bidirectional
rlabel metal5 s -2936 147056 147008 147656 6 vssd1
port 656 nsew ground bidirectional
rlabel metal5 s -2936 127828 147008 128428 6 vssd1
port 657 nsew ground bidirectional
rlabel metal5 s -2936 91828 147008 92428 6 vssd1
port 658 nsew ground bidirectional
rlabel metal5 s -2936 55828 147008 56428 6 vssd1
port 659 nsew ground bidirectional
rlabel metal5 s -2936 19828 147008 20428 6 vssd1
port 660 nsew ground bidirectional
rlabel metal5 s -2936 -1864 147008 -1264 8 vssd1
port 661 nsew ground bidirectional
rlabel metal4 s 112404 -3744 113004 149536 6 vccd2
port 662 nsew power bidirectional
rlabel metal4 s 76404 -3744 77004 149536 6 vccd2
port 663 nsew power bidirectional
rlabel metal4 s 40404 -3744 41004 149536 6 vccd2
port 664 nsew power bidirectional
rlabel metal4 s 4404 -3744 5004 149536 6 vccd2
port 665 nsew power bidirectional
rlabel metal4 s 147348 -2804 147948 148596 6 vccd2
port 666 nsew power bidirectional
rlabel metal4 s -3876 -2804 -3276 148596 4 vccd2
port 667 nsew power bidirectional
rlabel metal5 s -3876 147996 147948 148596 6 vccd2
port 668 nsew power bidirectional
rlabel metal5 s -4816 113476 148888 114076 6 vccd2
port 669 nsew power bidirectional
rlabel metal5 s -4816 77476 148888 78076 6 vccd2
port 670 nsew power bidirectional
rlabel metal5 s -4816 41476 148888 42076 6 vccd2
port 671 nsew power bidirectional
rlabel metal5 s -4816 5476 148888 6076 6 vccd2
port 672 nsew power bidirectional
rlabel metal5 s -3876 -2804 147948 -2204 8 vccd2
port 673 nsew power bidirectional
rlabel metal4 s 148288 -3744 148888 149536 6 vssd2
port 674 nsew ground bidirectional
rlabel metal4 s 130404 -3744 131004 149536 6 vssd2
port 675 nsew ground bidirectional
rlabel metal4 s 94404 -3744 95004 149536 6 vssd2
port 676 nsew ground bidirectional
rlabel metal4 s 58404 -3744 59004 149536 6 vssd2
port 677 nsew ground bidirectional
rlabel metal4 s 22404 -3744 23004 149536 6 vssd2
port 678 nsew ground bidirectional
rlabel metal4 s -4816 -3744 -4216 149536 4 vssd2
port 679 nsew ground bidirectional
rlabel metal5 s -4816 148936 148888 149536 6 vssd2
port 680 nsew ground bidirectional
rlabel metal5 s -4816 131476 148888 132076 6 vssd2
port 681 nsew ground bidirectional
rlabel metal5 s -4816 95476 148888 96076 6 vssd2
port 682 nsew ground bidirectional
rlabel metal5 s -4816 59476 148888 60076 6 vssd2
port 683 nsew ground bidirectional
rlabel metal5 s -4816 23476 148888 24076 6 vssd2
port 684 nsew ground bidirectional
rlabel metal5 s -4816 -3744 148888 -3144 8 vssd2
port 685 nsew ground bidirectional
rlabel metal4 s 116004 -5624 116604 151416 6 vdda1
port 686 nsew power bidirectional
rlabel metal4 s 80004 -5624 80604 151416 6 vdda1
port 687 nsew power bidirectional
rlabel metal4 s 44004 -5624 44604 151416 6 vdda1
port 688 nsew power bidirectional
rlabel metal4 s 8004 -5624 8604 151416 6 vdda1
port 689 nsew power bidirectional
rlabel metal4 s 149228 -4684 149828 150476 6 vdda1
port 690 nsew power bidirectional
rlabel metal4 s -5756 -4684 -5156 150476 4 vdda1
port 691 nsew power bidirectional
rlabel metal5 s -5756 149876 149828 150476 6 vdda1
port 692 nsew power bidirectional
rlabel metal5 s -6696 117076 150768 117676 6 vdda1
port 693 nsew power bidirectional
rlabel metal5 s -6696 81076 150768 81676 6 vdda1
port 694 nsew power bidirectional
rlabel metal5 s -6696 45076 150768 45676 6 vdda1
port 695 nsew power bidirectional
rlabel metal5 s -6696 9076 150768 9676 6 vdda1
port 696 nsew power bidirectional
rlabel metal5 s -5756 -4684 149828 -4084 8 vdda1
port 697 nsew power bidirectional
rlabel metal4 s 150168 -5624 150768 151416 6 vssa1
port 698 nsew ground bidirectional
rlabel metal4 s 134004 -5624 134604 151416 6 vssa1
port 699 nsew ground bidirectional
rlabel metal4 s 98004 -5624 98604 151416 6 vssa1
port 700 nsew ground bidirectional
rlabel metal4 s 62004 -5624 62604 151416 6 vssa1
port 701 nsew ground bidirectional
rlabel metal4 s 26004 -5624 26604 151416 6 vssa1
port 702 nsew ground bidirectional
rlabel metal4 s -6696 -5624 -6096 151416 4 vssa1
port 703 nsew ground bidirectional
rlabel metal5 s -6696 150816 150768 151416 6 vssa1
port 704 nsew ground bidirectional
rlabel metal5 s -6696 135076 150768 135676 6 vssa1
port 705 nsew ground bidirectional
rlabel metal5 s -6696 99076 150768 99676 6 vssa1
port 706 nsew ground bidirectional
rlabel metal5 s -6696 63076 150768 63676 6 vssa1
port 707 nsew ground bidirectional
rlabel metal5 s -6696 27076 150768 27676 6 vssa1
port 708 nsew ground bidirectional
rlabel metal5 s -6696 -5624 150768 -5024 8 vssa1
port 709 nsew ground bidirectional
rlabel metal4 s 119604 -7504 120204 153296 6 vdda2
port 710 nsew power bidirectional
rlabel metal4 s 83604 -7504 84204 153296 6 vdda2
port 711 nsew power bidirectional
rlabel metal4 s 47604 -7504 48204 153296 6 vdda2
port 712 nsew power bidirectional
rlabel metal4 s 11604 -7504 12204 153296 6 vdda2
port 713 nsew power bidirectional
rlabel metal4 s 151108 -6564 151708 152356 6 vdda2
port 714 nsew power bidirectional
rlabel metal4 s -7636 -6564 -7036 152356 4 vdda2
port 715 nsew power bidirectional
rlabel metal5 s -7636 151756 151708 152356 6 vdda2
port 716 nsew power bidirectional
rlabel metal5 s -8576 120676 152648 121276 6 vdda2
port 717 nsew power bidirectional
rlabel metal5 s -8576 84676 152648 85276 6 vdda2
port 718 nsew power bidirectional
rlabel metal5 s -8576 48676 152648 49276 6 vdda2
port 719 nsew power bidirectional
rlabel metal5 s -8576 12676 152648 13276 6 vdda2
port 720 nsew power bidirectional
rlabel metal5 s -7636 -6564 151708 -5964 8 vdda2
port 721 nsew power bidirectional
rlabel metal4 s 152048 -7504 152648 153296 6 vssa2
port 722 nsew ground bidirectional
rlabel metal4 s 137604 -7504 138204 153296 6 vssa2
port 723 nsew ground bidirectional
rlabel metal4 s 101604 -7504 102204 153296 6 vssa2
port 724 nsew ground bidirectional
rlabel metal4 s 65604 -7504 66204 153296 6 vssa2
port 725 nsew ground bidirectional
rlabel metal4 s 29604 -7504 30204 153296 6 vssa2
port 726 nsew ground bidirectional
rlabel metal4 s -8576 -7504 -7976 153296 4 vssa2
port 727 nsew ground bidirectional
rlabel metal5 s -8576 152696 152648 153296 6 vssa2
port 728 nsew ground bidirectional
rlabel metal5 s -8576 138676 152648 139276 6 vssa2
port 729 nsew ground bidirectional
rlabel metal5 s -8576 102676 152648 103276 6 vssa2
port 730 nsew ground bidirectional
rlabel metal5 s -8576 66676 152648 67276 6 vssa2
port 731 nsew ground bidirectional
rlabel metal5 s -8576 30676 152648 31276 6 vssa2
port 732 nsew ground bidirectional
rlabel metal5 s -8576 -7504 152648 -6904 8 vssa2
port 733 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 144084 146228
string LEFview TRUE
string GDS_FILE /project/openlane/user_project_wrapper/runs/user_project_wrapper/results/magic/user_project_wrapper.gds
string GDS_END 45072358
string GDS_START 130
<< end >>

