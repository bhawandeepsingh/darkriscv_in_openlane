VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 902.775 BY 913.495 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 909.495 23.370 913.495 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 703.840 902.775 704.440 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 0.000 699.570 4.000 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.840 4.000 874.440 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 717.440 902.775 718.040 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 0.000 805.370 4.000 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 0.000 614.470 4.000 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 909.495 547.770 913.495 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.490 0.000 846.770 4.000 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 0.000 533.970 4.000 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 370.640 902.775 371.240 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 909.495 593.770 913.495 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 0.000 552.370 4.000 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 909.495 674.270 913.495 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 591.640 902.775 592.240 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 843.240 902.775 843.840 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 4.000 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 880.640 4.000 881.240 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 0.000 428.170 4.000 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 909.495 731.770 913.495 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 469.240 902.775 469.840 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 0.000 814.570 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.890 909.495 842.170 913.495 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 909.495 313.170 913.495 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 909.495 161.370 913.495 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 0.000 717.970 4.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 533.840 902.775 534.440 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.390 909.495 807.670 913.495 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 13.640 902.775 14.240 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 0.000 324.670 4.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 0.000 510.970 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.790 909.495 527.070 913.495 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 909.495 556.970 913.495 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 909.495 343.070 913.495 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 428.440 902.775 429.040 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 909.495 232.670 913.495 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 909.495 237.270 913.495 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 909.495 750.170 913.495 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 78.240 902.775 78.840 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 47.640 902.775 48.240 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 909.495 71.670 913.495 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.840 4.000 908.440 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 673.240 902.775 673.840 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.990 0.000 881.270 4.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 909.495 423.570 913.495 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 909.495 119.970 913.495 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.390 0.000 600.670 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 146.240 902.775 146.840 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.990 0.000 490.270 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.490 909.495 846.770 913.495 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 809.240 902.775 809.840 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 0.000 538.570 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.690 0.000 832.970 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.590 0.000 747.870 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 909.495 299.370 913.495 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 520.240 902.775 520.840 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 909.495 789.270 913.495 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 204.040 902.775 204.640 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.790 909.495 826.070 913.495 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 336.640 902.775 337.240 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 0.000 662.770 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 547.440 902.775 548.040 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 909.495 76.270 913.495 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 0.000 784.670 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 153.040 902.775 153.640 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.240 4.000 860.840 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 909.495 409.770 913.495 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 909.495 186.670 913.495 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.240 4.000 690.840 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 125.840 902.775 126.440 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 909.495 267.170 913.495 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 909.495 124.570 913.495 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.390 0.000 899.670 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.190 0.000 775.470 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 909.495 195.870 913.495 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 0.000 566.170 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 909.495 414.370 913.495 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 0.000 448.870 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 554.240 902.775 554.840 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 0.000 529.370 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 909.495 793.870 913.495 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 870.440 902.775 871.040 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 909.495 53.270 913.495 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 132.640 902.775 133.240 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 0.000 439.670 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.290 909.495 607.570 913.495 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 909.495 400.570 913.495 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 778.640 902.775 779.240 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 909.495 821.470 913.495 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.590 0.000 770.870 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 0.000 543.170 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.590 0.000 632.870 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 909.495 317.770 913.495 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 540.640 902.775 541.240 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 909.495 352.270 913.495 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 909.495 18.770 913.495 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 408.040 902.775 408.640 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 909.495 62.470 913.495 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.090 909.495 874.370 913.495 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 909.495 708.770 913.495 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 909.495 855.970 913.495 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 909.495 798.470 913.495 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.890 0.000 819.170 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 744.640 4.000 745.240 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 0.000 809.970 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 231.240 902.775 231.840 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.790 909.495 665.070 913.495 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 693.640 902.775 694.240 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.240 4.000 724.840 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.490 0.000 823.770 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 909.495 485.670 913.495 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 210.840 902.775 211.440 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 567.840 902.775 568.440 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 357.040 902.775 357.640 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 0.000 205.070 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 909.495 717.970 913.495 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 909.495 276.370 913.495 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 98.640 902.775 99.240 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 909.495 99.270 913.495 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 909.495 393.670 913.495 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 877.240 902.775 877.840 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 909.495 4.970 913.495 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 909.495 67.070 913.495 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 380.840 902.775 381.440 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.590 909.495 655.870 913.495 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 909.495 552.370 913.495 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 401.240 902.775 401.840 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 829.640 902.775 830.240 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 0.000 382.170 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 909.495 602.970 913.495 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 0.000 713.370 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 0.000 343.070 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 170.040 902.775 170.640 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 909.495 481.070 913.495 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 302.640 902.775 303.240 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 85.040 902.775 85.640 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 909.495 175.170 913.495 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 836.440 902.775 837.040 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 329.840 902.775 330.440 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.890 909.495 727.170 913.495 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 183.640 902.775 184.240 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 909.495 869.770 913.495 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 224.440 902.775 225.040 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 909.495 766.270 913.495 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 909.495 285.570 913.495 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 909.495 642.070 913.495 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 909.495 451.170 913.495 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 909.495 214.270 913.495 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 909.495 152.170 913.495 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 771.840 902.775 772.440 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 909.495 32.570 913.495 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 561.040 902.775 561.640 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 816.040 4.000 816.640 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 909.495 418.970 913.495 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 652.840 902.775 653.440 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 785.440 902.775 786.040 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 909.495 303.970 913.495 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 909.495 322.370 913.495 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.090 0.000 851.370 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 909.495 837.570 913.495 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 323.040 902.775 323.640 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.790 909.495 803.070 913.495 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 909.495 446.570 913.495 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 909.495 784.670 913.495 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 0.000 504.070 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 909.495 384.470 913.495 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 909.495 460.370 913.495 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 0.000 561.570 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 258.440 902.775 259.040 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 890.840 902.775 891.440 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 731.040 902.775 731.640 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 799.040 902.775 799.640 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 909.495 598.370 913.495 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 0.000 586.870 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 909.495 200.470 913.495 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 462.440 902.775 463.040 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 909.495 103.870 913.495 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.190 909.495 775.470 913.495 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.490 909.495 892.770 913.495 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 4.000 803.040 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 909.495 504.070 913.495 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 909.495 147.570 913.495 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.990 909.495 490.270 913.495 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.690 0.000 694.970 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 581.440 902.775 582.040 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.590 909.495 678.870 913.495 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 909.495 329.270 913.495 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.390 0.000 738.670 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.190 0.000 890.470 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.990 909.495 651.270 913.495 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 499.840 902.775 500.440 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.390 909.495 761.670 913.495 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 0.000 690.370 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 618.840 902.775 619.440 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 909.495 513.270 913.495 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 6.840 902.775 7.440 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 909.495 271.770 913.495 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 909.495 170.570 913.495 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 0.000 520.170 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.290 909.495 722.570 913.495 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 909.495 570.770 913.495 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.840 4.000 500.440 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 909.495 241.870 913.495 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 909.495 218.870 913.495 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.090 909.495 897.370 913.495 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 680.040 902.775 680.640 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 909.495 883.570 913.495 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.190 0.000 867.470 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 513.440 902.775 514.040 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 0.000 800.770 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 394.440 902.775 395.040 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.390 0.000 876.670 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 909.495 308.570 913.495 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 0.000 453.470 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 0.000 377.570 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.390 0.000 623.670 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.390 909.495 669.670 913.495 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 659.640 902.775 660.240 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 909.495 361.470 913.495 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 909.495 333.870 913.495 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 816.040 902.775 816.640 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 54.440 902.775 55.040 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 0.000 646.670 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 244.840 902.775 245.440 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 0.000 315.470 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 414.840 902.775 415.440 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 909.495 182.070 913.495 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 435.240 902.775 435.840 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.790 0.000 872.070 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 0.000 757.070 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.890 909.495 865.170 913.495 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 486.240 902.775 486.840 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.190 0.000 729.470 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 0.000 828.370 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 197.240 902.775 197.840 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 119.040 902.775 119.640 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 40.840 902.775 41.440 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 527.040 902.775 527.640 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 909.495 637.470 913.495 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 455.640 902.775 456.240 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 884.040 902.775 884.640 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 904.440 902.775 905.040 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.390 0.000 761.670 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 909.495 389.070 913.495 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.790 909.495 780.070 913.495 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.790 0.000 780.070 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 251.640 902.775 252.240 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 316.240 902.775 316.840 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 139.440 902.775 140.040 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 909.495 499.470 913.495 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 176.840 902.775 177.440 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.590 909.495 494.870 913.495 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.240 4.000 775.840 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 909.495 262.570 913.495 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 822.840 902.775 823.440 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.290 909.495 860.570 913.495 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 909.495 522.470 913.495 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.690 909.495 878.970 913.495 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 605.240 902.775 605.840 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 159.840 902.775 160.440 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 909.495 432.770 913.495 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.990 0.000 743.270 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 350.240 902.775 350.840 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.590 909.495 816.870 913.495 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 909.495 628.270 913.495 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 909.495 142.970 913.495 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 909.495 129.170 913.495 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.390 909.495 623.670 913.495 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 909.495 699.570 913.495 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 309.440 902.775 310.040 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 909.495 290.170 913.495 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 666.440 902.775 667.040 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 0.000 481.070 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 34.040 902.775 34.640 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 909.495 223.470 913.495 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 909.495 531.670 913.495 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 0.000 642.070 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 909.495 257.970 913.495 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 909.495 347.670 913.495 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 856.840 902.775 857.440 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 909.495 280.970 913.495 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 744.640 902.775 745.240 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.990 909.495 812.270 913.495 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.190 0.000 752.470 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 632.440 902.775 633.040 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 91.840 902.775 92.440 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 0.000 524.770 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.290 0.000 860.570 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 909.495 39.470 913.495 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 737.840 902.775 738.440 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 612.040 902.775 612.640 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.090 909.495 736.370 913.495 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 625.640 902.775 626.240 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 0.000 356.870 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 909.495 110.770 913.495 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 574.640 902.775 575.240 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 0.000 789.270 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 901.040 4.000 901.640 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 476.040 902.775 476.640 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 909.495 471.870 913.495 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 909.495 338.470 913.495 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 909.495 704.170 913.495 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 909.495 80.870 913.495 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 71.440 902.775 72.040 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 0.000 671.970 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 493.040 902.775 493.640 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 363.840 902.775 364.440 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 909.495 464.970 913.495 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 289.040 902.775 289.640 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.790 0.000 895.070 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 792.240 902.775 792.840 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 710.640 4.000 711.240 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 909.495 561.570 913.495 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 387.640 902.775 388.240 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.240 4.000 809.840 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.790 0.000 734.070 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 343.440 902.775 344.040 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.090 909.495 851.370 913.495 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 909.495 366.070 913.495 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 909.495 9.570 913.495 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 190.440 902.775 191.040 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 442.040 902.775 442.640 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 0.000 476.470 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 909.495 209.670 913.495 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 0.000 766.270 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 909.495 476.470 913.495 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 909.495 614.470 913.495 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 0.000 619.070 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 282.240 902.775 282.840 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 909.495 57.870 913.495 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 112.240 902.775 112.840 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 0.000 462.670 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 909.495 517.870 913.495 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 0.000 704.170 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 909.495 646.670 913.495 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 909.495 251.070 913.495 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 0.000 676.570 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 909.495 405.170 913.495 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.040 4.000 850.640 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 909.495 94.670 913.495 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 27.240 902.775 27.840 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.240 4.000 894.840 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 217.640 902.775 218.240 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 758.240 902.775 758.840 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 909.495 683.470 913.495 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.890 0.000 681.170 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 421.640 902.775 422.240 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.590 909.495 770.870 913.495 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 909.495 379.870 913.495 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 863.640 902.775 864.240 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 686.840 902.775 687.440 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 0.000 414.370 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 909.495 579.970 913.495 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.890 909.495 888.170 913.495 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 751.440 902.775 752.040 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 909.495 455.770 913.495 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 909.495 754.770 913.495 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 909.495 133.770 913.495 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 909.495 660.470 913.495 ;
    END
  END user_irq[2]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 909.495 437.370 913.495 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 20.440 902.775 21.040 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 0.000 591.470 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 909.495 428.170 913.495 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 265.240 902.775 265.840 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 0.000 885.870 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.590 0.000 494.870 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 887.440 4.000 888.040 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 710.640 902.775 711.240 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 64.640 902.775 65.240 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 909.495 543.170 913.495 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 909.495 370.670 913.495 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 909.495 584.570 913.495 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 909.495 48.670 913.495 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 897.640 902.775 898.240 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 909.495 115.370 913.495 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 909.495 356.870 913.495 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 506.640 902.775 507.240 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 909.495 191.270 913.495 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 0.000 685.770 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.970 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 0.000 796.170 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 909.495 441.970 913.495 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 0.000 409.770 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 0.000 658.170 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 649.440 4.000 650.040 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 909.495 740.970 913.495 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 765.040 902.775 765.640 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 275.440 902.775 276.040 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 0.000 609.870 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 909.495 619.070 913.495 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.690 909.495 832.970 913.495 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 0.000 637.470 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 909.495 90.070 913.495 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 105.440 902.775 106.040 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 295.840 902.775 296.440 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 909.495 294.770 913.495 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 850.040 902.775 850.640 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 909.495 228.070 913.495 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 909.495 589.170 913.495 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 909.495 713.370 913.495 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 909.495 566.170 913.495 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 909.495 27.970 913.495 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 724.240 902.775 724.840 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 0.000 582.270 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.890 0.000 842.170 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 0.000 855.970 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.690 909.495 694.970 913.495 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 909.495 14.170 913.495 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 448.840 902.775 449.440 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 909.495 375.270 913.495 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 909.495 205.070 913.495 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 0.000 667.370 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 909.495 44.070 913.495 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.090 909.495 575.370 913.495 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 598.440 902.775 599.040 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.590 909.495 632.870 913.495 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 909.495 745.570 913.495 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 238.040 902.775 238.640 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 909.495 138.370 913.495 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 909.495 690.370 913.495 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 909.495 246.470 913.495 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 909.495 156.770 913.495 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.990 909.495 536.270 913.495 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 0.000 400.570 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 639.240 902.775 639.840 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 898.775 646.040 902.775 646.640 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 909.495 85.470 913.495 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 909.495 165.970 913.495 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 0.000 605.270 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 909.495 508.670 913.495 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 724.020 -9.320 727.020 920.520 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 544.020 -9.320 547.020 920.520 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 364.020 -9.320 367.020 920.520 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.020 -9.320 187.020 920.520 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 4.020 -9.320 7.020 920.520 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 909.500 -4.620 912.500 915.820 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 915.820 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -9.980 912.820 912.500 915.820 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 729.140 917.200 732.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 549.140 917.200 552.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 369.140 917.200 372.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 189.140 917.200 192.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 9.140 917.200 12.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -9.980 -4.620 912.500 -1.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 914.200 -9.320 917.200 920.520 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 814.020 -9.320 817.020 920.520 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 634.020 -9.320 637.020 920.520 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 454.020 -9.320 457.020 920.520 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 274.020 -9.320 277.020 920.520 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 94.020 -9.320 97.020 920.520 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 920.520 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 917.520 917.200 920.520 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 819.140 917.200 822.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 639.140 917.200 642.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 459.140 917.200 462.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 279.140 917.200 282.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 99.140 917.200 102.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 -9.320 917.200 -6.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 742.020 -18.720 745.020 929.920 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 562.020 -18.720 565.020 929.920 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 382.020 -18.720 385.020 929.920 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 202.020 -18.720 205.020 929.920 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.020 -18.720 25.020 929.920 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 918.900 -14.020 921.900 925.220 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 925.220 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -19.380 922.220 921.900 925.220 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 747.380 926.600 750.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 567.380 926.600 570.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 387.380 926.600 390.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 207.380 926.600 210.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 27.380 926.600 30.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -19.380 -14.020 921.900 -11.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 923.600 -18.720 926.600 929.920 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 832.020 -18.720 835.020 929.920 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 652.020 -18.720 655.020 929.920 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 472.020 -18.720 475.020 929.920 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 292.020 -18.720 295.020 929.920 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 112.020 -18.720 115.020 929.920 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 929.920 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 926.920 926.600 929.920 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 837.380 926.600 840.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 657.380 926.600 660.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 477.380 926.600 480.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 297.380 926.600 300.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 117.380 926.600 120.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 -18.720 926.600 -15.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 760.020 -28.120 763.020 939.320 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 580.020 -28.120 583.020 939.320 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 400.020 -28.120 403.020 939.320 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 220.020 -28.120 223.020 939.320 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 40.020 -28.120 43.020 939.320 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 928.300 -23.420 931.300 934.620 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 934.620 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -28.780 931.620 931.300 934.620 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 765.380 936.000 768.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 585.380 936.000 588.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 405.380 936.000 408.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 225.380 936.000 228.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 45.380 936.000 48.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -28.780 -23.420 931.300 -20.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 933.000 -28.120 936.000 939.320 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 850.020 -28.120 853.020 939.320 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 670.020 -28.120 673.020 939.320 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 490.020 -28.120 493.020 939.320 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 310.020 -28.120 313.020 939.320 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 130.020 -28.120 133.020 939.320 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 939.320 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 936.320 936.000 939.320 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 855.380 936.000 858.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 675.380 936.000 678.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 495.380 936.000 498.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 315.380 936.000 318.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 135.380 936.000 138.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 -28.120 936.000 -25.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 778.020 -37.520 781.020 948.720 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 598.020 -37.520 601.020 948.720 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 418.020 -37.520 421.020 948.720 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 238.020 -37.520 241.020 948.720 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 58.020 -37.520 61.020 948.720 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 937.700 -32.820 940.700 944.020 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 944.020 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -38.180 941.020 940.700 944.020 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 783.380 945.400 786.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 603.380 945.400 606.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 423.380 945.400 426.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 243.380 945.400 246.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 63.380 945.400 66.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -38.180 -32.820 940.700 -29.820 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 942.400 -37.520 945.400 948.720 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 868.020 -37.520 871.020 948.720 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 688.020 -37.520 691.020 948.720 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 508.020 -37.520 511.020 948.720 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 328.020 -37.520 331.020 948.720 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 148.020 -37.520 151.020 948.720 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 948.720 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 945.720 945.400 948.720 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 873.380 945.400 876.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 693.380 945.400 696.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 513.380 945.400 516.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 333.380 945.400 336.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 153.380 945.400 156.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 -37.520 945.400 -34.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 4.745 11.305 896.395 899.215 ;
      LAYER met1 ;
        RECT 4.685 10.640 899.690 900.560 ;
      LAYER met2 ;
        RECT 6.080 909.215 9.010 909.495 ;
        RECT 9.850 909.215 13.610 909.495 ;
        RECT 14.450 909.215 18.210 909.495 ;
        RECT 19.050 909.215 22.810 909.495 ;
        RECT 23.650 909.215 27.410 909.495 ;
        RECT 28.250 909.215 32.010 909.495 ;
        RECT 32.850 909.215 38.910 909.495 ;
        RECT 39.750 909.215 43.510 909.495 ;
        RECT 44.350 909.215 48.110 909.495 ;
        RECT 48.950 909.215 52.710 909.495 ;
        RECT 53.550 909.215 57.310 909.495 ;
        RECT 58.150 909.215 61.910 909.495 ;
        RECT 62.750 909.215 66.510 909.495 ;
        RECT 67.350 909.215 71.110 909.495 ;
        RECT 71.950 909.215 75.710 909.495 ;
        RECT 76.550 909.215 80.310 909.495 ;
        RECT 81.150 909.215 84.910 909.495 ;
        RECT 85.750 909.215 89.510 909.495 ;
        RECT 90.350 909.215 94.110 909.495 ;
        RECT 94.950 909.215 98.710 909.495 ;
        RECT 99.550 909.215 103.310 909.495 ;
        RECT 104.150 909.215 110.210 909.495 ;
        RECT 111.050 909.215 114.810 909.495 ;
        RECT 115.650 909.215 119.410 909.495 ;
        RECT 120.250 909.215 124.010 909.495 ;
        RECT 124.850 909.215 128.610 909.495 ;
        RECT 129.450 909.215 133.210 909.495 ;
        RECT 134.050 909.215 137.810 909.495 ;
        RECT 138.650 909.215 142.410 909.495 ;
        RECT 143.250 909.215 147.010 909.495 ;
        RECT 147.850 909.215 151.610 909.495 ;
        RECT 152.450 909.215 156.210 909.495 ;
        RECT 157.050 909.215 160.810 909.495 ;
        RECT 161.650 909.215 165.410 909.495 ;
        RECT 166.250 909.215 170.010 909.495 ;
        RECT 170.850 909.215 174.610 909.495 ;
        RECT 175.450 909.215 181.510 909.495 ;
        RECT 182.350 909.215 186.110 909.495 ;
        RECT 186.950 909.215 190.710 909.495 ;
        RECT 191.550 909.215 195.310 909.495 ;
        RECT 196.150 909.215 199.910 909.495 ;
        RECT 200.750 909.215 204.510 909.495 ;
        RECT 205.350 909.215 209.110 909.495 ;
        RECT 209.950 909.215 213.710 909.495 ;
        RECT 214.550 909.215 218.310 909.495 ;
        RECT 219.150 909.215 222.910 909.495 ;
        RECT 223.750 909.215 227.510 909.495 ;
        RECT 228.350 909.215 232.110 909.495 ;
        RECT 232.950 909.215 236.710 909.495 ;
        RECT 237.550 909.215 241.310 909.495 ;
        RECT 242.150 909.215 245.910 909.495 ;
        RECT 246.750 909.215 250.510 909.495 ;
        RECT 251.350 909.215 257.410 909.495 ;
        RECT 258.250 909.215 262.010 909.495 ;
        RECT 262.850 909.215 266.610 909.495 ;
        RECT 267.450 909.215 271.210 909.495 ;
        RECT 272.050 909.215 275.810 909.495 ;
        RECT 276.650 909.215 280.410 909.495 ;
        RECT 281.250 909.215 285.010 909.495 ;
        RECT 285.850 909.215 289.610 909.495 ;
        RECT 290.450 909.215 294.210 909.495 ;
        RECT 295.050 909.215 298.810 909.495 ;
        RECT 299.650 909.215 303.410 909.495 ;
        RECT 304.250 909.215 308.010 909.495 ;
        RECT 308.850 909.215 312.610 909.495 ;
        RECT 313.450 909.215 317.210 909.495 ;
        RECT 318.050 909.215 321.810 909.495 ;
        RECT 322.650 909.215 328.710 909.495 ;
        RECT 329.550 909.215 333.310 909.495 ;
        RECT 334.150 909.215 337.910 909.495 ;
        RECT 338.750 909.215 342.510 909.495 ;
        RECT 343.350 909.215 347.110 909.495 ;
        RECT 347.950 909.215 351.710 909.495 ;
        RECT 352.550 909.215 356.310 909.495 ;
        RECT 357.150 909.215 360.910 909.495 ;
        RECT 361.750 909.215 365.510 909.495 ;
        RECT 366.350 909.215 370.110 909.495 ;
        RECT 370.950 909.215 374.710 909.495 ;
        RECT 375.550 909.215 379.310 909.495 ;
        RECT 380.150 909.215 383.910 909.495 ;
        RECT 384.750 909.215 388.510 909.495 ;
        RECT 389.350 909.215 393.110 909.495 ;
        RECT 393.950 909.215 400.010 909.495 ;
        RECT 400.850 909.215 404.610 909.495 ;
        RECT 405.450 909.215 409.210 909.495 ;
        RECT 410.050 909.215 413.810 909.495 ;
        RECT 414.650 909.215 418.410 909.495 ;
        RECT 419.250 909.215 423.010 909.495 ;
        RECT 423.850 909.215 427.610 909.495 ;
        RECT 428.450 909.215 432.210 909.495 ;
        RECT 433.050 909.215 436.810 909.495 ;
        RECT 437.650 909.215 441.410 909.495 ;
        RECT 442.250 909.215 446.010 909.495 ;
        RECT 446.850 909.215 450.610 909.495 ;
        RECT 451.450 909.215 455.210 909.495 ;
        RECT 456.050 909.215 459.810 909.495 ;
        RECT 460.650 909.215 464.410 909.495 ;
        RECT 465.250 909.215 471.310 909.495 ;
        RECT 472.150 909.215 475.910 909.495 ;
        RECT 476.750 909.215 480.510 909.495 ;
        RECT 481.350 909.215 485.110 909.495 ;
        RECT 485.950 909.215 489.710 909.495 ;
        RECT 490.550 909.215 494.310 909.495 ;
        RECT 495.150 909.215 498.910 909.495 ;
        RECT 499.750 909.215 503.510 909.495 ;
        RECT 504.350 909.215 508.110 909.495 ;
        RECT 508.950 909.215 512.710 909.495 ;
        RECT 513.550 909.215 517.310 909.495 ;
        RECT 518.150 909.215 521.910 909.495 ;
        RECT 522.750 909.215 526.510 909.495 ;
        RECT 527.350 909.215 531.110 909.495 ;
        RECT 531.950 909.215 535.710 909.495 ;
        RECT 536.550 909.215 542.610 909.495 ;
        RECT 543.450 909.215 547.210 909.495 ;
        RECT 548.050 909.215 551.810 909.495 ;
        RECT 552.650 909.215 556.410 909.495 ;
        RECT 557.250 909.215 561.010 909.495 ;
        RECT 561.850 909.215 565.610 909.495 ;
        RECT 566.450 909.215 570.210 909.495 ;
        RECT 571.050 909.215 574.810 909.495 ;
        RECT 575.650 909.215 579.410 909.495 ;
        RECT 580.250 909.215 584.010 909.495 ;
        RECT 584.850 909.215 588.610 909.495 ;
        RECT 589.450 909.215 593.210 909.495 ;
        RECT 594.050 909.215 597.810 909.495 ;
        RECT 598.650 909.215 602.410 909.495 ;
        RECT 603.250 909.215 607.010 909.495 ;
        RECT 607.850 909.215 613.910 909.495 ;
        RECT 614.750 909.215 618.510 909.495 ;
        RECT 619.350 909.215 623.110 909.495 ;
        RECT 623.950 909.215 627.710 909.495 ;
        RECT 628.550 909.215 632.310 909.495 ;
        RECT 633.150 909.215 636.910 909.495 ;
        RECT 637.750 909.215 641.510 909.495 ;
        RECT 642.350 909.215 646.110 909.495 ;
        RECT 646.950 909.215 650.710 909.495 ;
        RECT 651.550 909.215 655.310 909.495 ;
        RECT 656.150 909.215 659.910 909.495 ;
        RECT 660.750 909.215 664.510 909.495 ;
        RECT 665.350 909.215 669.110 909.495 ;
        RECT 669.950 909.215 673.710 909.495 ;
        RECT 674.550 909.215 678.310 909.495 ;
        RECT 679.150 909.215 682.910 909.495 ;
        RECT 683.750 909.215 689.810 909.495 ;
        RECT 690.650 909.215 694.410 909.495 ;
        RECT 695.250 909.215 699.010 909.495 ;
        RECT 699.850 909.215 703.610 909.495 ;
        RECT 704.450 909.215 708.210 909.495 ;
        RECT 709.050 909.215 712.810 909.495 ;
        RECT 713.650 909.215 717.410 909.495 ;
        RECT 718.250 909.215 722.010 909.495 ;
        RECT 722.850 909.215 726.610 909.495 ;
        RECT 727.450 909.215 731.210 909.495 ;
        RECT 732.050 909.215 735.810 909.495 ;
        RECT 736.650 909.215 740.410 909.495 ;
        RECT 741.250 909.215 745.010 909.495 ;
        RECT 745.850 909.215 749.610 909.495 ;
        RECT 750.450 909.215 754.210 909.495 ;
        RECT 755.050 909.215 761.110 909.495 ;
        RECT 761.950 909.215 765.710 909.495 ;
        RECT 766.550 909.215 770.310 909.495 ;
        RECT 771.150 909.215 774.910 909.495 ;
        RECT 775.750 909.215 779.510 909.495 ;
        RECT 780.350 909.215 784.110 909.495 ;
        RECT 784.950 909.215 788.710 909.495 ;
        RECT 789.550 909.215 793.310 909.495 ;
        RECT 794.150 909.215 797.910 909.495 ;
        RECT 798.750 909.215 802.510 909.495 ;
        RECT 803.350 909.215 807.110 909.495 ;
        RECT 807.950 909.215 811.710 909.495 ;
        RECT 812.550 909.215 816.310 909.495 ;
        RECT 817.150 909.215 820.910 909.495 ;
        RECT 821.750 909.215 825.510 909.495 ;
        RECT 826.350 909.215 832.410 909.495 ;
        RECT 833.250 909.215 837.010 909.495 ;
        RECT 837.850 909.215 841.610 909.495 ;
        RECT 842.450 909.215 846.210 909.495 ;
        RECT 847.050 909.215 850.810 909.495 ;
        RECT 851.650 909.215 855.410 909.495 ;
        RECT 856.250 909.215 860.010 909.495 ;
        RECT 860.850 909.215 864.610 909.495 ;
        RECT 865.450 909.215 869.210 909.495 ;
        RECT 870.050 909.215 873.810 909.495 ;
        RECT 874.650 909.215 878.410 909.495 ;
        RECT 879.250 909.215 883.010 909.495 ;
        RECT 883.850 909.215 887.610 909.495 ;
        RECT 888.450 909.215 892.210 909.495 ;
        RECT 893.050 909.215 896.810 909.495 ;
        RECT 897.650 909.215 899.660 909.495 ;
        RECT 6.080 4.280 899.660 909.215 ;
        RECT 6.080 4.000 6.710 4.280 ;
        RECT 7.550 4.000 11.310 4.280 ;
        RECT 12.150 4.000 15.910 4.280 ;
        RECT 16.750 4.000 20.510 4.280 ;
        RECT 21.350 4.000 25.110 4.280 ;
        RECT 25.950 4.000 29.710 4.280 ;
        RECT 30.550 4.000 34.310 4.280 ;
        RECT 35.150 4.000 38.910 4.280 ;
        RECT 39.750 4.000 43.510 4.280 ;
        RECT 44.350 4.000 48.110 4.280 ;
        RECT 48.950 4.000 52.710 4.280 ;
        RECT 53.550 4.000 57.310 4.280 ;
        RECT 58.150 4.000 61.910 4.280 ;
        RECT 62.750 4.000 66.510 4.280 ;
        RECT 67.350 4.000 71.110 4.280 ;
        RECT 71.950 4.000 78.010 4.280 ;
        RECT 78.850 4.000 82.610 4.280 ;
        RECT 83.450 4.000 87.210 4.280 ;
        RECT 88.050 4.000 91.810 4.280 ;
        RECT 92.650 4.000 96.410 4.280 ;
        RECT 97.250 4.000 101.010 4.280 ;
        RECT 101.850 4.000 105.610 4.280 ;
        RECT 106.450 4.000 110.210 4.280 ;
        RECT 111.050 4.000 114.810 4.280 ;
        RECT 115.650 4.000 119.410 4.280 ;
        RECT 120.250 4.000 124.010 4.280 ;
        RECT 124.850 4.000 128.610 4.280 ;
        RECT 129.450 4.000 133.210 4.280 ;
        RECT 134.050 4.000 137.810 4.280 ;
        RECT 138.650 4.000 142.410 4.280 ;
        RECT 143.250 4.000 149.310 4.280 ;
        RECT 150.150 4.000 153.910 4.280 ;
        RECT 154.750 4.000 158.510 4.280 ;
        RECT 159.350 4.000 163.110 4.280 ;
        RECT 163.950 4.000 167.710 4.280 ;
        RECT 168.550 4.000 172.310 4.280 ;
        RECT 173.150 4.000 176.910 4.280 ;
        RECT 177.750 4.000 181.510 4.280 ;
        RECT 182.350 4.000 186.110 4.280 ;
        RECT 186.950 4.000 190.710 4.280 ;
        RECT 191.550 4.000 195.310 4.280 ;
        RECT 196.150 4.000 199.910 4.280 ;
        RECT 200.750 4.000 204.510 4.280 ;
        RECT 205.350 4.000 209.110 4.280 ;
        RECT 209.950 4.000 213.710 4.280 ;
        RECT 214.550 4.000 220.610 4.280 ;
        RECT 221.450 4.000 225.210 4.280 ;
        RECT 226.050 4.000 229.810 4.280 ;
        RECT 230.650 4.000 234.410 4.280 ;
        RECT 235.250 4.000 239.010 4.280 ;
        RECT 239.850 4.000 243.610 4.280 ;
        RECT 244.450 4.000 248.210 4.280 ;
        RECT 249.050 4.000 252.810 4.280 ;
        RECT 253.650 4.000 257.410 4.280 ;
        RECT 258.250 4.000 262.010 4.280 ;
        RECT 262.850 4.000 266.610 4.280 ;
        RECT 267.450 4.000 271.210 4.280 ;
        RECT 272.050 4.000 275.810 4.280 ;
        RECT 276.650 4.000 280.410 4.280 ;
        RECT 281.250 4.000 285.010 4.280 ;
        RECT 285.850 4.000 291.910 4.280 ;
        RECT 292.750 4.000 296.510 4.280 ;
        RECT 297.350 4.000 301.110 4.280 ;
        RECT 301.950 4.000 305.710 4.280 ;
        RECT 306.550 4.000 310.310 4.280 ;
        RECT 311.150 4.000 314.910 4.280 ;
        RECT 315.750 4.000 319.510 4.280 ;
        RECT 320.350 4.000 324.110 4.280 ;
        RECT 324.950 4.000 328.710 4.280 ;
        RECT 329.550 4.000 333.310 4.280 ;
        RECT 334.150 4.000 337.910 4.280 ;
        RECT 338.750 4.000 342.510 4.280 ;
        RECT 343.350 4.000 347.110 4.280 ;
        RECT 347.950 4.000 351.710 4.280 ;
        RECT 352.550 4.000 356.310 4.280 ;
        RECT 357.150 4.000 363.210 4.280 ;
        RECT 364.050 4.000 367.810 4.280 ;
        RECT 368.650 4.000 372.410 4.280 ;
        RECT 373.250 4.000 377.010 4.280 ;
        RECT 377.850 4.000 381.610 4.280 ;
        RECT 382.450 4.000 386.210 4.280 ;
        RECT 387.050 4.000 390.810 4.280 ;
        RECT 391.650 4.000 395.410 4.280 ;
        RECT 396.250 4.000 400.010 4.280 ;
        RECT 400.850 4.000 404.610 4.280 ;
        RECT 405.450 4.000 409.210 4.280 ;
        RECT 410.050 4.000 413.810 4.280 ;
        RECT 414.650 4.000 418.410 4.280 ;
        RECT 419.250 4.000 423.010 4.280 ;
        RECT 423.850 4.000 427.610 4.280 ;
        RECT 428.450 4.000 434.510 4.280 ;
        RECT 435.350 4.000 439.110 4.280 ;
        RECT 439.950 4.000 443.710 4.280 ;
        RECT 444.550 4.000 448.310 4.280 ;
        RECT 449.150 4.000 452.910 4.280 ;
        RECT 453.750 4.000 457.510 4.280 ;
        RECT 458.350 4.000 462.110 4.280 ;
        RECT 462.950 4.000 466.710 4.280 ;
        RECT 467.550 4.000 471.310 4.280 ;
        RECT 472.150 4.000 475.910 4.280 ;
        RECT 476.750 4.000 480.510 4.280 ;
        RECT 481.350 4.000 485.110 4.280 ;
        RECT 485.950 4.000 489.710 4.280 ;
        RECT 490.550 4.000 494.310 4.280 ;
        RECT 495.150 4.000 498.910 4.280 ;
        RECT 499.750 4.000 503.510 4.280 ;
        RECT 504.350 4.000 510.410 4.280 ;
        RECT 511.250 4.000 515.010 4.280 ;
        RECT 515.850 4.000 519.610 4.280 ;
        RECT 520.450 4.000 524.210 4.280 ;
        RECT 525.050 4.000 528.810 4.280 ;
        RECT 529.650 4.000 533.410 4.280 ;
        RECT 534.250 4.000 538.010 4.280 ;
        RECT 538.850 4.000 542.610 4.280 ;
        RECT 543.450 4.000 547.210 4.280 ;
        RECT 548.050 4.000 551.810 4.280 ;
        RECT 552.650 4.000 556.410 4.280 ;
        RECT 557.250 4.000 561.010 4.280 ;
        RECT 561.850 4.000 565.610 4.280 ;
        RECT 566.450 4.000 570.210 4.280 ;
        RECT 571.050 4.000 574.810 4.280 ;
        RECT 575.650 4.000 581.710 4.280 ;
        RECT 582.550 4.000 586.310 4.280 ;
        RECT 587.150 4.000 590.910 4.280 ;
        RECT 591.750 4.000 595.510 4.280 ;
        RECT 596.350 4.000 600.110 4.280 ;
        RECT 600.950 4.000 604.710 4.280 ;
        RECT 605.550 4.000 609.310 4.280 ;
        RECT 610.150 4.000 613.910 4.280 ;
        RECT 614.750 4.000 618.510 4.280 ;
        RECT 619.350 4.000 623.110 4.280 ;
        RECT 623.950 4.000 627.710 4.280 ;
        RECT 628.550 4.000 632.310 4.280 ;
        RECT 633.150 4.000 636.910 4.280 ;
        RECT 637.750 4.000 641.510 4.280 ;
        RECT 642.350 4.000 646.110 4.280 ;
        RECT 646.950 4.000 653.010 4.280 ;
        RECT 653.850 4.000 657.610 4.280 ;
        RECT 658.450 4.000 662.210 4.280 ;
        RECT 663.050 4.000 666.810 4.280 ;
        RECT 667.650 4.000 671.410 4.280 ;
        RECT 672.250 4.000 676.010 4.280 ;
        RECT 676.850 4.000 680.610 4.280 ;
        RECT 681.450 4.000 685.210 4.280 ;
        RECT 686.050 4.000 689.810 4.280 ;
        RECT 690.650 4.000 694.410 4.280 ;
        RECT 695.250 4.000 699.010 4.280 ;
        RECT 699.850 4.000 703.610 4.280 ;
        RECT 704.450 4.000 708.210 4.280 ;
        RECT 709.050 4.000 712.810 4.280 ;
        RECT 713.650 4.000 717.410 4.280 ;
        RECT 718.250 4.000 724.310 4.280 ;
        RECT 725.150 4.000 728.910 4.280 ;
        RECT 729.750 4.000 733.510 4.280 ;
        RECT 734.350 4.000 738.110 4.280 ;
        RECT 738.950 4.000 742.710 4.280 ;
        RECT 743.550 4.000 747.310 4.280 ;
        RECT 748.150 4.000 751.910 4.280 ;
        RECT 752.750 4.000 756.510 4.280 ;
        RECT 757.350 4.000 761.110 4.280 ;
        RECT 761.950 4.000 765.710 4.280 ;
        RECT 766.550 4.000 770.310 4.280 ;
        RECT 771.150 4.000 774.910 4.280 ;
        RECT 775.750 4.000 779.510 4.280 ;
        RECT 780.350 4.000 784.110 4.280 ;
        RECT 784.950 4.000 788.710 4.280 ;
        RECT 789.550 4.000 795.610 4.280 ;
        RECT 796.450 4.000 800.210 4.280 ;
        RECT 801.050 4.000 804.810 4.280 ;
        RECT 805.650 4.000 809.410 4.280 ;
        RECT 810.250 4.000 814.010 4.280 ;
        RECT 814.850 4.000 818.610 4.280 ;
        RECT 819.450 4.000 823.210 4.280 ;
        RECT 824.050 4.000 827.810 4.280 ;
        RECT 828.650 4.000 832.410 4.280 ;
        RECT 833.250 4.000 837.010 4.280 ;
        RECT 837.850 4.000 841.610 4.280 ;
        RECT 842.450 4.000 846.210 4.280 ;
        RECT 847.050 4.000 850.810 4.280 ;
        RECT 851.650 4.000 855.410 4.280 ;
        RECT 856.250 4.000 860.010 4.280 ;
        RECT 860.850 4.000 866.910 4.280 ;
        RECT 867.750 4.000 871.510 4.280 ;
        RECT 872.350 4.000 876.110 4.280 ;
        RECT 876.950 4.000 880.710 4.280 ;
        RECT 881.550 4.000 885.310 4.280 ;
        RECT 886.150 4.000 889.910 4.280 ;
        RECT 890.750 4.000 894.510 4.280 ;
        RECT 895.350 4.000 899.110 4.280 ;
      LAYER met3 ;
        RECT 4.000 904.040 898.375 904.905 ;
        RECT 4.000 902.040 898.775 904.040 ;
        RECT 4.400 900.640 898.775 902.040 ;
        RECT 4.000 898.640 898.775 900.640 ;
        RECT 4.000 897.240 898.375 898.640 ;
        RECT 4.000 895.240 898.775 897.240 ;
        RECT 4.400 893.840 898.775 895.240 ;
        RECT 4.000 891.840 898.775 893.840 ;
        RECT 4.000 890.440 898.375 891.840 ;
        RECT 4.000 888.440 898.775 890.440 ;
        RECT 4.400 887.040 898.775 888.440 ;
        RECT 4.000 885.040 898.775 887.040 ;
        RECT 4.000 883.640 898.375 885.040 ;
        RECT 4.000 881.640 898.775 883.640 ;
        RECT 4.400 880.240 898.775 881.640 ;
        RECT 4.000 878.240 898.775 880.240 ;
        RECT 4.000 876.840 898.375 878.240 ;
        RECT 4.000 874.840 898.775 876.840 ;
        RECT 4.400 873.440 898.775 874.840 ;
        RECT 4.000 871.440 898.775 873.440 ;
        RECT 4.000 870.040 898.375 871.440 ;
        RECT 4.000 868.040 898.775 870.040 ;
        RECT 4.400 866.640 898.775 868.040 ;
        RECT 4.000 864.640 898.775 866.640 ;
        RECT 4.000 863.240 898.375 864.640 ;
        RECT 4.000 861.240 898.775 863.240 ;
        RECT 4.400 859.840 898.775 861.240 ;
        RECT 4.000 857.840 898.775 859.840 ;
        RECT 4.000 856.440 898.375 857.840 ;
        RECT 4.000 851.040 898.775 856.440 ;
        RECT 4.400 849.640 898.375 851.040 ;
        RECT 4.000 844.240 898.775 849.640 ;
        RECT 4.400 842.840 898.375 844.240 ;
        RECT 4.000 837.440 898.775 842.840 ;
        RECT 4.400 836.040 898.375 837.440 ;
        RECT 4.000 830.640 898.775 836.040 ;
        RECT 4.400 829.240 898.375 830.640 ;
        RECT 4.000 823.840 898.775 829.240 ;
        RECT 4.400 822.440 898.375 823.840 ;
        RECT 4.000 817.040 898.775 822.440 ;
        RECT 4.400 815.640 898.375 817.040 ;
        RECT 4.000 810.240 898.775 815.640 ;
        RECT 4.400 808.840 898.375 810.240 ;
        RECT 4.000 803.440 898.775 808.840 ;
        RECT 4.400 802.040 898.775 803.440 ;
        RECT 4.000 800.040 898.775 802.040 ;
        RECT 4.000 798.640 898.375 800.040 ;
        RECT 4.000 796.640 898.775 798.640 ;
        RECT 4.400 795.240 898.775 796.640 ;
        RECT 4.000 793.240 898.775 795.240 ;
        RECT 4.000 791.840 898.375 793.240 ;
        RECT 4.000 789.840 898.775 791.840 ;
        RECT 4.400 788.440 898.775 789.840 ;
        RECT 4.000 786.440 898.775 788.440 ;
        RECT 4.000 785.040 898.375 786.440 ;
        RECT 4.000 783.040 898.775 785.040 ;
        RECT 4.400 781.640 898.775 783.040 ;
        RECT 4.000 779.640 898.775 781.640 ;
        RECT 4.000 778.240 898.375 779.640 ;
        RECT 4.000 776.240 898.775 778.240 ;
        RECT 4.400 774.840 898.775 776.240 ;
        RECT 4.000 772.840 898.775 774.840 ;
        RECT 4.000 771.440 898.375 772.840 ;
        RECT 4.000 769.440 898.775 771.440 ;
        RECT 4.400 768.040 898.775 769.440 ;
        RECT 4.000 766.040 898.775 768.040 ;
        RECT 4.000 764.640 898.375 766.040 ;
        RECT 4.000 762.640 898.775 764.640 ;
        RECT 4.400 761.240 898.775 762.640 ;
        RECT 4.000 759.240 898.775 761.240 ;
        RECT 4.000 757.840 898.375 759.240 ;
        RECT 4.000 755.840 898.775 757.840 ;
        RECT 4.400 754.440 898.775 755.840 ;
        RECT 4.000 752.440 898.775 754.440 ;
        RECT 4.000 751.040 898.375 752.440 ;
        RECT 4.000 745.640 898.775 751.040 ;
        RECT 4.400 744.240 898.375 745.640 ;
        RECT 4.000 738.840 898.775 744.240 ;
        RECT 4.400 737.440 898.375 738.840 ;
        RECT 4.000 732.040 898.775 737.440 ;
        RECT 4.400 730.640 898.375 732.040 ;
        RECT 4.000 725.240 898.775 730.640 ;
        RECT 4.400 723.840 898.375 725.240 ;
        RECT 4.000 718.440 898.775 723.840 ;
        RECT 4.400 717.040 898.375 718.440 ;
        RECT 4.000 711.640 898.775 717.040 ;
        RECT 4.400 710.240 898.375 711.640 ;
        RECT 4.000 704.840 898.775 710.240 ;
        RECT 4.400 703.440 898.375 704.840 ;
        RECT 4.000 698.040 898.775 703.440 ;
        RECT 4.400 696.640 898.775 698.040 ;
        RECT 4.000 694.640 898.775 696.640 ;
        RECT 4.000 693.240 898.375 694.640 ;
        RECT 4.000 691.240 898.775 693.240 ;
        RECT 4.400 689.840 898.775 691.240 ;
        RECT 4.000 687.840 898.775 689.840 ;
        RECT 4.000 686.440 898.375 687.840 ;
        RECT 4.000 684.440 898.775 686.440 ;
        RECT 4.400 683.040 898.775 684.440 ;
        RECT 4.000 681.040 898.775 683.040 ;
        RECT 4.000 679.640 898.375 681.040 ;
        RECT 4.000 677.640 898.775 679.640 ;
        RECT 4.400 676.240 898.775 677.640 ;
        RECT 4.000 674.240 898.775 676.240 ;
        RECT 4.000 672.840 898.375 674.240 ;
        RECT 4.000 670.840 898.775 672.840 ;
        RECT 4.400 669.440 898.775 670.840 ;
        RECT 4.000 667.440 898.775 669.440 ;
        RECT 4.000 666.040 898.375 667.440 ;
        RECT 4.000 664.040 898.775 666.040 ;
        RECT 4.400 662.640 898.775 664.040 ;
        RECT 4.000 660.640 898.775 662.640 ;
        RECT 4.000 659.240 898.375 660.640 ;
        RECT 4.000 657.240 898.775 659.240 ;
        RECT 4.400 655.840 898.775 657.240 ;
        RECT 4.000 653.840 898.775 655.840 ;
        RECT 4.000 652.440 898.375 653.840 ;
        RECT 4.000 650.440 898.775 652.440 ;
        RECT 4.400 649.040 898.775 650.440 ;
        RECT 4.000 647.040 898.775 649.040 ;
        RECT 4.000 645.640 898.375 647.040 ;
        RECT 4.000 640.240 898.775 645.640 ;
        RECT 4.400 638.840 898.375 640.240 ;
        RECT 4.000 633.440 898.775 638.840 ;
        RECT 4.400 632.040 898.375 633.440 ;
        RECT 4.000 626.640 898.775 632.040 ;
        RECT 4.400 625.240 898.375 626.640 ;
        RECT 4.000 619.840 898.775 625.240 ;
        RECT 4.400 618.440 898.375 619.840 ;
        RECT 4.000 613.040 898.775 618.440 ;
        RECT 4.400 611.640 898.375 613.040 ;
        RECT 4.000 606.240 898.775 611.640 ;
        RECT 4.400 604.840 898.375 606.240 ;
        RECT 4.000 599.440 898.775 604.840 ;
        RECT 4.400 598.040 898.375 599.440 ;
        RECT 4.000 592.640 898.775 598.040 ;
        RECT 4.400 591.240 898.375 592.640 ;
        RECT 4.000 585.840 898.775 591.240 ;
        RECT 4.400 584.440 898.775 585.840 ;
        RECT 4.000 582.440 898.775 584.440 ;
        RECT 4.000 581.040 898.375 582.440 ;
        RECT 4.000 579.040 898.775 581.040 ;
        RECT 4.400 577.640 898.775 579.040 ;
        RECT 4.000 575.640 898.775 577.640 ;
        RECT 4.000 574.240 898.375 575.640 ;
        RECT 4.000 572.240 898.775 574.240 ;
        RECT 4.400 570.840 898.775 572.240 ;
        RECT 4.000 568.840 898.775 570.840 ;
        RECT 4.000 567.440 898.375 568.840 ;
        RECT 4.000 565.440 898.775 567.440 ;
        RECT 4.400 564.040 898.775 565.440 ;
        RECT 4.000 562.040 898.775 564.040 ;
        RECT 4.000 560.640 898.375 562.040 ;
        RECT 4.000 558.640 898.775 560.640 ;
        RECT 4.400 557.240 898.775 558.640 ;
        RECT 4.000 555.240 898.775 557.240 ;
        RECT 4.000 553.840 898.375 555.240 ;
        RECT 4.000 551.840 898.775 553.840 ;
        RECT 4.400 550.440 898.775 551.840 ;
        RECT 4.000 548.440 898.775 550.440 ;
        RECT 4.000 547.040 898.375 548.440 ;
        RECT 4.000 545.040 898.775 547.040 ;
        RECT 4.400 543.640 898.775 545.040 ;
        RECT 4.000 541.640 898.775 543.640 ;
        RECT 4.000 540.240 898.375 541.640 ;
        RECT 4.000 538.240 898.775 540.240 ;
        RECT 4.400 536.840 898.775 538.240 ;
        RECT 4.000 534.840 898.775 536.840 ;
        RECT 4.000 533.440 898.375 534.840 ;
        RECT 4.000 528.040 898.775 533.440 ;
        RECT 4.400 526.640 898.375 528.040 ;
        RECT 4.000 521.240 898.775 526.640 ;
        RECT 4.400 519.840 898.375 521.240 ;
        RECT 4.000 514.440 898.775 519.840 ;
        RECT 4.400 513.040 898.375 514.440 ;
        RECT 4.000 507.640 898.775 513.040 ;
        RECT 4.400 506.240 898.375 507.640 ;
        RECT 4.000 500.840 898.775 506.240 ;
        RECT 4.400 499.440 898.375 500.840 ;
        RECT 4.000 494.040 898.775 499.440 ;
        RECT 4.400 492.640 898.375 494.040 ;
        RECT 4.000 487.240 898.775 492.640 ;
        RECT 4.400 485.840 898.375 487.240 ;
        RECT 4.000 480.440 898.775 485.840 ;
        RECT 4.400 479.040 898.775 480.440 ;
        RECT 4.000 477.040 898.775 479.040 ;
        RECT 4.000 475.640 898.375 477.040 ;
        RECT 4.000 473.640 898.775 475.640 ;
        RECT 4.400 472.240 898.775 473.640 ;
        RECT 4.000 470.240 898.775 472.240 ;
        RECT 4.000 468.840 898.375 470.240 ;
        RECT 4.000 466.840 898.775 468.840 ;
        RECT 4.400 465.440 898.775 466.840 ;
        RECT 4.000 463.440 898.775 465.440 ;
        RECT 4.000 462.040 898.375 463.440 ;
        RECT 4.000 460.040 898.775 462.040 ;
        RECT 4.400 458.640 898.775 460.040 ;
        RECT 4.000 456.640 898.775 458.640 ;
        RECT 4.000 455.240 898.375 456.640 ;
        RECT 4.000 453.240 898.775 455.240 ;
        RECT 4.400 451.840 898.775 453.240 ;
        RECT 4.000 449.840 898.775 451.840 ;
        RECT 4.000 448.440 898.375 449.840 ;
        RECT 4.000 446.440 898.775 448.440 ;
        RECT 4.400 445.040 898.775 446.440 ;
        RECT 4.000 443.040 898.775 445.040 ;
        RECT 4.000 441.640 898.375 443.040 ;
        RECT 4.000 439.640 898.775 441.640 ;
        RECT 4.400 438.240 898.775 439.640 ;
        RECT 4.000 436.240 898.775 438.240 ;
        RECT 4.000 434.840 898.375 436.240 ;
        RECT 4.000 432.840 898.775 434.840 ;
        RECT 4.400 431.440 898.775 432.840 ;
        RECT 4.000 429.440 898.775 431.440 ;
        RECT 4.000 428.040 898.375 429.440 ;
        RECT 4.000 422.640 898.775 428.040 ;
        RECT 4.400 421.240 898.375 422.640 ;
        RECT 4.000 415.840 898.775 421.240 ;
        RECT 4.400 414.440 898.375 415.840 ;
        RECT 4.000 409.040 898.775 414.440 ;
        RECT 4.400 407.640 898.375 409.040 ;
        RECT 4.000 402.240 898.775 407.640 ;
        RECT 4.400 400.840 898.375 402.240 ;
        RECT 4.000 395.440 898.775 400.840 ;
        RECT 4.400 394.040 898.375 395.440 ;
        RECT 4.000 388.640 898.775 394.040 ;
        RECT 4.400 387.240 898.375 388.640 ;
        RECT 4.000 381.840 898.775 387.240 ;
        RECT 4.400 380.440 898.375 381.840 ;
        RECT 4.000 375.040 898.775 380.440 ;
        RECT 4.400 373.640 898.775 375.040 ;
        RECT 4.000 371.640 898.775 373.640 ;
        RECT 4.000 370.240 898.375 371.640 ;
        RECT 4.000 368.240 898.775 370.240 ;
        RECT 4.400 366.840 898.775 368.240 ;
        RECT 4.000 364.840 898.775 366.840 ;
        RECT 4.000 363.440 898.375 364.840 ;
        RECT 4.000 361.440 898.775 363.440 ;
        RECT 4.400 360.040 898.775 361.440 ;
        RECT 4.000 358.040 898.775 360.040 ;
        RECT 4.000 356.640 898.375 358.040 ;
        RECT 4.000 354.640 898.775 356.640 ;
        RECT 4.400 353.240 898.775 354.640 ;
        RECT 4.000 351.240 898.775 353.240 ;
        RECT 4.000 349.840 898.375 351.240 ;
        RECT 4.000 347.840 898.775 349.840 ;
        RECT 4.400 346.440 898.775 347.840 ;
        RECT 4.000 344.440 898.775 346.440 ;
        RECT 4.000 343.040 898.375 344.440 ;
        RECT 4.000 341.040 898.775 343.040 ;
        RECT 4.400 339.640 898.775 341.040 ;
        RECT 4.000 337.640 898.775 339.640 ;
        RECT 4.000 336.240 898.375 337.640 ;
        RECT 4.000 334.240 898.775 336.240 ;
        RECT 4.400 332.840 898.775 334.240 ;
        RECT 4.000 330.840 898.775 332.840 ;
        RECT 4.000 329.440 898.375 330.840 ;
        RECT 4.000 327.440 898.775 329.440 ;
        RECT 4.400 326.040 898.775 327.440 ;
        RECT 4.000 324.040 898.775 326.040 ;
        RECT 4.000 322.640 898.375 324.040 ;
        RECT 4.000 317.240 898.775 322.640 ;
        RECT 4.400 315.840 898.375 317.240 ;
        RECT 4.000 310.440 898.775 315.840 ;
        RECT 4.400 309.040 898.375 310.440 ;
        RECT 4.000 303.640 898.775 309.040 ;
        RECT 4.400 302.240 898.375 303.640 ;
        RECT 4.000 296.840 898.775 302.240 ;
        RECT 4.400 295.440 898.375 296.840 ;
        RECT 4.000 290.040 898.775 295.440 ;
        RECT 4.400 288.640 898.375 290.040 ;
        RECT 4.000 283.240 898.775 288.640 ;
        RECT 4.400 281.840 898.375 283.240 ;
        RECT 4.000 276.440 898.775 281.840 ;
        RECT 4.400 275.040 898.375 276.440 ;
        RECT 4.000 269.640 898.775 275.040 ;
        RECT 4.400 268.240 898.775 269.640 ;
        RECT 4.000 266.240 898.775 268.240 ;
        RECT 4.000 264.840 898.375 266.240 ;
        RECT 4.000 262.840 898.775 264.840 ;
        RECT 4.400 261.440 898.775 262.840 ;
        RECT 4.000 259.440 898.775 261.440 ;
        RECT 4.000 258.040 898.375 259.440 ;
        RECT 4.000 256.040 898.775 258.040 ;
        RECT 4.400 254.640 898.775 256.040 ;
        RECT 4.000 252.640 898.775 254.640 ;
        RECT 4.000 251.240 898.375 252.640 ;
        RECT 4.000 249.240 898.775 251.240 ;
        RECT 4.400 247.840 898.775 249.240 ;
        RECT 4.000 245.840 898.775 247.840 ;
        RECT 4.000 244.440 898.375 245.840 ;
        RECT 4.000 242.440 898.775 244.440 ;
        RECT 4.400 241.040 898.775 242.440 ;
        RECT 4.000 239.040 898.775 241.040 ;
        RECT 4.000 237.640 898.375 239.040 ;
        RECT 4.000 235.640 898.775 237.640 ;
        RECT 4.400 234.240 898.775 235.640 ;
        RECT 4.000 232.240 898.775 234.240 ;
        RECT 4.000 230.840 898.375 232.240 ;
        RECT 4.000 228.840 898.775 230.840 ;
        RECT 4.400 227.440 898.775 228.840 ;
        RECT 4.000 225.440 898.775 227.440 ;
        RECT 4.000 224.040 898.375 225.440 ;
        RECT 4.000 222.040 898.775 224.040 ;
        RECT 4.400 220.640 898.775 222.040 ;
        RECT 4.000 218.640 898.775 220.640 ;
        RECT 4.000 217.240 898.375 218.640 ;
        RECT 4.000 211.840 898.775 217.240 ;
        RECT 4.400 210.440 898.375 211.840 ;
        RECT 4.000 205.040 898.775 210.440 ;
        RECT 4.400 203.640 898.375 205.040 ;
        RECT 4.000 198.240 898.775 203.640 ;
        RECT 4.400 196.840 898.375 198.240 ;
        RECT 4.000 191.440 898.775 196.840 ;
        RECT 4.400 190.040 898.375 191.440 ;
        RECT 4.000 184.640 898.775 190.040 ;
        RECT 4.400 183.240 898.375 184.640 ;
        RECT 4.000 177.840 898.775 183.240 ;
        RECT 4.400 176.440 898.375 177.840 ;
        RECT 4.000 171.040 898.775 176.440 ;
        RECT 4.400 169.640 898.375 171.040 ;
        RECT 4.000 164.240 898.775 169.640 ;
        RECT 4.400 162.840 898.775 164.240 ;
        RECT 4.000 160.840 898.775 162.840 ;
        RECT 4.000 159.440 898.375 160.840 ;
        RECT 4.000 157.440 898.775 159.440 ;
        RECT 4.400 156.040 898.775 157.440 ;
        RECT 4.000 154.040 898.775 156.040 ;
        RECT 4.000 152.640 898.375 154.040 ;
        RECT 4.000 150.640 898.775 152.640 ;
        RECT 4.400 149.240 898.775 150.640 ;
        RECT 4.000 147.240 898.775 149.240 ;
        RECT 4.000 145.840 898.375 147.240 ;
        RECT 4.000 143.840 898.775 145.840 ;
        RECT 4.400 142.440 898.775 143.840 ;
        RECT 4.000 140.440 898.775 142.440 ;
        RECT 4.000 139.040 898.375 140.440 ;
        RECT 4.000 137.040 898.775 139.040 ;
        RECT 4.400 135.640 898.775 137.040 ;
        RECT 4.000 133.640 898.775 135.640 ;
        RECT 4.000 132.240 898.375 133.640 ;
        RECT 4.000 130.240 898.775 132.240 ;
        RECT 4.400 128.840 898.775 130.240 ;
        RECT 4.000 126.840 898.775 128.840 ;
        RECT 4.000 125.440 898.375 126.840 ;
        RECT 4.000 123.440 898.775 125.440 ;
        RECT 4.400 122.040 898.775 123.440 ;
        RECT 4.000 120.040 898.775 122.040 ;
        RECT 4.000 118.640 898.375 120.040 ;
        RECT 4.000 116.640 898.775 118.640 ;
        RECT 4.400 115.240 898.775 116.640 ;
        RECT 4.000 113.240 898.775 115.240 ;
        RECT 4.000 111.840 898.375 113.240 ;
        RECT 4.000 106.440 898.775 111.840 ;
        RECT 4.400 105.040 898.375 106.440 ;
        RECT 4.000 99.640 898.775 105.040 ;
        RECT 4.400 98.240 898.375 99.640 ;
        RECT 4.000 92.840 898.775 98.240 ;
        RECT 4.400 91.440 898.375 92.840 ;
        RECT 4.000 86.040 898.775 91.440 ;
        RECT 4.400 84.640 898.375 86.040 ;
        RECT 4.000 79.240 898.775 84.640 ;
        RECT 4.400 77.840 898.375 79.240 ;
        RECT 4.000 72.440 898.775 77.840 ;
        RECT 4.400 71.040 898.375 72.440 ;
        RECT 4.000 65.640 898.775 71.040 ;
        RECT 4.400 64.240 898.375 65.640 ;
        RECT 4.000 58.840 898.775 64.240 ;
        RECT 4.400 57.440 898.775 58.840 ;
        RECT 4.000 55.440 898.775 57.440 ;
        RECT 4.000 54.040 898.375 55.440 ;
        RECT 4.000 52.040 898.775 54.040 ;
        RECT 4.400 50.640 898.775 52.040 ;
        RECT 4.000 48.640 898.775 50.640 ;
        RECT 4.000 47.240 898.375 48.640 ;
        RECT 4.000 45.240 898.775 47.240 ;
        RECT 4.400 43.840 898.775 45.240 ;
        RECT 4.000 41.840 898.775 43.840 ;
        RECT 4.000 40.440 898.375 41.840 ;
        RECT 4.000 38.440 898.775 40.440 ;
        RECT 4.400 37.040 898.775 38.440 ;
        RECT 4.000 35.040 898.775 37.040 ;
        RECT 4.000 33.640 898.375 35.040 ;
        RECT 4.000 31.640 898.775 33.640 ;
        RECT 4.400 30.240 898.775 31.640 ;
        RECT 4.000 28.240 898.775 30.240 ;
        RECT 4.000 26.840 898.375 28.240 ;
        RECT 4.000 24.840 898.775 26.840 ;
        RECT 4.400 23.440 898.775 24.840 ;
        RECT 4.000 21.440 898.775 23.440 ;
        RECT 4.000 20.040 898.375 21.440 ;
        RECT 4.000 18.040 898.775 20.040 ;
        RECT 4.400 16.640 898.775 18.040 ;
        RECT 4.000 14.640 898.775 16.640 ;
        RECT 4.000 13.240 898.375 14.640 ;
        RECT 4.000 11.240 898.775 13.240 ;
        RECT 4.400 9.840 898.775 11.240 ;
        RECT 4.000 7.840 898.775 9.840 ;
        RECT 4.000 6.975 898.375 7.840 ;
      LAYER met4 ;
        RECT 33.415 17.175 39.620 894.705 ;
        RECT 43.420 17.175 57.620 894.705 ;
        RECT 61.420 17.175 93.620 894.705 ;
        RECT 97.420 17.175 111.620 894.705 ;
        RECT 115.420 17.175 129.620 894.705 ;
        RECT 133.420 17.175 147.620 894.705 ;
        RECT 151.420 17.175 183.620 894.705 ;
        RECT 187.420 17.175 201.620 894.705 ;
        RECT 205.420 17.175 219.620 894.705 ;
        RECT 223.420 17.175 237.620 894.705 ;
        RECT 241.420 17.175 273.620 894.705 ;
        RECT 277.420 17.175 291.620 894.705 ;
        RECT 295.420 17.175 309.620 894.705 ;
        RECT 313.420 17.175 327.620 894.705 ;
        RECT 331.420 17.175 363.620 894.705 ;
        RECT 367.420 17.175 381.620 894.705 ;
        RECT 385.420 17.175 399.620 894.705 ;
        RECT 403.420 17.175 417.620 894.705 ;
        RECT 421.420 17.175 453.620 894.705 ;
        RECT 457.420 17.175 471.620 894.705 ;
        RECT 475.420 17.175 489.620 894.705 ;
        RECT 493.420 17.175 507.620 894.705 ;
        RECT 511.420 17.175 543.620 894.705 ;
        RECT 547.420 17.175 561.620 894.705 ;
        RECT 565.420 17.175 579.620 894.705 ;
        RECT 583.420 17.175 597.620 894.705 ;
        RECT 601.420 17.175 633.620 894.705 ;
        RECT 637.420 17.175 651.620 894.705 ;
        RECT 655.420 17.175 669.620 894.705 ;
        RECT 673.420 17.175 687.620 894.705 ;
        RECT 691.420 17.175 723.620 894.705 ;
        RECT 727.420 17.175 741.620 894.705 ;
        RECT 745.420 17.175 759.620 894.705 ;
        RECT 763.420 17.175 777.620 894.705 ;
        RECT 781.420 17.175 813.620 894.705 ;
        RECT 817.420 17.175 831.620 894.705 ;
        RECT 835.420 17.175 849.620 894.705 ;
        RECT 853.420 17.175 867.620 894.705 ;
        RECT 871.420 17.175 889.345 894.705 ;
      LAYER met5 ;
        RECT -42.880 948.720 -39.880 948.730 ;
        RECT 148.020 948.720 151.020 948.730 ;
        RECT 328.020 948.720 331.020 948.730 ;
        RECT 508.020 948.720 511.020 948.730 ;
        RECT 688.020 948.720 691.020 948.730 ;
        RECT 868.020 948.720 871.020 948.730 ;
        RECT 942.400 948.720 945.400 948.730 ;
        RECT -42.880 945.710 -39.880 945.720 ;
        RECT 148.020 945.710 151.020 945.720 ;
        RECT 328.020 945.710 331.020 945.720 ;
        RECT 508.020 945.710 511.020 945.720 ;
        RECT 688.020 945.710 691.020 945.720 ;
        RECT 868.020 945.710 871.020 945.720 ;
        RECT 942.400 945.710 945.400 945.720 ;
        RECT -38.180 944.020 -35.180 944.030 ;
        RECT 58.020 944.020 61.020 944.030 ;
        RECT 238.020 944.020 241.020 944.030 ;
        RECT 418.020 944.020 421.020 944.030 ;
        RECT 598.020 944.020 601.020 944.030 ;
        RECT 778.020 944.020 781.020 944.030 ;
        RECT 937.700 944.020 940.700 944.030 ;
        RECT -38.180 941.010 -35.180 941.020 ;
        RECT 58.020 941.010 61.020 941.020 ;
        RECT 238.020 941.010 241.020 941.020 ;
        RECT 418.020 941.010 421.020 941.020 ;
        RECT 598.020 941.010 601.020 941.020 ;
        RECT 778.020 941.010 781.020 941.020 ;
        RECT 937.700 941.010 940.700 941.020 ;
        RECT -33.480 939.320 -30.480 939.330 ;
        RECT 130.020 939.320 133.020 939.330 ;
        RECT 310.020 939.320 313.020 939.330 ;
        RECT 490.020 939.320 493.020 939.330 ;
        RECT 670.020 939.320 673.020 939.330 ;
        RECT 850.020 939.320 853.020 939.330 ;
        RECT 933.000 939.320 936.000 939.330 ;
        RECT -33.480 936.310 -30.480 936.320 ;
        RECT 130.020 936.310 133.020 936.320 ;
        RECT 310.020 936.310 313.020 936.320 ;
        RECT 490.020 936.310 493.020 936.320 ;
        RECT 670.020 936.310 673.020 936.320 ;
        RECT 850.020 936.310 853.020 936.320 ;
        RECT 933.000 936.310 936.000 936.320 ;
        RECT -28.780 934.620 -25.780 934.630 ;
        RECT 40.020 934.620 43.020 934.630 ;
        RECT 220.020 934.620 223.020 934.630 ;
        RECT 400.020 934.620 403.020 934.630 ;
        RECT 580.020 934.620 583.020 934.630 ;
        RECT 760.020 934.620 763.020 934.630 ;
        RECT 928.300 934.620 931.300 934.630 ;
        RECT -28.780 931.610 -25.780 931.620 ;
        RECT 40.020 931.610 43.020 931.620 ;
        RECT 220.020 931.610 223.020 931.620 ;
        RECT 400.020 931.610 403.020 931.620 ;
        RECT 580.020 931.610 583.020 931.620 ;
        RECT 760.020 931.610 763.020 931.620 ;
        RECT 928.300 931.610 931.300 931.620 ;
        RECT -24.080 929.920 -21.080 929.930 ;
        RECT 112.020 929.920 115.020 929.930 ;
        RECT 292.020 929.920 295.020 929.930 ;
        RECT 472.020 929.920 475.020 929.930 ;
        RECT 652.020 929.920 655.020 929.930 ;
        RECT 832.020 929.920 835.020 929.930 ;
        RECT 923.600 929.920 926.600 929.930 ;
        RECT -24.080 926.910 -21.080 926.920 ;
        RECT 112.020 926.910 115.020 926.920 ;
        RECT 292.020 926.910 295.020 926.920 ;
        RECT 472.020 926.910 475.020 926.920 ;
        RECT 652.020 926.910 655.020 926.920 ;
        RECT 832.020 926.910 835.020 926.920 ;
        RECT 923.600 926.910 926.600 926.920 ;
        RECT -19.380 925.220 -16.380 925.230 ;
        RECT 22.020 925.220 25.020 925.230 ;
        RECT 202.020 925.220 205.020 925.230 ;
        RECT 382.020 925.220 385.020 925.230 ;
        RECT 562.020 925.220 565.020 925.230 ;
        RECT 742.020 925.220 745.020 925.230 ;
        RECT 918.900 925.220 921.900 925.230 ;
        RECT -19.380 922.210 -16.380 922.220 ;
        RECT 22.020 922.210 25.020 922.220 ;
        RECT 202.020 922.210 205.020 922.220 ;
        RECT 382.020 922.210 385.020 922.220 ;
        RECT 562.020 922.210 565.020 922.220 ;
        RECT 742.020 922.210 745.020 922.220 ;
        RECT 918.900 922.210 921.900 922.220 ;
        RECT -14.680 920.520 -11.680 920.530 ;
        RECT 94.020 920.520 97.020 920.530 ;
        RECT 274.020 920.520 277.020 920.530 ;
        RECT 454.020 920.520 457.020 920.530 ;
        RECT 634.020 920.520 637.020 920.530 ;
        RECT 814.020 920.520 817.020 920.530 ;
        RECT 914.200 920.520 917.200 920.530 ;
        RECT -14.680 917.510 -11.680 917.520 ;
        RECT 94.020 917.510 97.020 917.520 ;
        RECT 274.020 917.510 277.020 917.520 ;
        RECT 454.020 917.510 457.020 917.520 ;
        RECT 634.020 917.510 637.020 917.520 ;
        RECT 814.020 917.510 817.020 917.520 ;
        RECT 914.200 917.510 917.200 917.520 ;
        RECT -9.980 915.820 -6.980 915.830 ;
        RECT 4.020 915.820 7.020 915.830 ;
        RECT 184.020 915.820 187.020 915.830 ;
        RECT 364.020 915.820 367.020 915.830 ;
        RECT 544.020 915.820 547.020 915.830 ;
        RECT 724.020 915.820 727.020 915.830 ;
        RECT 909.500 915.820 912.500 915.830 ;
        RECT -9.980 912.810 -6.980 912.820 ;
        RECT 909.500 912.810 912.500 912.820 ;
        RECT 0.000 877.980 902.775 911.220 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 942.400 876.380 945.400 876.390 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 942.400 873.370 945.400 873.380 ;
        RECT 0.000 859.980 902.775 871.780 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 933.000 858.380 936.000 858.390 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 933.000 855.370 936.000 855.380 ;
        RECT 0.000 841.980 902.775 853.780 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 923.600 840.380 926.600 840.390 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 923.600 837.370 926.600 837.380 ;
        RECT 0.000 823.740 902.775 835.780 ;
        RECT -14.680 822.140 -11.680 822.150 ;
        RECT 914.200 822.140 917.200 822.150 ;
        RECT -14.680 819.130 -11.680 819.140 ;
        RECT 914.200 819.130 917.200 819.140 ;
        RECT 0.000 787.980 902.775 817.540 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 937.700 786.380 940.700 786.390 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 937.700 783.370 940.700 783.380 ;
        RECT 0.000 769.980 902.775 781.780 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 928.300 768.380 931.300 768.390 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 928.300 765.370 931.300 765.380 ;
        RECT 0.000 751.980 902.775 763.780 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 918.900 750.380 921.900 750.390 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 918.900 747.370 921.900 747.380 ;
        RECT 0.000 733.740 902.775 745.780 ;
        RECT -9.980 732.140 -6.980 732.150 ;
        RECT 909.500 732.140 912.500 732.150 ;
        RECT -9.980 729.130 -6.980 729.140 ;
        RECT 909.500 729.130 912.500 729.140 ;
        RECT 0.000 697.980 902.775 727.540 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 942.400 696.380 945.400 696.390 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 942.400 693.370 945.400 693.380 ;
        RECT 0.000 679.980 902.775 691.780 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 933.000 678.380 936.000 678.390 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 933.000 675.370 936.000 675.380 ;
        RECT 0.000 661.980 902.775 673.780 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 923.600 660.380 926.600 660.390 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 923.600 657.370 926.600 657.380 ;
        RECT 0.000 643.740 902.775 655.780 ;
        RECT -14.680 642.140 -11.680 642.150 ;
        RECT 914.200 642.140 917.200 642.150 ;
        RECT -14.680 639.130 -11.680 639.140 ;
        RECT 914.200 639.130 917.200 639.140 ;
        RECT 0.000 607.980 902.775 637.540 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 937.700 606.380 940.700 606.390 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 937.700 603.370 940.700 603.380 ;
        RECT 0.000 589.980 902.775 601.780 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 928.300 588.380 931.300 588.390 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 928.300 585.370 931.300 585.380 ;
        RECT 0.000 571.980 902.775 583.780 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 918.900 570.380 921.900 570.390 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 918.900 567.370 921.900 567.380 ;
        RECT 0.000 553.740 902.775 565.780 ;
        RECT -9.980 552.140 -6.980 552.150 ;
        RECT 909.500 552.140 912.500 552.150 ;
        RECT -9.980 549.130 -6.980 549.140 ;
        RECT 909.500 549.130 912.500 549.140 ;
        RECT 0.000 517.980 902.775 547.540 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 942.400 516.380 945.400 516.390 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 942.400 513.370 945.400 513.380 ;
        RECT 0.000 499.980 902.775 511.780 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 933.000 498.380 936.000 498.390 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 933.000 495.370 936.000 495.380 ;
        RECT 0.000 481.980 902.775 493.780 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 923.600 480.380 926.600 480.390 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 923.600 477.370 926.600 477.380 ;
        RECT 0.000 463.740 902.775 475.780 ;
        RECT -14.680 462.140 -11.680 462.150 ;
        RECT 914.200 462.140 917.200 462.150 ;
        RECT -14.680 459.130 -11.680 459.140 ;
        RECT 914.200 459.130 917.200 459.140 ;
        RECT 0.000 427.980 902.775 457.540 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 937.700 426.380 940.700 426.390 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 937.700 423.370 940.700 423.380 ;
        RECT 0.000 409.980 902.775 421.780 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 928.300 408.380 931.300 408.390 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 928.300 405.370 931.300 405.380 ;
        RECT 0.000 391.980 902.775 403.780 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 918.900 390.380 921.900 390.390 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 918.900 387.370 921.900 387.380 ;
        RECT 0.000 373.740 902.775 385.780 ;
        RECT -9.980 372.140 -6.980 372.150 ;
        RECT 909.500 372.140 912.500 372.150 ;
        RECT -9.980 369.130 -6.980 369.140 ;
        RECT 909.500 369.130 912.500 369.140 ;
        RECT 0.000 337.980 902.775 367.540 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 942.400 336.380 945.400 336.390 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 942.400 333.370 945.400 333.380 ;
        RECT 0.000 319.980 902.775 331.780 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 933.000 318.380 936.000 318.390 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 933.000 315.370 936.000 315.380 ;
        RECT 0.000 301.980 902.775 313.780 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 923.600 300.380 926.600 300.390 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 923.600 297.370 926.600 297.380 ;
        RECT 0.000 283.740 902.775 295.780 ;
        RECT -14.680 282.140 -11.680 282.150 ;
        RECT 914.200 282.140 917.200 282.150 ;
        RECT -14.680 279.130 -11.680 279.140 ;
        RECT 914.200 279.130 917.200 279.140 ;
        RECT 0.000 247.980 902.775 277.540 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 937.700 246.380 940.700 246.390 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 937.700 243.370 940.700 243.380 ;
        RECT 0.000 229.980 902.775 241.780 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 928.300 228.380 931.300 228.390 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 928.300 225.370 931.300 225.380 ;
        RECT 0.000 211.980 902.775 223.780 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 918.900 210.380 921.900 210.390 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 918.900 207.370 921.900 207.380 ;
        RECT 0.000 193.740 902.775 205.780 ;
        RECT -9.980 192.140 -6.980 192.150 ;
        RECT 909.500 192.140 912.500 192.150 ;
        RECT -9.980 189.130 -6.980 189.140 ;
        RECT 909.500 189.130 912.500 189.140 ;
        RECT 0.000 157.980 902.775 187.540 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 942.400 156.380 945.400 156.390 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 942.400 153.370 945.400 153.380 ;
        RECT 0.000 139.980 902.775 151.780 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 933.000 138.380 936.000 138.390 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 933.000 135.370 936.000 135.380 ;
        RECT 0.000 121.980 902.775 133.780 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 923.600 120.380 926.600 120.390 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 923.600 117.370 926.600 117.380 ;
        RECT 0.000 103.740 902.775 115.780 ;
        RECT -14.680 102.140 -11.680 102.150 ;
        RECT 914.200 102.140 917.200 102.150 ;
        RECT -14.680 99.130 -11.680 99.140 ;
        RECT 914.200 99.130 917.200 99.140 ;
        RECT 0.000 67.980 902.775 97.540 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 937.700 66.380 940.700 66.390 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 937.700 63.370 940.700 63.380 ;
        RECT 0.000 49.980 902.775 61.780 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 928.300 48.380 931.300 48.390 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 928.300 45.370 931.300 45.380 ;
        RECT 0.000 31.980 902.775 43.780 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 918.900 30.380 921.900 30.390 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 918.900 27.370 921.900 27.380 ;
        RECT 0.000 13.740 902.775 25.780 ;
        RECT -9.980 12.140 -6.980 12.150 ;
        RECT 909.500 12.140 912.500 12.150 ;
        RECT -9.980 9.130 -6.980 9.140 ;
        RECT 909.500 9.130 912.500 9.140 ;
        RECT 0.000 0.000 902.775 7.540 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 909.500 -1.620 912.500 -1.610 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 909.500 -4.630 912.500 -4.620 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 914.200 -6.320 917.200 -6.310 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 914.200 -9.330 917.200 -9.320 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 918.900 -11.020 921.900 -11.010 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 918.900 -14.030 921.900 -14.020 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 923.600 -15.720 926.600 -15.710 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 923.600 -18.730 926.600 -18.720 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 928.300 -20.420 931.300 -20.410 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 928.300 -23.430 931.300 -23.420 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 933.000 -25.120 936.000 -25.110 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 933.000 -28.130 936.000 -28.120 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 937.700 -29.820 940.700 -29.810 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 937.700 -32.830 940.700 -32.820 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 942.400 -34.520 945.400 -34.510 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 942.400 -37.530 945.400 -37.520 ;
  END
END user_project_wrapper
END LIBRARY

