magic
tech sky130A
magscale 1 2
timestamp 1622199858
<< obsli1 >>
rect 949 2261 179279 179843
<< obsm1 >>
rect 937 2128 179938 180112
<< metal2 >>
rect 938 181899 994 182699
rect 1858 181899 1914 182699
rect 2778 181899 2834 182699
rect 3698 181899 3754 182699
rect 4618 181899 4674 182699
rect 5538 181899 5594 182699
rect 6458 181899 6514 182699
rect 7838 181899 7894 182699
rect 8758 181899 8814 182699
rect 9678 181899 9734 182699
rect 10598 181899 10654 182699
rect 11518 181899 11574 182699
rect 12438 181899 12494 182699
rect 13358 181899 13414 182699
rect 14278 181899 14334 182699
rect 15198 181899 15254 182699
rect 16118 181899 16174 182699
rect 17038 181899 17094 182699
rect 17958 181899 18014 182699
rect 18878 181899 18934 182699
rect 19798 181899 19854 182699
rect 20718 181899 20774 182699
rect 22098 181899 22154 182699
rect 23018 181899 23074 182699
rect 23938 181899 23994 182699
rect 24858 181899 24914 182699
rect 25778 181899 25834 182699
rect 26698 181899 26754 182699
rect 27618 181899 27674 182699
rect 28538 181899 28594 182699
rect 29458 181899 29514 182699
rect 30378 181899 30434 182699
rect 31298 181899 31354 182699
rect 32218 181899 32274 182699
rect 33138 181899 33194 182699
rect 34058 181899 34114 182699
rect 34978 181899 35034 182699
rect 36358 181899 36414 182699
rect 37278 181899 37334 182699
rect 38198 181899 38254 182699
rect 39118 181899 39174 182699
rect 40038 181899 40094 182699
rect 40958 181899 41014 182699
rect 41878 181899 41934 182699
rect 42798 181899 42854 182699
rect 43718 181899 43774 182699
rect 44638 181899 44694 182699
rect 45558 181899 45614 182699
rect 46478 181899 46534 182699
rect 47398 181899 47454 182699
rect 48318 181899 48374 182699
rect 49238 181899 49294 182699
rect 50158 181899 50214 182699
rect 51538 181899 51594 182699
rect 52458 181899 52514 182699
rect 53378 181899 53434 182699
rect 54298 181899 54354 182699
rect 55218 181899 55274 182699
rect 56138 181899 56194 182699
rect 57058 181899 57114 182699
rect 57978 181899 58034 182699
rect 58898 181899 58954 182699
rect 59818 181899 59874 182699
rect 60738 181899 60794 182699
rect 61658 181899 61714 182699
rect 62578 181899 62634 182699
rect 63498 181899 63554 182699
rect 64418 181899 64474 182699
rect 65798 181899 65854 182699
rect 66718 181899 66774 182699
rect 67638 181899 67694 182699
rect 68558 181899 68614 182699
rect 69478 181899 69534 182699
rect 70398 181899 70454 182699
rect 71318 181899 71374 182699
rect 72238 181899 72294 182699
rect 73158 181899 73214 182699
rect 74078 181899 74134 182699
rect 74998 181899 75054 182699
rect 75918 181899 75974 182699
rect 76838 181899 76894 182699
rect 77758 181899 77814 182699
rect 78678 181899 78734 182699
rect 80058 181899 80114 182699
rect 80978 181899 81034 182699
rect 81898 181899 81954 182699
rect 82818 181899 82874 182699
rect 83738 181899 83794 182699
rect 84658 181899 84714 182699
rect 85578 181899 85634 182699
rect 86498 181899 86554 182699
rect 87418 181899 87474 182699
rect 88338 181899 88394 182699
rect 89258 181899 89314 182699
rect 90178 181899 90234 182699
rect 91098 181899 91154 182699
rect 92018 181899 92074 182699
rect 92938 181899 92994 182699
rect 94318 181899 94374 182699
rect 95238 181899 95294 182699
rect 96158 181899 96214 182699
rect 97078 181899 97134 182699
rect 97998 181899 98054 182699
rect 98918 181899 98974 182699
rect 99838 181899 99894 182699
rect 100758 181899 100814 182699
rect 101678 181899 101734 182699
rect 102598 181899 102654 182699
rect 103518 181899 103574 182699
rect 104438 181899 104494 182699
rect 105358 181899 105414 182699
rect 106278 181899 106334 182699
rect 107198 181899 107254 182699
rect 108578 181899 108634 182699
rect 109498 181899 109554 182699
rect 110418 181899 110474 182699
rect 111338 181899 111394 182699
rect 112258 181899 112314 182699
rect 113178 181899 113234 182699
rect 114098 181899 114154 182699
rect 115018 181899 115074 182699
rect 115938 181899 115994 182699
rect 116858 181899 116914 182699
rect 117778 181899 117834 182699
rect 118698 181899 118754 182699
rect 119618 181899 119674 182699
rect 120538 181899 120594 182699
rect 121458 181899 121514 182699
rect 122838 181899 122894 182699
rect 123758 181899 123814 182699
rect 124678 181899 124734 182699
rect 125598 181899 125654 182699
rect 126518 181899 126574 182699
rect 127438 181899 127494 182699
rect 128358 181899 128414 182699
rect 129278 181899 129334 182699
rect 130198 181899 130254 182699
rect 131118 181899 131174 182699
rect 132038 181899 132094 182699
rect 132958 181899 133014 182699
rect 133878 181899 133934 182699
rect 134798 181899 134854 182699
rect 135718 181899 135774 182699
rect 136638 181899 136694 182699
rect 138018 181899 138074 182699
rect 138938 181899 138994 182699
rect 139858 181899 139914 182699
rect 140778 181899 140834 182699
rect 141698 181899 141754 182699
rect 142618 181899 142674 182699
rect 143538 181899 143594 182699
rect 144458 181899 144514 182699
rect 145378 181899 145434 182699
rect 146298 181899 146354 182699
rect 147218 181899 147274 182699
rect 148138 181899 148194 182699
rect 149058 181899 149114 182699
rect 149978 181899 150034 182699
rect 150898 181899 150954 182699
rect 152278 181899 152334 182699
rect 153198 181899 153254 182699
rect 154118 181899 154174 182699
rect 155038 181899 155094 182699
rect 155958 181899 156014 182699
rect 156878 181899 156934 182699
rect 157798 181899 157854 182699
rect 158718 181899 158774 182699
rect 159638 181899 159694 182699
rect 160558 181899 160614 182699
rect 161478 181899 161534 182699
rect 162398 181899 162454 182699
rect 163318 181899 163374 182699
rect 164238 181899 164294 182699
rect 165158 181899 165214 182699
rect 166538 181899 166594 182699
rect 167458 181899 167514 182699
rect 168378 181899 168434 182699
rect 169298 181899 169354 182699
rect 170218 181899 170274 182699
rect 171138 181899 171194 182699
rect 172058 181899 172114 182699
rect 172978 181899 173034 182699
rect 173898 181899 173954 182699
rect 174818 181899 174874 182699
rect 175738 181899 175794 182699
rect 176658 181899 176714 182699
rect 177578 181899 177634 182699
rect 178498 181899 178554 182699
rect 179418 181899 179474 182699
rect 478 0 534 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 3238 0 3294 800
rect 4158 0 4214 800
rect 5078 0 5134 800
rect 5998 0 6054 800
rect 6918 0 6974 800
rect 7838 0 7894 800
rect 8758 0 8814 800
rect 9678 0 9734 800
rect 10598 0 10654 800
rect 11518 0 11574 800
rect 12438 0 12494 800
rect 13358 0 13414 800
rect 14278 0 14334 800
rect 15658 0 15714 800
rect 16578 0 16634 800
rect 17498 0 17554 800
rect 18418 0 18474 800
rect 19338 0 19394 800
rect 20258 0 20314 800
rect 21178 0 21234 800
rect 22098 0 22154 800
rect 23018 0 23074 800
rect 23938 0 23994 800
rect 24858 0 24914 800
rect 25778 0 25834 800
rect 26698 0 26754 800
rect 27618 0 27674 800
rect 28538 0 28594 800
rect 29918 0 29974 800
rect 30838 0 30894 800
rect 31758 0 31814 800
rect 32678 0 32734 800
rect 33598 0 33654 800
rect 34518 0 34574 800
rect 35438 0 35494 800
rect 36358 0 36414 800
rect 37278 0 37334 800
rect 38198 0 38254 800
rect 39118 0 39174 800
rect 40038 0 40094 800
rect 40958 0 41014 800
rect 41878 0 41934 800
rect 42798 0 42854 800
rect 44178 0 44234 800
rect 45098 0 45154 800
rect 46018 0 46074 800
rect 46938 0 46994 800
rect 47858 0 47914 800
rect 48778 0 48834 800
rect 49698 0 49754 800
rect 50618 0 50674 800
rect 51538 0 51594 800
rect 52458 0 52514 800
rect 53378 0 53434 800
rect 54298 0 54354 800
rect 55218 0 55274 800
rect 56138 0 56194 800
rect 57058 0 57114 800
rect 58438 0 58494 800
rect 59358 0 59414 800
rect 60278 0 60334 800
rect 61198 0 61254 800
rect 62118 0 62174 800
rect 63038 0 63094 800
rect 63958 0 64014 800
rect 64878 0 64934 800
rect 65798 0 65854 800
rect 66718 0 66774 800
rect 67638 0 67694 800
rect 68558 0 68614 800
rect 69478 0 69534 800
rect 70398 0 70454 800
rect 71318 0 71374 800
rect 72698 0 72754 800
rect 73618 0 73674 800
rect 74538 0 74594 800
rect 75458 0 75514 800
rect 76378 0 76434 800
rect 77298 0 77354 800
rect 78218 0 78274 800
rect 79138 0 79194 800
rect 80058 0 80114 800
rect 80978 0 81034 800
rect 81898 0 81954 800
rect 82818 0 82874 800
rect 83738 0 83794 800
rect 84658 0 84714 800
rect 85578 0 85634 800
rect 86958 0 87014 800
rect 87878 0 87934 800
rect 88798 0 88854 800
rect 89718 0 89774 800
rect 90638 0 90694 800
rect 91558 0 91614 800
rect 92478 0 92534 800
rect 93398 0 93454 800
rect 94318 0 94374 800
rect 95238 0 95294 800
rect 96158 0 96214 800
rect 97078 0 97134 800
rect 97998 0 98054 800
rect 98918 0 98974 800
rect 99838 0 99894 800
rect 100758 0 100814 800
rect 102138 0 102194 800
rect 103058 0 103114 800
rect 103978 0 104034 800
rect 104898 0 104954 800
rect 105818 0 105874 800
rect 106738 0 106794 800
rect 107658 0 107714 800
rect 108578 0 108634 800
rect 109498 0 109554 800
rect 110418 0 110474 800
rect 111338 0 111394 800
rect 112258 0 112314 800
rect 113178 0 113234 800
rect 114098 0 114154 800
rect 115018 0 115074 800
rect 116398 0 116454 800
rect 117318 0 117374 800
rect 118238 0 118294 800
rect 119158 0 119214 800
rect 120078 0 120134 800
rect 120998 0 121054 800
rect 121918 0 121974 800
rect 122838 0 122894 800
rect 123758 0 123814 800
rect 124678 0 124734 800
rect 125598 0 125654 800
rect 126518 0 126574 800
rect 127438 0 127494 800
rect 128358 0 128414 800
rect 129278 0 129334 800
rect 130658 0 130714 800
rect 131578 0 131634 800
rect 132498 0 132554 800
rect 133418 0 133474 800
rect 134338 0 134394 800
rect 135258 0 135314 800
rect 136178 0 136234 800
rect 137098 0 137154 800
rect 138018 0 138074 800
rect 138938 0 138994 800
rect 139858 0 139914 800
rect 140778 0 140834 800
rect 141698 0 141754 800
rect 142618 0 142674 800
rect 143538 0 143594 800
rect 144918 0 144974 800
rect 145838 0 145894 800
rect 146758 0 146814 800
rect 147678 0 147734 800
rect 148598 0 148654 800
rect 149518 0 149574 800
rect 150438 0 150494 800
rect 151358 0 151414 800
rect 152278 0 152334 800
rect 153198 0 153254 800
rect 154118 0 154174 800
rect 155038 0 155094 800
rect 155958 0 156014 800
rect 156878 0 156934 800
rect 157798 0 157854 800
rect 159178 0 159234 800
rect 160098 0 160154 800
rect 161018 0 161074 800
rect 161938 0 161994 800
rect 162858 0 162914 800
rect 163778 0 163834 800
rect 164698 0 164754 800
rect 165618 0 165674 800
rect 166538 0 166594 800
rect 167458 0 167514 800
rect 168378 0 168434 800
rect 169298 0 169354 800
rect 170218 0 170274 800
rect 171138 0 171194 800
rect 172058 0 172114 800
rect 173438 0 173494 800
rect 174358 0 174414 800
rect 175278 0 175334 800
rect 176198 0 176254 800
rect 177118 0 177174 800
rect 178038 0 178094 800
rect 178958 0 179014 800
rect 179878 0 179934 800
<< obsm2 >>
rect 1216 181843 1802 181899
rect 1970 181843 2722 181899
rect 2890 181843 3642 181899
rect 3810 181843 4562 181899
rect 4730 181843 5482 181899
rect 5650 181843 6402 181899
rect 6570 181843 7782 181899
rect 7950 181843 8702 181899
rect 8870 181843 9622 181899
rect 9790 181843 10542 181899
rect 10710 181843 11462 181899
rect 11630 181843 12382 181899
rect 12550 181843 13302 181899
rect 13470 181843 14222 181899
rect 14390 181843 15142 181899
rect 15310 181843 16062 181899
rect 16230 181843 16982 181899
rect 17150 181843 17902 181899
rect 18070 181843 18822 181899
rect 18990 181843 19742 181899
rect 19910 181843 20662 181899
rect 20830 181843 22042 181899
rect 22210 181843 22962 181899
rect 23130 181843 23882 181899
rect 24050 181843 24802 181899
rect 24970 181843 25722 181899
rect 25890 181843 26642 181899
rect 26810 181843 27562 181899
rect 27730 181843 28482 181899
rect 28650 181843 29402 181899
rect 29570 181843 30322 181899
rect 30490 181843 31242 181899
rect 31410 181843 32162 181899
rect 32330 181843 33082 181899
rect 33250 181843 34002 181899
rect 34170 181843 34922 181899
rect 35090 181843 36302 181899
rect 36470 181843 37222 181899
rect 37390 181843 38142 181899
rect 38310 181843 39062 181899
rect 39230 181843 39982 181899
rect 40150 181843 40902 181899
rect 41070 181843 41822 181899
rect 41990 181843 42742 181899
rect 42910 181843 43662 181899
rect 43830 181843 44582 181899
rect 44750 181843 45502 181899
rect 45670 181843 46422 181899
rect 46590 181843 47342 181899
rect 47510 181843 48262 181899
rect 48430 181843 49182 181899
rect 49350 181843 50102 181899
rect 50270 181843 51482 181899
rect 51650 181843 52402 181899
rect 52570 181843 53322 181899
rect 53490 181843 54242 181899
rect 54410 181843 55162 181899
rect 55330 181843 56082 181899
rect 56250 181843 57002 181899
rect 57170 181843 57922 181899
rect 58090 181843 58842 181899
rect 59010 181843 59762 181899
rect 59930 181843 60682 181899
rect 60850 181843 61602 181899
rect 61770 181843 62522 181899
rect 62690 181843 63442 181899
rect 63610 181843 64362 181899
rect 64530 181843 65742 181899
rect 65910 181843 66662 181899
rect 66830 181843 67582 181899
rect 67750 181843 68502 181899
rect 68670 181843 69422 181899
rect 69590 181843 70342 181899
rect 70510 181843 71262 181899
rect 71430 181843 72182 181899
rect 72350 181843 73102 181899
rect 73270 181843 74022 181899
rect 74190 181843 74942 181899
rect 75110 181843 75862 181899
rect 76030 181843 76782 181899
rect 76950 181843 77702 181899
rect 77870 181843 78622 181899
rect 78790 181843 80002 181899
rect 80170 181843 80922 181899
rect 81090 181843 81842 181899
rect 82010 181843 82762 181899
rect 82930 181843 83682 181899
rect 83850 181843 84602 181899
rect 84770 181843 85522 181899
rect 85690 181843 86442 181899
rect 86610 181843 87362 181899
rect 87530 181843 88282 181899
rect 88450 181843 89202 181899
rect 89370 181843 90122 181899
rect 90290 181843 91042 181899
rect 91210 181843 91962 181899
rect 92130 181843 92882 181899
rect 93050 181843 94262 181899
rect 94430 181843 95182 181899
rect 95350 181843 96102 181899
rect 96270 181843 97022 181899
rect 97190 181843 97942 181899
rect 98110 181843 98862 181899
rect 99030 181843 99782 181899
rect 99950 181843 100702 181899
rect 100870 181843 101622 181899
rect 101790 181843 102542 181899
rect 102710 181843 103462 181899
rect 103630 181843 104382 181899
rect 104550 181843 105302 181899
rect 105470 181843 106222 181899
rect 106390 181843 107142 181899
rect 107310 181843 108522 181899
rect 108690 181843 109442 181899
rect 109610 181843 110362 181899
rect 110530 181843 111282 181899
rect 111450 181843 112202 181899
rect 112370 181843 113122 181899
rect 113290 181843 114042 181899
rect 114210 181843 114962 181899
rect 115130 181843 115882 181899
rect 116050 181843 116802 181899
rect 116970 181843 117722 181899
rect 117890 181843 118642 181899
rect 118810 181843 119562 181899
rect 119730 181843 120482 181899
rect 120650 181843 121402 181899
rect 121570 181843 122782 181899
rect 122950 181843 123702 181899
rect 123870 181843 124622 181899
rect 124790 181843 125542 181899
rect 125710 181843 126462 181899
rect 126630 181843 127382 181899
rect 127550 181843 128302 181899
rect 128470 181843 129222 181899
rect 129390 181843 130142 181899
rect 130310 181843 131062 181899
rect 131230 181843 131982 181899
rect 132150 181843 132902 181899
rect 133070 181843 133822 181899
rect 133990 181843 134742 181899
rect 134910 181843 135662 181899
rect 135830 181843 136582 181899
rect 136750 181843 137962 181899
rect 138130 181843 138882 181899
rect 139050 181843 139802 181899
rect 139970 181843 140722 181899
rect 140890 181843 141642 181899
rect 141810 181843 142562 181899
rect 142730 181843 143482 181899
rect 143650 181843 144402 181899
rect 144570 181843 145322 181899
rect 145490 181843 146242 181899
rect 146410 181843 147162 181899
rect 147330 181843 148082 181899
rect 148250 181843 149002 181899
rect 149170 181843 149922 181899
rect 150090 181843 150842 181899
rect 151010 181843 152222 181899
rect 152390 181843 153142 181899
rect 153310 181843 154062 181899
rect 154230 181843 154982 181899
rect 155150 181843 155902 181899
rect 156070 181843 156822 181899
rect 156990 181843 157742 181899
rect 157910 181843 158662 181899
rect 158830 181843 159582 181899
rect 159750 181843 160502 181899
rect 160670 181843 161422 181899
rect 161590 181843 162342 181899
rect 162510 181843 163262 181899
rect 163430 181843 164182 181899
rect 164350 181843 165102 181899
rect 165270 181843 166482 181899
rect 166650 181843 167402 181899
rect 167570 181843 168322 181899
rect 168490 181843 169242 181899
rect 169410 181843 170162 181899
rect 170330 181843 171082 181899
rect 171250 181843 172002 181899
rect 172170 181843 172922 181899
rect 173090 181843 173842 181899
rect 174010 181843 174762 181899
rect 174930 181843 175682 181899
rect 175850 181843 176602 181899
rect 176770 181843 177522 181899
rect 177690 181843 178442 181899
rect 178610 181843 179362 181899
rect 179530 181843 179932 181899
rect 1216 856 179932 181843
rect 1216 800 1342 856
rect 1510 800 2262 856
rect 2430 800 3182 856
rect 3350 800 4102 856
rect 4270 800 5022 856
rect 5190 800 5942 856
rect 6110 800 6862 856
rect 7030 800 7782 856
rect 7950 800 8702 856
rect 8870 800 9622 856
rect 9790 800 10542 856
rect 10710 800 11462 856
rect 11630 800 12382 856
rect 12550 800 13302 856
rect 13470 800 14222 856
rect 14390 800 15602 856
rect 15770 800 16522 856
rect 16690 800 17442 856
rect 17610 800 18362 856
rect 18530 800 19282 856
rect 19450 800 20202 856
rect 20370 800 21122 856
rect 21290 800 22042 856
rect 22210 800 22962 856
rect 23130 800 23882 856
rect 24050 800 24802 856
rect 24970 800 25722 856
rect 25890 800 26642 856
rect 26810 800 27562 856
rect 27730 800 28482 856
rect 28650 800 29862 856
rect 30030 800 30782 856
rect 30950 800 31702 856
rect 31870 800 32622 856
rect 32790 800 33542 856
rect 33710 800 34462 856
rect 34630 800 35382 856
rect 35550 800 36302 856
rect 36470 800 37222 856
rect 37390 800 38142 856
rect 38310 800 39062 856
rect 39230 800 39982 856
rect 40150 800 40902 856
rect 41070 800 41822 856
rect 41990 800 42742 856
rect 42910 800 44122 856
rect 44290 800 45042 856
rect 45210 800 45962 856
rect 46130 800 46882 856
rect 47050 800 47802 856
rect 47970 800 48722 856
rect 48890 800 49642 856
rect 49810 800 50562 856
rect 50730 800 51482 856
rect 51650 800 52402 856
rect 52570 800 53322 856
rect 53490 800 54242 856
rect 54410 800 55162 856
rect 55330 800 56082 856
rect 56250 800 57002 856
rect 57170 800 58382 856
rect 58550 800 59302 856
rect 59470 800 60222 856
rect 60390 800 61142 856
rect 61310 800 62062 856
rect 62230 800 62982 856
rect 63150 800 63902 856
rect 64070 800 64822 856
rect 64990 800 65742 856
rect 65910 800 66662 856
rect 66830 800 67582 856
rect 67750 800 68502 856
rect 68670 800 69422 856
rect 69590 800 70342 856
rect 70510 800 71262 856
rect 71430 800 72642 856
rect 72810 800 73562 856
rect 73730 800 74482 856
rect 74650 800 75402 856
rect 75570 800 76322 856
rect 76490 800 77242 856
rect 77410 800 78162 856
rect 78330 800 79082 856
rect 79250 800 80002 856
rect 80170 800 80922 856
rect 81090 800 81842 856
rect 82010 800 82762 856
rect 82930 800 83682 856
rect 83850 800 84602 856
rect 84770 800 85522 856
rect 85690 800 86902 856
rect 87070 800 87822 856
rect 87990 800 88742 856
rect 88910 800 89662 856
rect 89830 800 90582 856
rect 90750 800 91502 856
rect 91670 800 92422 856
rect 92590 800 93342 856
rect 93510 800 94262 856
rect 94430 800 95182 856
rect 95350 800 96102 856
rect 96270 800 97022 856
rect 97190 800 97942 856
rect 98110 800 98862 856
rect 99030 800 99782 856
rect 99950 800 100702 856
rect 100870 800 102082 856
rect 102250 800 103002 856
rect 103170 800 103922 856
rect 104090 800 104842 856
rect 105010 800 105762 856
rect 105930 800 106682 856
rect 106850 800 107602 856
rect 107770 800 108522 856
rect 108690 800 109442 856
rect 109610 800 110362 856
rect 110530 800 111282 856
rect 111450 800 112202 856
rect 112370 800 113122 856
rect 113290 800 114042 856
rect 114210 800 114962 856
rect 115130 800 116342 856
rect 116510 800 117262 856
rect 117430 800 118182 856
rect 118350 800 119102 856
rect 119270 800 120022 856
rect 120190 800 120942 856
rect 121110 800 121862 856
rect 122030 800 122782 856
rect 122950 800 123702 856
rect 123870 800 124622 856
rect 124790 800 125542 856
rect 125710 800 126462 856
rect 126630 800 127382 856
rect 127550 800 128302 856
rect 128470 800 129222 856
rect 129390 800 130602 856
rect 130770 800 131522 856
rect 131690 800 132442 856
rect 132610 800 133362 856
rect 133530 800 134282 856
rect 134450 800 135202 856
rect 135370 800 136122 856
rect 136290 800 137042 856
rect 137210 800 137962 856
rect 138130 800 138882 856
rect 139050 800 139802 856
rect 139970 800 140722 856
rect 140890 800 141642 856
rect 141810 800 142562 856
rect 142730 800 143482 856
rect 143650 800 144862 856
rect 145030 800 145782 856
rect 145950 800 146702 856
rect 146870 800 147622 856
rect 147790 800 148542 856
rect 148710 800 149462 856
rect 149630 800 150382 856
rect 150550 800 151302 856
rect 151470 800 152222 856
rect 152390 800 153142 856
rect 153310 800 154062 856
rect 154230 800 154982 856
rect 155150 800 155902 856
rect 156070 800 156822 856
rect 156990 800 157742 856
rect 157910 800 159122 856
rect 159290 800 160042 856
rect 160210 800 160962 856
rect 161130 800 161882 856
rect 162050 800 162802 856
rect 162970 800 163722 856
rect 163890 800 164642 856
rect 164810 800 165562 856
rect 165730 800 166482 856
rect 166650 800 167402 856
rect 167570 800 168322 856
rect 168490 800 169242 856
rect 169410 800 170162 856
rect 170330 800 171082 856
rect 171250 800 172002 856
rect 172170 800 173382 856
rect 173550 800 174302 856
rect 174470 800 175222 856
rect 175390 800 176142 856
rect 176310 800 177062 856
rect 177230 800 177982 856
rect 178150 800 178902 856
rect 179070 800 179822 856
<< metal3 >>
rect 0 181568 800 181688
rect 179755 180888 180555 181008
rect 0 180208 800 180328
rect 179755 179528 180555 179648
rect 0 178848 800 178968
rect 179755 178168 180555 178288
rect 0 177488 800 177608
rect 179755 176808 180555 176928
rect 0 176128 800 176248
rect 179755 175448 180555 175568
rect 0 174768 800 174888
rect 179755 174088 180555 174208
rect 0 173408 800 173528
rect 179755 172728 180555 172848
rect 0 172048 800 172168
rect 179755 171368 180555 171488
rect 0 170008 800 170128
rect 179755 170008 180555 170128
rect 0 168648 800 168768
rect 179755 168648 180555 168768
rect 0 167288 800 167408
rect 179755 167288 180555 167408
rect 0 165928 800 166048
rect 179755 165928 180555 166048
rect 0 164568 800 164688
rect 179755 164568 180555 164688
rect 0 163208 800 163328
rect 179755 163208 180555 163328
rect 0 161848 800 161968
rect 179755 161848 180555 161968
rect 0 160488 800 160608
rect 179755 159808 180555 159928
rect 0 159128 800 159248
rect 179755 158448 180555 158568
rect 0 157768 800 157888
rect 179755 157088 180555 157208
rect 0 156408 800 156528
rect 179755 155728 180555 155848
rect 0 155048 800 155168
rect 179755 154368 180555 154488
rect 0 153688 800 153808
rect 179755 153008 180555 153128
rect 0 152328 800 152448
rect 179755 151648 180555 151768
rect 0 150968 800 151088
rect 179755 150288 180555 150408
rect 0 148928 800 149048
rect 179755 148928 180555 149048
rect 0 147568 800 147688
rect 179755 147568 180555 147688
rect 0 146208 800 146328
rect 179755 146208 180555 146328
rect 0 144848 800 144968
rect 179755 144848 180555 144968
rect 0 143488 800 143608
rect 179755 143488 180555 143608
rect 0 142128 800 142248
rect 179755 142128 180555 142248
rect 0 140768 800 140888
rect 179755 140768 180555 140888
rect 0 139408 800 139528
rect 179755 138728 180555 138848
rect 0 138048 800 138168
rect 179755 137368 180555 137488
rect 0 136688 800 136808
rect 179755 136008 180555 136128
rect 0 135328 800 135448
rect 179755 134648 180555 134768
rect 0 133968 800 134088
rect 179755 133288 180555 133408
rect 0 132608 800 132728
rect 179755 131928 180555 132048
rect 0 131248 800 131368
rect 179755 130568 180555 130688
rect 0 129888 800 130008
rect 179755 129208 180555 129328
rect 0 127848 800 127968
rect 179755 127848 180555 127968
rect 0 126488 800 126608
rect 179755 126488 180555 126608
rect 0 125128 800 125248
rect 179755 125128 180555 125248
rect 0 123768 800 123888
rect 179755 123768 180555 123888
rect 0 122408 800 122528
rect 179755 122408 180555 122528
rect 0 121048 800 121168
rect 179755 121048 180555 121168
rect 0 119688 800 119808
rect 179755 119688 180555 119808
rect 0 118328 800 118448
rect 179755 118328 180555 118448
rect 0 116968 800 117088
rect 179755 116288 180555 116408
rect 0 115608 800 115728
rect 179755 114928 180555 115048
rect 0 114248 800 114368
rect 179755 113568 180555 113688
rect 0 112888 800 113008
rect 179755 112208 180555 112328
rect 0 111528 800 111648
rect 179755 110848 180555 110968
rect 0 110168 800 110288
rect 179755 109488 180555 109608
rect 0 108808 800 108928
rect 179755 108128 180555 108248
rect 0 107448 800 107568
rect 179755 106768 180555 106888
rect 0 105408 800 105528
rect 179755 105408 180555 105528
rect 0 104048 800 104168
rect 179755 104048 180555 104168
rect 0 102688 800 102808
rect 179755 102688 180555 102808
rect 0 101328 800 101448
rect 179755 101328 180555 101448
rect 0 99968 800 100088
rect 179755 99968 180555 100088
rect 0 98608 800 98728
rect 179755 98608 180555 98728
rect 0 97248 800 97368
rect 179755 97248 180555 97368
rect 0 95888 800 96008
rect 179755 95208 180555 95328
rect 0 94528 800 94648
rect 179755 93848 180555 93968
rect 0 93168 800 93288
rect 179755 92488 180555 92608
rect 0 91808 800 91928
rect 179755 91128 180555 91248
rect 0 90448 800 90568
rect 179755 89768 180555 89888
rect 0 89088 800 89208
rect 179755 88408 180555 88528
rect 0 87728 800 87848
rect 179755 87048 180555 87168
rect 0 86368 800 86488
rect 179755 85688 180555 85808
rect 0 84328 800 84448
rect 179755 84328 180555 84448
rect 0 82968 800 83088
rect 179755 82968 180555 83088
rect 0 81608 800 81728
rect 179755 81608 180555 81728
rect 0 80248 800 80368
rect 179755 80248 180555 80368
rect 0 78888 800 79008
rect 179755 78888 180555 79008
rect 0 77528 800 77648
rect 179755 77528 180555 77648
rect 0 76168 800 76288
rect 179755 76168 180555 76288
rect 0 74808 800 74928
rect 179755 74128 180555 74248
rect 0 73448 800 73568
rect 179755 72768 180555 72888
rect 0 72088 800 72208
rect 179755 71408 180555 71528
rect 0 70728 800 70848
rect 179755 70048 180555 70168
rect 0 69368 800 69488
rect 179755 68688 180555 68808
rect 0 68008 800 68128
rect 179755 67328 180555 67448
rect 0 66648 800 66768
rect 179755 65968 180555 66088
rect 0 65288 800 65408
rect 179755 64608 180555 64728
rect 0 63248 800 63368
rect 179755 63248 180555 63368
rect 0 61888 800 62008
rect 179755 61888 180555 62008
rect 0 60528 800 60648
rect 179755 60528 180555 60648
rect 0 59168 800 59288
rect 179755 59168 180555 59288
rect 0 57808 800 57928
rect 179755 57808 180555 57928
rect 0 56448 800 56568
rect 179755 56448 180555 56568
rect 0 55088 800 55208
rect 179755 55088 180555 55208
rect 0 53728 800 53848
rect 179755 53048 180555 53168
rect 0 52368 800 52488
rect 179755 51688 180555 51808
rect 0 51008 800 51128
rect 179755 50328 180555 50448
rect 0 49648 800 49768
rect 179755 48968 180555 49088
rect 0 48288 800 48408
rect 179755 47608 180555 47728
rect 0 46928 800 47048
rect 179755 46248 180555 46368
rect 0 45568 800 45688
rect 179755 44888 180555 45008
rect 0 44208 800 44328
rect 179755 43528 180555 43648
rect 0 42168 800 42288
rect 179755 42168 180555 42288
rect 0 40808 800 40928
rect 179755 40808 180555 40928
rect 0 39448 800 39568
rect 179755 39448 180555 39568
rect 0 38088 800 38208
rect 179755 38088 180555 38208
rect 0 36728 800 36848
rect 179755 36728 180555 36848
rect 0 35368 800 35488
rect 179755 35368 180555 35488
rect 0 34008 800 34128
rect 179755 34008 180555 34128
rect 0 32648 800 32768
rect 179755 31968 180555 32088
rect 0 31288 800 31408
rect 179755 30608 180555 30728
rect 0 29928 800 30048
rect 179755 29248 180555 29368
rect 0 28568 800 28688
rect 179755 27888 180555 28008
rect 0 27208 800 27328
rect 179755 26528 180555 26648
rect 0 25848 800 25968
rect 179755 25168 180555 25288
rect 0 24488 800 24608
rect 179755 23808 180555 23928
rect 0 23128 800 23248
rect 179755 22448 180555 22568
rect 0 21088 800 21208
rect 179755 21088 180555 21208
rect 0 19728 800 19848
rect 179755 19728 180555 19848
rect 0 18368 800 18488
rect 179755 18368 180555 18488
rect 0 17008 800 17128
rect 179755 17008 180555 17128
rect 0 15648 800 15768
rect 179755 15648 180555 15768
rect 0 14288 800 14408
rect 179755 14288 180555 14408
rect 0 12928 800 13048
rect 179755 12928 180555 13048
rect 0 11568 800 11688
rect 179755 10888 180555 11008
rect 0 10208 800 10328
rect 179755 9528 180555 9648
rect 0 8848 800 8968
rect 179755 8168 180555 8288
rect 0 7488 800 7608
rect 179755 6808 180555 6928
rect 0 6128 800 6248
rect 179755 5448 180555 5568
rect 0 4768 800 4888
rect 179755 4088 180555 4208
rect 0 3408 800 3528
rect 179755 2728 180555 2848
rect 0 2048 800 2168
rect 179755 1368 180555 1488
<< obsm3 >>
rect 800 180808 179675 180981
rect 800 180408 179755 180808
rect 880 180128 179755 180408
rect 800 179728 179755 180128
rect 800 179448 179675 179728
rect 800 179048 179755 179448
rect 880 178768 179755 179048
rect 800 178368 179755 178768
rect 800 178088 179675 178368
rect 800 177688 179755 178088
rect 880 177408 179755 177688
rect 800 177008 179755 177408
rect 800 176728 179675 177008
rect 800 176328 179755 176728
rect 880 176048 179755 176328
rect 800 175648 179755 176048
rect 800 175368 179675 175648
rect 800 174968 179755 175368
rect 880 174688 179755 174968
rect 800 174288 179755 174688
rect 800 174008 179675 174288
rect 800 173608 179755 174008
rect 880 173328 179755 173608
rect 800 172928 179755 173328
rect 800 172648 179675 172928
rect 800 172248 179755 172648
rect 880 171968 179755 172248
rect 800 171568 179755 171968
rect 800 171288 179675 171568
rect 800 170208 179755 171288
rect 880 169928 179675 170208
rect 800 168848 179755 169928
rect 880 168568 179675 168848
rect 800 167488 179755 168568
rect 880 167208 179675 167488
rect 800 166128 179755 167208
rect 880 165848 179675 166128
rect 800 164768 179755 165848
rect 880 164488 179675 164768
rect 800 163408 179755 164488
rect 880 163128 179675 163408
rect 800 162048 179755 163128
rect 880 161768 179675 162048
rect 800 160688 179755 161768
rect 880 160408 179755 160688
rect 800 160008 179755 160408
rect 800 159728 179675 160008
rect 800 159328 179755 159728
rect 880 159048 179755 159328
rect 800 158648 179755 159048
rect 800 158368 179675 158648
rect 800 157968 179755 158368
rect 880 157688 179755 157968
rect 800 157288 179755 157688
rect 800 157008 179675 157288
rect 800 156608 179755 157008
rect 880 156328 179755 156608
rect 800 155928 179755 156328
rect 800 155648 179675 155928
rect 800 155248 179755 155648
rect 880 154968 179755 155248
rect 800 154568 179755 154968
rect 800 154288 179675 154568
rect 800 153888 179755 154288
rect 880 153608 179755 153888
rect 800 153208 179755 153608
rect 800 152928 179675 153208
rect 800 152528 179755 152928
rect 880 152248 179755 152528
rect 800 151848 179755 152248
rect 800 151568 179675 151848
rect 800 151168 179755 151568
rect 880 150888 179755 151168
rect 800 150488 179755 150888
rect 800 150208 179675 150488
rect 800 149128 179755 150208
rect 880 148848 179675 149128
rect 800 147768 179755 148848
rect 880 147488 179675 147768
rect 800 146408 179755 147488
rect 880 146128 179675 146408
rect 800 145048 179755 146128
rect 880 144768 179675 145048
rect 800 143688 179755 144768
rect 880 143408 179675 143688
rect 800 142328 179755 143408
rect 880 142048 179675 142328
rect 800 140968 179755 142048
rect 880 140688 179675 140968
rect 800 139608 179755 140688
rect 880 139328 179755 139608
rect 800 138928 179755 139328
rect 800 138648 179675 138928
rect 800 138248 179755 138648
rect 880 137968 179755 138248
rect 800 137568 179755 137968
rect 800 137288 179675 137568
rect 800 136888 179755 137288
rect 880 136608 179755 136888
rect 800 136208 179755 136608
rect 800 135928 179675 136208
rect 800 135528 179755 135928
rect 880 135248 179755 135528
rect 800 134848 179755 135248
rect 800 134568 179675 134848
rect 800 134168 179755 134568
rect 880 133888 179755 134168
rect 800 133488 179755 133888
rect 800 133208 179675 133488
rect 800 132808 179755 133208
rect 880 132528 179755 132808
rect 800 132128 179755 132528
rect 800 131848 179675 132128
rect 800 131448 179755 131848
rect 880 131168 179755 131448
rect 800 130768 179755 131168
rect 800 130488 179675 130768
rect 800 130088 179755 130488
rect 880 129808 179755 130088
rect 800 129408 179755 129808
rect 800 129128 179675 129408
rect 800 128048 179755 129128
rect 880 127768 179675 128048
rect 800 126688 179755 127768
rect 880 126408 179675 126688
rect 800 125328 179755 126408
rect 880 125048 179675 125328
rect 800 123968 179755 125048
rect 880 123688 179675 123968
rect 800 122608 179755 123688
rect 880 122328 179675 122608
rect 800 121248 179755 122328
rect 880 120968 179675 121248
rect 800 119888 179755 120968
rect 880 119608 179675 119888
rect 800 118528 179755 119608
rect 880 118248 179675 118528
rect 800 117168 179755 118248
rect 880 116888 179755 117168
rect 800 116488 179755 116888
rect 800 116208 179675 116488
rect 800 115808 179755 116208
rect 880 115528 179755 115808
rect 800 115128 179755 115528
rect 800 114848 179675 115128
rect 800 114448 179755 114848
rect 880 114168 179755 114448
rect 800 113768 179755 114168
rect 800 113488 179675 113768
rect 800 113088 179755 113488
rect 880 112808 179755 113088
rect 800 112408 179755 112808
rect 800 112128 179675 112408
rect 800 111728 179755 112128
rect 880 111448 179755 111728
rect 800 111048 179755 111448
rect 800 110768 179675 111048
rect 800 110368 179755 110768
rect 880 110088 179755 110368
rect 800 109688 179755 110088
rect 800 109408 179675 109688
rect 800 109008 179755 109408
rect 880 108728 179755 109008
rect 800 108328 179755 108728
rect 800 108048 179675 108328
rect 800 107648 179755 108048
rect 880 107368 179755 107648
rect 800 106968 179755 107368
rect 800 106688 179675 106968
rect 800 105608 179755 106688
rect 880 105328 179675 105608
rect 800 104248 179755 105328
rect 880 103968 179675 104248
rect 800 102888 179755 103968
rect 880 102608 179675 102888
rect 800 101528 179755 102608
rect 880 101248 179675 101528
rect 800 100168 179755 101248
rect 880 99888 179675 100168
rect 800 98808 179755 99888
rect 880 98528 179675 98808
rect 800 97448 179755 98528
rect 880 97168 179675 97448
rect 800 96088 179755 97168
rect 880 95808 179755 96088
rect 800 95408 179755 95808
rect 800 95128 179675 95408
rect 800 94728 179755 95128
rect 880 94448 179755 94728
rect 800 94048 179755 94448
rect 800 93768 179675 94048
rect 800 93368 179755 93768
rect 880 93088 179755 93368
rect 800 92688 179755 93088
rect 800 92408 179675 92688
rect 800 92008 179755 92408
rect 880 91728 179755 92008
rect 800 91328 179755 91728
rect 800 91048 179675 91328
rect 800 90648 179755 91048
rect 880 90368 179755 90648
rect 800 89968 179755 90368
rect 800 89688 179675 89968
rect 800 89288 179755 89688
rect 880 89008 179755 89288
rect 800 88608 179755 89008
rect 800 88328 179675 88608
rect 800 87928 179755 88328
rect 880 87648 179755 87928
rect 800 87248 179755 87648
rect 800 86968 179675 87248
rect 800 86568 179755 86968
rect 880 86288 179755 86568
rect 800 85888 179755 86288
rect 800 85608 179675 85888
rect 800 84528 179755 85608
rect 880 84248 179675 84528
rect 800 83168 179755 84248
rect 880 82888 179675 83168
rect 800 81808 179755 82888
rect 880 81528 179675 81808
rect 800 80448 179755 81528
rect 880 80168 179675 80448
rect 800 79088 179755 80168
rect 880 78808 179675 79088
rect 800 77728 179755 78808
rect 880 77448 179675 77728
rect 800 76368 179755 77448
rect 880 76088 179675 76368
rect 800 75008 179755 76088
rect 880 74728 179755 75008
rect 800 74328 179755 74728
rect 800 74048 179675 74328
rect 800 73648 179755 74048
rect 880 73368 179755 73648
rect 800 72968 179755 73368
rect 800 72688 179675 72968
rect 800 72288 179755 72688
rect 880 72008 179755 72288
rect 800 71608 179755 72008
rect 800 71328 179675 71608
rect 800 70928 179755 71328
rect 880 70648 179755 70928
rect 800 70248 179755 70648
rect 800 69968 179675 70248
rect 800 69568 179755 69968
rect 880 69288 179755 69568
rect 800 68888 179755 69288
rect 800 68608 179675 68888
rect 800 68208 179755 68608
rect 880 67928 179755 68208
rect 800 67528 179755 67928
rect 800 67248 179675 67528
rect 800 66848 179755 67248
rect 880 66568 179755 66848
rect 800 66168 179755 66568
rect 800 65888 179675 66168
rect 800 65488 179755 65888
rect 880 65208 179755 65488
rect 800 64808 179755 65208
rect 800 64528 179675 64808
rect 800 63448 179755 64528
rect 880 63168 179675 63448
rect 800 62088 179755 63168
rect 880 61808 179675 62088
rect 800 60728 179755 61808
rect 880 60448 179675 60728
rect 800 59368 179755 60448
rect 880 59088 179675 59368
rect 800 58008 179755 59088
rect 880 57728 179675 58008
rect 800 56648 179755 57728
rect 880 56368 179675 56648
rect 800 55288 179755 56368
rect 880 55008 179675 55288
rect 800 53928 179755 55008
rect 880 53648 179755 53928
rect 800 53248 179755 53648
rect 800 52968 179675 53248
rect 800 52568 179755 52968
rect 880 52288 179755 52568
rect 800 51888 179755 52288
rect 800 51608 179675 51888
rect 800 51208 179755 51608
rect 880 50928 179755 51208
rect 800 50528 179755 50928
rect 800 50248 179675 50528
rect 800 49848 179755 50248
rect 880 49568 179755 49848
rect 800 49168 179755 49568
rect 800 48888 179675 49168
rect 800 48488 179755 48888
rect 880 48208 179755 48488
rect 800 47808 179755 48208
rect 800 47528 179675 47808
rect 800 47128 179755 47528
rect 880 46848 179755 47128
rect 800 46448 179755 46848
rect 800 46168 179675 46448
rect 800 45768 179755 46168
rect 880 45488 179755 45768
rect 800 45088 179755 45488
rect 800 44808 179675 45088
rect 800 44408 179755 44808
rect 880 44128 179755 44408
rect 800 43728 179755 44128
rect 800 43448 179675 43728
rect 800 42368 179755 43448
rect 880 42088 179675 42368
rect 800 41008 179755 42088
rect 880 40728 179675 41008
rect 800 39648 179755 40728
rect 880 39368 179675 39648
rect 800 38288 179755 39368
rect 880 38008 179675 38288
rect 800 36928 179755 38008
rect 880 36648 179675 36928
rect 800 35568 179755 36648
rect 880 35288 179675 35568
rect 800 34208 179755 35288
rect 880 33928 179675 34208
rect 800 32848 179755 33928
rect 880 32568 179755 32848
rect 800 32168 179755 32568
rect 800 31888 179675 32168
rect 800 31488 179755 31888
rect 880 31208 179755 31488
rect 800 30808 179755 31208
rect 800 30528 179675 30808
rect 800 30128 179755 30528
rect 880 29848 179755 30128
rect 800 29448 179755 29848
rect 800 29168 179675 29448
rect 800 28768 179755 29168
rect 880 28488 179755 28768
rect 800 28088 179755 28488
rect 800 27808 179675 28088
rect 800 27408 179755 27808
rect 880 27128 179755 27408
rect 800 26728 179755 27128
rect 800 26448 179675 26728
rect 800 26048 179755 26448
rect 880 25768 179755 26048
rect 800 25368 179755 25768
rect 800 25088 179675 25368
rect 800 24688 179755 25088
rect 880 24408 179755 24688
rect 800 24008 179755 24408
rect 800 23728 179675 24008
rect 800 23328 179755 23728
rect 880 23048 179755 23328
rect 800 22648 179755 23048
rect 800 22368 179675 22648
rect 800 21288 179755 22368
rect 880 21008 179675 21288
rect 800 19928 179755 21008
rect 880 19648 179675 19928
rect 800 18568 179755 19648
rect 880 18288 179675 18568
rect 800 17208 179755 18288
rect 880 16928 179675 17208
rect 800 15848 179755 16928
rect 880 15568 179675 15848
rect 800 14488 179755 15568
rect 880 14208 179675 14488
rect 800 13128 179755 14208
rect 880 12848 179675 13128
rect 800 11768 179755 12848
rect 880 11488 179755 11768
rect 800 11088 179755 11488
rect 800 10808 179675 11088
rect 800 10408 179755 10808
rect 880 10128 179755 10408
rect 800 9728 179755 10128
rect 800 9448 179675 9728
rect 800 9048 179755 9448
rect 880 8768 179755 9048
rect 800 8368 179755 8768
rect 800 8088 179675 8368
rect 800 7688 179755 8088
rect 880 7408 179755 7688
rect 800 7008 179755 7408
rect 800 6728 179675 7008
rect 800 6328 179755 6728
rect 880 6048 179755 6328
rect 800 5648 179755 6048
rect 800 5368 179675 5648
rect 800 4968 179755 5368
rect 880 4688 179755 4968
rect 800 4288 179755 4688
rect 800 4008 179675 4288
rect 800 3608 179755 4008
rect 880 3328 179755 3608
rect 800 2928 179755 3328
rect 800 2648 179675 2928
rect 800 2248 179755 2648
rect 880 1968 179755 2248
rect 800 1568 179755 1968
rect 800 1395 179675 1568
<< metal4 >>
rect -8576 -7504 -7976 189744
rect -7636 -6564 -7036 188804
rect -6696 -5624 -6096 187864
rect -5756 -4684 -5156 186924
rect -4816 -3744 -4216 185984
rect -3876 -2804 -3276 185044
rect -2936 -1864 -2336 184104
rect -1996 -924 -1396 183164
rect 804 -1864 1404 184104
rect 4404 -3744 5004 185984
rect 8004 -5624 8604 187864
rect 11604 -7504 12204 189744
rect 18804 -1864 19404 184104
rect 22404 -3744 23004 185984
rect 26004 -5624 26604 187864
rect 29604 -7504 30204 189744
rect 36804 -1864 37404 184104
rect 40404 -3744 41004 185984
rect 44004 -5624 44604 187864
rect 47604 -7504 48204 189744
rect 54804 -1864 55404 184104
rect 58404 -3744 59004 185984
rect 62004 -5624 62604 187864
rect 65604 -7504 66204 189744
rect 72804 -1864 73404 184104
rect 76404 -3744 77004 185984
rect 80004 -5624 80604 187864
rect 83604 -7504 84204 189744
rect 90804 -1864 91404 184104
rect 94404 -3744 95004 185984
rect 98004 -5624 98604 187864
rect 101604 -7504 102204 189744
rect 108804 -1864 109404 184104
rect 112404 -3744 113004 185984
rect 116004 -5624 116604 187864
rect 119604 -7504 120204 189744
rect 126804 -1864 127404 184104
rect 130404 -3744 131004 185984
rect 134004 -5624 134604 187864
rect 137604 -7504 138204 189744
rect 144804 -1864 145404 184104
rect 148404 -3744 149004 185984
rect 152004 -5624 152604 187864
rect 155604 -7504 156204 189744
rect 162804 -1864 163404 184104
rect 166404 -3744 167004 185984
rect 170004 -5624 170604 187864
rect 173604 -7504 174204 189744
rect 181900 -924 182500 183164
rect 182840 -1864 183440 184104
rect 183780 -2804 184380 185044
rect 184720 -3744 185320 185984
rect 185660 -4684 186260 186924
rect 186600 -5624 187200 187864
rect 187540 -6564 188140 188804
rect 188480 -7504 189080 189744
<< obsm4 >>
rect 6683 3435 7924 178941
rect 8684 3435 11524 178941
rect 12284 3435 18724 178941
rect 19484 3435 22324 178941
rect 23084 3435 25924 178941
rect 26684 3435 29524 178941
rect 30284 3435 36724 178941
rect 37484 3435 40324 178941
rect 41084 3435 43924 178941
rect 44684 3435 47524 178941
rect 48284 3435 54724 178941
rect 55484 3435 58324 178941
rect 59084 3435 61924 178941
rect 62684 3435 65524 178941
rect 66284 3435 72724 178941
rect 73484 3435 76324 178941
rect 77084 3435 79924 178941
rect 80684 3435 83524 178941
rect 84284 3435 90724 178941
rect 91484 3435 94324 178941
rect 95084 3435 97924 178941
rect 98684 3435 101524 178941
rect 102284 3435 108724 178941
rect 109484 3435 112324 178941
rect 113084 3435 115924 178941
rect 116684 3435 119524 178941
rect 120284 3435 126724 178941
rect 127484 3435 130324 178941
rect 131084 3435 133924 178941
rect 134684 3435 137524 178941
rect 138284 3435 144724 178941
rect 145484 3435 148324 178941
rect 149084 3435 151924 178941
rect 152684 3435 155524 178941
rect 156284 3435 162724 178941
rect 163484 3435 166324 178941
rect 167084 3435 169924 178941
rect 170684 3435 173524 178941
rect 174284 3435 177869 178941
<< metal5 >>
rect -8576 189144 189080 189744
rect -7636 188204 188140 188804
rect -6696 187264 187200 187864
rect -5756 186324 186260 186924
rect -4816 185384 185320 185984
rect -3876 184444 184380 185044
rect -2936 183504 183440 184104
rect -1996 182564 182500 183164
rect -8576 174676 189080 175276
rect -6696 171076 187200 171676
rect -4816 167476 185320 168076
rect -2936 163828 183440 164428
rect -8576 156676 189080 157276
rect -6696 153076 187200 153676
rect -4816 149476 185320 150076
rect -2936 145828 183440 146428
rect -8576 138676 189080 139276
rect -6696 135076 187200 135676
rect -4816 131476 185320 132076
rect -2936 127828 183440 128428
rect -8576 120676 189080 121276
rect -6696 117076 187200 117676
rect -4816 113476 185320 114076
rect -2936 109828 183440 110428
rect -8576 102676 189080 103276
rect -6696 99076 187200 99676
rect -4816 95476 185320 96076
rect -2936 91828 183440 92428
rect -8576 84676 189080 85276
rect -6696 81076 187200 81676
rect -4816 77476 185320 78076
rect -2936 73828 183440 74428
rect -8576 66676 189080 67276
rect -6696 63076 187200 63676
rect -4816 59476 185320 60076
rect -2936 55828 183440 56428
rect -8576 48676 189080 49276
rect -6696 45076 187200 45676
rect -4816 41476 185320 42076
rect -2936 37828 183440 38428
rect -8576 30676 189080 31276
rect -6696 27076 187200 27676
rect -4816 23476 185320 24076
rect -2936 19828 183440 20428
rect -8576 12676 189080 13276
rect -6696 9076 187200 9676
rect -4816 5476 185320 6076
rect -2936 1828 183440 2428
rect -1996 -924 182500 -324
rect -2936 -1864 183440 -1264
rect -3876 -2804 184380 -2204
rect -4816 -3744 185320 -3144
rect -5756 -4684 186260 -4084
rect -6696 -5624 187200 -5024
rect -7636 -6564 188140 -5964
rect -8576 -7504 189080 -6904
<< obsm5 >>
rect -8576 189744 -7976 189746
rect 29604 189744 30204 189746
rect 65604 189744 66204 189746
rect 101604 189744 102204 189746
rect 137604 189744 138204 189746
rect 173604 189744 174204 189746
rect 188480 189744 189080 189746
rect -8576 189142 -7976 189144
rect 29604 189142 30204 189144
rect 65604 189142 66204 189144
rect 101604 189142 102204 189144
rect 137604 189142 138204 189144
rect 173604 189142 174204 189144
rect 188480 189142 189080 189144
rect -7636 188804 -7036 188806
rect 11604 188804 12204 188806
rect 47604 188804 48204 188806
rect 83604 188804 84204 188806
rect 119604 188804 120204 188806
rect 155604 188804 156204 188806
rect 187540 188804 188140 188806
rect -7636 188202 -7036 188204
rect 11604 188202 12204 188204
rect 47604 188202 48204 188204
rect 83604 188202 84204 188204
rect 119604 188202 120204 188204
rect 155604 188202 156204 188204
rect 187540 188202 188140 188204
rect -6696 187864 -6096 187866
rect 26004 187864 26604 187866
rect 62004 187864 62604 187866
rect 98004 187864 98604 187866
rect 134004 187864 134604 187866
rect 170004 187864 170604 187866
rect 186600 187864 187200 187866
rect -6696 187262 -6096 187264
rect 26004 187262 26604 187264
rect 62004 187262 62604 187264
rect 98004 187262 98604 187264
rect 134004 187262 134604 187264
rect 170004 187262 170604 187264
rect 186600 187262 187200 187264
rect -5756 186924 -5156 186926
rect 8004 186924 8604 186926
rect 44004 186924 44604 186926
rect 80004 186924 80604 186926
rect 116004 186924 116604 186926
rect 152004 186924 152604 186926
rect 185660 186924 186260 186926
rect -5756 186322 -5156 186324
rect 8004 186322 8604 186324
rect 44004 186322 44604 186324
rect 80004 186322 80604 186324
rect 116004 186322 116604 186324
rect 152004 186322 152604 186324
rect 185660 186322 186260 186324
rect -4816 185984 -4216 185986
rect 22404 185984 23004 185986
rect 58404 185984 59004 185986
rect 94404 185984 95004 185986
rect 130404 185984 131004 185986
rect 166404 185984 167004 185986
rect 184720 185984 185320 185986
rect -4816 185382 -4216 185384
rect 22404 185382 23004 185384
rect 58404 185382 59004 185384
rect 94404 185382 95004 185384
rect 130404 185382 131004 185384
rect 166404 185382 167004 185384
rect 184720 185382 185320 185384
rect -3876 185044 -3276 185046
rect 4404 185044 5004 185046
rect 40404 185044 41004 185046
rect 76404 185044 77004 185046
rect 112404 185044 113004 185046
rect 148404 185044 149004 185046
rect 183780 185044 184380 185046
rect -3876 184442 -3276 184444
rect 4404 184442 5004 184444
rect 40404 184442 41004 184444
rect 76404 184442 77004 184444
rect 112404 184442 113004 184444
rect 148404 184442 149004 184444
rect 183780 184442 184380 184444
rect -2936 184104 -2336 184106
rect 18804 184104 19404 184106
rect 54804 184104 55404 184106
rect 90804 184104 91404 184106
rect 126804 184104 127404 184106
rect 162804 184104 163404 184106
rect 182840 184104 183440 184106
rect -2936 183502 -2336 183504
rect 18804 183502 19404 183504
rect 54804 183502 55404 183504
rect 90804 183502 91404 183504
rect 126804 183502 127404 183504
rect 162804 183502 163404 183504
rect 182840 183502 183440 183504
rect -1996 183164 -1396 183166
rect 804 183164 1404 183166
rect 36804 183164 37404 183166
rect 72804 183164 73404 183166
rect 108804 183164 109404 183166
rect 144804 183164 145404 183166
rect 181900 183164 182500 183166
rect -1996 182562 -1396 182564
rect 181900 182562 182500 182564
rect 0 175596 180555 182244
rect -8576 175276 -7976 175278
rect 188480 175276 189080 175278
rect -8576 174674 -7976 174676
rect 188480 174674 189080 174676
rect 0 171996 180555 174356
rect -6696 171676 -6096 171678
rect 186600 171676 187200 171678
rect -6696 171074 -6096 171076
rect 186600 171074 187200 171076
rect 0 168396 180555 170756
rect -4816 168076 -4216 168078
rect 184720 168076 185320 168078
rect -4816 167474 -4216 167476
rect 184720 167474 185320 167476
rect 0 164748 180555 167156
rect -2936 164428 -2336 164430
rect 182840 164428 183440 164430
rect -2936 163826 -2336 163828
rect 182840 163826 183440 163828
rect 0 157596 180555 163508
rect -7636 157276 -7036 157278
rect 187540 157276 188140 157278
rect -7636 156674 -7036 156676
rect 187540 156674 188140 156676
rect 0 153996 180555 156356
rect -5756 153676 -5156 153678
rect 185660 153676 186260 153678
rect -5756 153074 -5156 153076
rect 185660 153074 186260 153076
rect 0 150396 180555 152756
rect -3876 150076 -3276 150078
rect 183780 150076 184380 150078
rect -3876 149474 -3276 149476
rect 183780 149474 184380 149476
rect 0 146748 180555 149156
rect -1996 146428 -1396 146430
rect 181900 146428 182500 146430
rect -1996 145826 -1396 145828
rect 181900 145826 182500 145828
rect 0 139596 180555 145508
rect -8576 139276 -7976 139278
rect 188480 139276 189080 139278
rect -8576 138674 -7976 138676
rect 188480 138674 189080 138676
rect 0 135996 180555 138356
rect -6696 135676 -6096 135678
rect 186600 135676 187200 135678
rect -6696 135074 -6096 135076
rect 186600 135074 187200 135076
rect 0 132396 180555 134756
rect -4816 132076 -4216 132078
rect 184720 132076 185320 132078
rect -4816 131474 -4216 131476
rect 184720 131474 185320 131476
rect 0 128748 180555 131156
rect -2936 128428 -2336 128430
rect 182840 128428 183440 128430
rect -2936 127826 -2336 127828
rect 182840 127826 183440 127828
rect 0 121596 180555 127508
rect -7636 121276 -7036 121278
rect 187540 121276 188140 121278
rect -7636 120674 -7036 120676
rect 187540 120674 188140 120676
rect 0 117996 180555 120356
rect -5756 117676 -5156 117678
rect 185660 117676 186260 117678
rect -5756 117074 -5156 117076
rect 185660 117074 186260 117076
rect 0 114396 180555 116756
rect -3876 114076 -3276 114078
rect 183780 114076 184380 114078
rect -3876 113474 -3276 113476
rect 183780 113474 184380 113476
rect 0 110748 180555 113156
rect -1996 110428 -1396 110430
rect 181900 110428 182500 110430
rect -1996 109826 -1396 109828
rect 181900 109826 182500 109828
rect 0 103596 180555 109508
rect -8576 103276 -7976 103278
rect 188480 103276 189080 103278
rect -8576 102674 -7976 102676
rect 188480 102674 189080 102676
rect 0 99996 180555 102356
rect -6696 99676 -6096 99678
rect 186600 99676 187200 99678
rect -6696 99074 -6096 99076
rect 186600 99074 187200 99076
rect 0 96396 180555 98756
rect -4816 96076 -4216 96078
rect 184720 96076 185320 96078
rect -4816 95474 -4216 95476
rect 184720 95474 185320 95476
rect 0 92748 180555 95156
rect -2936 92428 -2336 92430
rect 182840 92428 183440 92430
rect -2936 91826 -2336 91828
rect 182840 91826 183440 91828
rect 0 85596 180555 91508
rect -7636 85276 -7036 85278
rect 187540 85276 188140 85278
rect -7636 84674 -7036 84676
rect 187540 84674 188140 84676
rect 0 81996 180555 84356
rect -5756 81676 -5156 81678
rect 185660 81676 186260 81678
rect -5756 81074 -5156 81076
rect 185660 81074 186260 81076
rect 0 78396 180555 80756
rect -3876 78076 -3276 78078
rect 183780 78076 184380 78078
rect -3876 77474 -3276 77476
rect 183780 77474 184380 77476
rect 0 74748 180555 77156
rect -1996 74428 -1396 74430
rect 181900 74428 182500 74430
rect -1996 73826 -1396 73828
rect 181900 73826 182500 73828
rect 0 67596 180555 73508
rect -8576 67276 -7976 67278
rect 188480 67276 189080 67278
rect -8576 66674 -7976 66676
rect 188480 66674 189080 66676
rect 0 63996 180555 66356
rect -6696 63676 -6096 63678
rect 186600 63676 187200 63678
rect -6696 63074 -6096 63076
rect 186600 63074 187200 63076
rect 0 60396 180555 62756
rect -4816 60076 -4216 60078
rect 184720 60076 185320 60078
rect -4816 59474 -4216 59476
rect 184720 59474 185320 59476
rect 0 56748 180555 59156
rect -2936 56428 -2336 56430
rect 182840 56428 183440 56430
rect -2936 55826 -2336 55828
rect 182840 55826 183440 55828
rect 0 49596 180555 55508
rect -7636 49276 -7036 49278
rect 187540 49276 188140 49278
rect -7636 48674 -7036 48676
rect 187540 48674 188140 48676
rect 0 45996 180555 48356
rect -5756 45676 -5156 45678
rect 185660 45676 186260 45678
rect -5756 45074 -5156 45076
rect 185660 45074 186260 45076
rect 0 42396 180555 44756
rect -3876 42076 -3276 42078
rect 183780 42076 184380 42078
rect -3876 41474 -3276 41476
rect 183780 41474 184380 41476
rect 0 38748 180555 41156
rect -1996 38428 -1396 38430
rect 181900 38428 182500 38430
rect -1996 37826 -1396 37828
rect 181900 37826 182500 37828
rect 0 31596 180555 37508
rect -8576 31276 -7976 31278
rect 188480 31276 189080 31278
rect -8576 30674 -7976 30676
rect 188480 30674 189080 30676
rect 0 27996 180555 30356
rect -6696 27676 -6096 27678
rect 186600 27676 187200 27678
rect -6696 27074 -6096 27076
rect 186600 27074 187200 27076
rect 0 24396 180555 26756
rect -4816 24076 -4216 24078
rect 184720 24076 185320 24078
rect -4816 23474 -4216 23476
rect 184720 23474 185320 23476
rect 0 20748 180555 23156
rect -2936 20428 -2336 20430
rect 182840 20428 183440 20430
rect -2936 19826 -2336 19828
rect 182840 19826 183440 19828
rect 0 13596 180555 19508
rect -7636 13276 -7036 13278
rect 187540 13276 188140 13278
rect -7636 12674 -7036 12676
rect 187540 12674 188140 12676
rect 0 9996 180555 12356
rect -5756 9676 -5156 9678
rect 185660 9676 186260 9678
rect -5756 9074 -5156 9076
rect 185660 9074 186260 9076
rect 0 6396 180555 8756
rect -3876 6076 -3276 6078
rect 183780 6076 184380 6078
rect -3876 5474 -3276 5476
rect 183780 5474 184380 5476
rect 0 2748 180555 5156
rect -1996 2428 -1396 2430
rect 181900 2428 182500 2430
rect -1996 1826 -1396 1828
rect 181900 1826 182500 1828
rect 0 0 180555 1508
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 181900 -324 182500 -322
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 181900 -926 182500 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 182840 -1264 183440 -1262
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 182840 -1866 183440 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 183780 -2204 184380 -2202
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 183780 -2806 184380 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 184720 -3144 185320 -3142
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 184720 -3746 185320 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 185660 -4084 186260 -4082
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 185660 -4686 186260 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 186600 -5024 187200 -5022
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 186600 -5626 187200 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 187540 -5964 188140 -5962
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 187540 -6566 188140 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 188480 -6904 189080 -6902
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 188480 -7506 189080 -7504
<< labels >>
rlabel metal2 s 4618 181899 4674 182699 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 179755 140768 180555 140888 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 139858 0 139914 800 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal3 s 0 174768 800 174888 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal3 s 179755 143488 180555 143608 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 161018 0 161074 800 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal3 s 0 131248 800 131368 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 8758 0 8814 800 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 122838 0 122894 800 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal2 s 97078 0 97134 800 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 109498 181899 109554 182699 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal2 s 169298 0 169354 800 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 0 2048 800 2168 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal2 s 106738 0 106794 800 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 179755 74128 180555 74248 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 118698 181899 118754 182699 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal2 s 110418 0 110474 800 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal2 s 134798 181899 134854 182699 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal2 s 10598 0 10654 800 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 0 59168 800 59288 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 179755 118328 180555 118448 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 0 78888 800 79008 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 179755 168648 180555 168768 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal2 s 114098 0 114154 800 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 0 176128 800 176248 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal2 s 51538 0 51594 800 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal2 s 85578 0 85634 800 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 146298 181899 146354 182699 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal3 s 179755 93848 180555 93968 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal2 s 162858 0 162914 800 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 io_in[10]
port 31 nsew signal input
rlabel metal2 s 168378 181899 168434 182699 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 io_in[12]
port 33 nsew signal input
rlabel metal2 s 62578 181899 62634 182699 6 io_in[13]
port 34 nsew signal input
rlabel metal2 s 32218 181899 32274 182699 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 143538 0 143594 800 6 io_in[15]
port 36 nsew signal input
rlabel metal3 s 0 115608 800 115728 6 io_in[16]
port 37 nsew signal input
rlabel metal3 s 179755 106768 180555 106888 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 161478 181899 161534 182699 6 io_in[18]
port 39 nsew signal input
rlabel metal3 s 179755 2728 180555 2848 6 io_in[19]
port 40 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 105358 181899 105414 182699 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 111338 181899 111394 182699 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 68558 181899 68614 182699 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s 0 114248 800 114368 6 io_in[24]
port 46 nsew signal input
rlabel metal3 s 179755 85688 180555 85808 6 io_in[25]
port 47 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 io_in[26]
port 48 nsew signal input
rlabel metal2 s 46478 181899 46534 182699 6 io_in[27]
port 49 nsew signal input
rlabel metal2 s 47398 181899 47454 182699 6 io_in[28]
port 50 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 io_in[29]
port 51 nsew signal input
rlabel metal2 s 149978 181899 150034 182699 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s 179755 15648 180555 15768 6 io_in[30]
port 53 nsew signal input
rlabel metal3 s 179755 9528 180555 9648 6 io_in[31]
port 54 nsew signal input
rlabel metal2 s 14278 181899 14334 182699 6 io_in[32]
port 55 nsew signal input
rlabel metal3 s 0 181568 800 181688 6 io_in[33]
port 56 nsew signal input
rlabel metal3 s 179755 134648 180555 134768 6 io_in[34]
port 57 nsew signal input
rlabel metal2 s 176198 0 176254 800 6 io_in[35]
port 58 nsew signal input
rlabel metal2 s 84658 181899 84714 182699 6 io_in[36]
port 59 nsew signal input
rlabel metal2 s 23938 181899 23994 182699 6 io_in[37]
port 60 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 io_in[3]
port 61 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 179755 29248 180555 29368 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 0 152328 800 152448 6 io_in[6]
port 64 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 io_in[7]
port 65 nsew signal input
rlabel metal2 s 169298 181899 169354 182699 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 179755 161848 180555 161968 6 io_in[9]
port 67 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 io_oeb[0]
port 68 nsew signal output
rlabel metal2 s 166538 0 166594 800 6 io_oeb[10]
port 69 nsew signal output
rlabel metal2 s 149518 0 149574 800 6 io_oeb[11]
port 70 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 io_oeb[12]
port 71 nsew signal output
rlabel metal2 s 59818 181899 59874 182699 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 179755 104048 180555 104168 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 157798 181899 157854 182699 6 io_oeb[15]
port 74 nsew signal output
rlabel metal3 s 179755 40808 180555 40928 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 165158 181899 165214 182699 6 io_oeb[18]
port 77 nsew signal output
rlabel metal3 s 179755 67328 180555 67448 6 io_oeb[19]
port 78 nsew signal output
rlabel metal2 s 132498 0 132554 800 6 io_oeb[1]
port 79 nsew signal output
rlabel metal3 s 179755 109488 180555 109608 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 15198 181899 15254 182699 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 156878 0 156934 800 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s 179755 30608 180555 30728 6 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s 0 172048 800 172168 6 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s 0 87728 800 87848 6 io_oeb[26]
port 86 nsew signal output
rlabel metal2 s 81898 181899 81954 182699 6 io_oeb[27]
port 87 nsew signal output
rlabel metal2 s 37278 181899 37334 182699 6 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 io_oeb[29]
port 89 nsew signal output
rlabel metal2 s 86958 0 87014 800 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s 0 138048 800 138168 6 io_oeb[30]
port 91 nsew signal output
rlabel metal2 s 37278 0 37334 800 6 io_oeb[31]
port 92 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s 179755 25168 180555 25288 6 io_oeb[33]
port 94 nsew signal output
rlabel metal2 s 53378 181899 53434 182699 6 io_oeb[34]
port 95 nsew signal output
rlabel metal2 s 73618 0 73674 800 6 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 io_oeb[36]
port 97 nsew signal output
rlabel metal2 s 24858 181899 24914 182699 6 io_oeb[37]
port 98 nsew signal output
rlabel metal2 s 179878 0 179934 800 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 0 46928 800 47048 6 io_oeb[4]
port 100 nsew signal output
rlabel metal2 s 155038 0 155094 800 6 io_oeb[5]
port 101 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 io_oeb[6]
port 102 nsew signal output
rlabel metal2 s 39118 181899 39174 182699 6 io_oeb[7]
port 103 nsew signal output
rlabel metal2 s 113178 0 113234 800 6 io_oeb[8]
port 104 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 io_oeb[9]
port 105 nsew signal output
rlabel metal2 s 82818 181899 82874 182699 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 io_out[10]
port 107 nsew signal output
rlabel metal2 s 89718 0 89774 800 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 179755 110848 180555 110968 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 0 108808 800 108928 6 io_out[13]
port 110 nsew signal output
rlabel metal2 s 105818 0 105874 800 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 158718 181899 158774 182699 6 io_out[15]
port 112 nsew signal output
rlabel metal3 s 179755 174088 180555 174208 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 10598 181899 10654 182699 6 io_out[17]
port 114 nsew signal output
rlabel metal3 s 179755 26528 180555 26648 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 0 157768 800 157888 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 121458 181899 121514 182699 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 80058 181899 80114 182699 6 io_out[21]
port 119 nsew signal output
rlabel metal3 s 0 132608 800 132728 6 io_out[22]
port 120 nsew signal output
rlabel metal3 s 0 72088 800 72208 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s 179755 155728 180555 155848 6 io_out[24]
port 122 nsew signal output
rlabel metal2 s 78218 0 78274 800 6 io_out[25]
port 123 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 io_out[26]
port 124 nsew signal output
rlabel metal2 s 164238 181899 164294 182699 6 io_out[27]
port 125 nsew signal output
rlabel metal2 s 154118 0 154174 800 6 io_out[28]
port 126 nsew signal output
rlabel metal2 s 108578 0 108634 800 6 io_out[29]
port 127 nsew signal output
rlabel metal2 s 126518 0 126574 800 6 io_out[2]
port 128 nsew signal output
rlabel metal2 s 63498 181899 63554 182699 6 io_out[30]
port 129 nsew signal output
rlabel metal3 s 179755 108128 180555 108248 6 io_out[31]
port 130 nsew signal output
rlabel metal3 s 0 143488 800 143608 6 io_out[32]
port 131 nsew signal output
rlabel metal2 s 70398 181899 70454 182699 6 io_out[33]
port 132 nsew signal output
rlabel metal2 s 3698 181899 3754 182699 6 io_out[34]
port 133 nsew signal output
rlabel metal3 s 179755 81608 180555 81728 6 io_out[35]
port 134 nsew signal output
rlabel metal2 s 12438 181899 12494 182699 6 io_out[36]
port 135 nsew signal output
rlabel metal3 s 0 102688 800 102808 6 io_out[37]
port 136 nsew signal output
rlabel metal2 s 174818 181899 174874 182699 6 io_out[3]
port 137 nsew signal output
rlabel metal2 s 141698 181899 141754 182699 6 io_out[4]
port 138 nsew signal output
rlabel metal2 s 171138 181899 171194 182699 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 0 104048 800 104168 6 io_out[6]
port 140 nsew signal output
rlabel metal2 s 159638 181899 159694 182699 6 io_out[7]
port 141 nsew signal output
rlabel metal2 s 163778 0 163834 800 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 0 101328 800 101448 6 io_out[9]
port 143 nsew signal output
rlabel metal3 s 0 148928 800 149048 6 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 161938 0 161994 800 6 la_data_in[100]
port 145 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 la_data_in[101]
port 146 nsew signal input
rlabel metal3 s 179755 46248 180555 46368 6 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 132958 181899 133014 182699 6 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 la_data_in[104]
port 149 nsew signal input
rlabel metal3 s 0 127848 800 127968 6 la_data_in[105]
port 150 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 la_data_in[106]
port 151 nsew signal input
rlabel metal3 s 179755 138728 180555 138848 6 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 141698 0 141754 800 6 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_data_in[109]
port 154 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 la_data_in[10]
port 155 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 la_data_in[110]
port 156 nsew signal input
rlabel metal3 s 0 139408 800 139528 6 la_data_in[111]
port 157 nsew signal input
rlabel metal3 s 0 144848 800 144968 6 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 164698 0 164754 800 6 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 97078 181899 97134 182699 6 la_data_in[114]
port 160 nsew signal input
rlabel metal3 s 179755 42168 180555 42288 6 la_data_in[115]
port 161 nsew signal input
rlabel metal3 s 179755 113568 180555 113688 6 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 la_data_in[118]
port 164 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 la_data_in[119]
port 165 nsew signal input
rlabel metal3 s 179755 71408 180555 71528 6 la_data_in[11]
port 166 nsew signal input
rlabel metal3 s 0 56448 800 56568 6 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 143538 181899 143594 182699 6 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 55218 181899 55274 182699 6 la_data_in[124]
port 171 nsew signal input
rlabel metal3 s 179755 19728 180555 19848 6 la_data_in[125]
port 172 nsew signal input
rlabel metal3 s 0 90448 800 90568 6 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 19798 181899 19854 182699 6 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 78678 181899 78734 182699 6 la_data_in[12]
port 175 nsew signal input
rlabel metal3 s 0 86368 800 86488 6 la_data_in[13]
port 176 nsew signal input
rlabel metal3 s 179755 175448 180555 175568 6 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 la_data_in[15]
port 178 nsew signal input
rlabel metal3 s 0 147568 800 147688 6 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 938 181899 994 182699 6 la_data_in[17]
port 180 nsew signal input
rlabel metal3 s 0 146208 800 146328 6 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 13358 181899 13414 182699 6 la_data_in[19]
port 182 nsew signal input
rlabel metal3 s 179755 76168 180555 76288 6 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 131118 181899 131174 182699 6 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 110418 181899 110474 182699 6 la_data_in[21]
port 185 nsew signal input
rlabel metal3 s 179755 80248 180555 80368 6 la_data_in[22]
port 186 nsew signal input
rlabel metal3 s 179755 165928 180555 166048 6 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 120538 181899 120594 182699 6 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 142618 0 142674 800 6 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_data_in[27]
port 191 nsew signal input
rlabel metal3 s 179755 34008 180555 34128 6 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 96158 181899 96214 182699 6 la_data_in[2]
port 194 nsew signal input
rlabel metal3 s 179755 60528 180555 60648 6 la_data_in[30]
port 195 nsew signal input
rlabel metal3 s 179755 17008 180555 17128 6 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 34978 181899 35034 182699 6 la_data_in[32]
port 197 nsew signal input
rlabel metal3 s 179755 167288 180555 167408 6 la_data_in[33]
port 198 nsew signal input
rlabel metal3 s 179755 65968 180555 66088 6 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 145378 181899 145434 182699 6 la_data_in[35]
port 200 nsew signal input
rlabel metal3 s 179755 36728 180555 36848 6 la_data_in[36]
port 201 nsew signal input
rlabel metal3 s 0 118328 800 118448 6 la_data_in[37]
port 202 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 173898 181899 173954 182699 6 la_data_in[39]
port 204 nsew signal input
rlabel metal3 s 179755 44888 180555 45008 6 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 153198 181899 153254 182699 6 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_data_in[41]
port 207 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 57058 181899 57114 182699 6 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 128358 181899 128414 182699 6 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 90178 181899 90234 182699 6 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 42798 181899 42854 182699 6 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 30378 181899 30434 182699 6 la_data_in[47]
port 213 nsew signal input
rlabel metal3 s 179755 154368 180555 154488 6 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 6458 181899 6514 182699 6 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 la_data_in[4]
port 216 nsew signal input
rlabel metal3 s 179755 112208 180555 112328 6 la_data_in[50]
port 217 nsew signal input
rlabel metal3 s 0 163208 800 163328 6 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 83738 181899 83794 182699 6 la_data_in[52]
port 219 nsew signal input
rlabel metal3 s 179755 130568 180555 130688 6 la_data_in[53]
port 220 nsew signal input
rlabel metal3 s 179755 157088 180555 157208 6 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 60738 181899 60794 182699 6 la_data_in[55]
port 222 nsew signal input
rlabel metal3 s 0 121048 800 121168 6 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 64418 181899 64474 182699 6 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 170218 0 170274 800 6 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 167458 181899 167514 182699 6 la_data_in[59]
port 226 nsew signal input
rlabel metal3 s 179755 64608 180555 64728 6 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 160558 181899 160614 182699 6 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 89258 181899 89314 182699 6 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 156878 181899 156934 182699 6 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 76838 181899 76894 182699 6 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 92018 181899 92074 182699 6 la_data_in[65]
port 233 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 112258 0 112314 800 6 la_data_in[67]
port 235 nsew signal input
rlabel metal3 s 179755 51688 180555 51808 6 la_data_in[68]
port 236 nsew signal input
rlabel metal3 s 179755 178168 180555 178288 6 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 la_data_in[6]
port 238 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 la_data_in[70]
port 239 nsew signal input
rlabel metal3 s 179755 146208 180555 146328 6 la_data_in[71]
port 240 nsew signal input
rlabel metal3 s 179755 159808 180555 159928 6 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 119618 181899 119674 182699 6 la_data_in[73]
port 242 nsew signal input
rlabel metal3 s 0 91808 800 91928 6 la_data_in[74]
port 243 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 40038 181899 40094 182699 6 la_data_in[78]
port 247 nsew signal input
rlabel metal3 s 179755 92488 180555 92608 6 la_data_in[79]
port 248 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 20718 181899 20774 182699 6 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 155038 181899 155094 182699 6 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 178498 181899 178554 182699 6 la_data_in[84]
port 254 nsew signal input
rlabel metal3 s 0 160488 800 160608 6 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 100758 181899 100814 182699 6 la_data_in[86]
port 256 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 29458 181899 29514 182699 6 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 97998 181899 98054 182699 6 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 138938 0 138994 800 6 la_data_in[8]
port 260 nsew signal input
rlabel metal3 s 179755 116288 180555 116408 6 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 135718 181899 135774 182699 6 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 65798 181899 65854 182699 6 la_data_in[93]
port 264 nsew signal input
rlabel metal3 s 0 168648 800 168768 6 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 147678 0 147734 800 6 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 178038 0 178094 800 6 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 130198 181899 130254 182699 6 la_data_in[98]
port 269 nsew signal input
rlabel metal3 s 179755 99968 180555 100088 6 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 152278 181899 152334 182699 6 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 138018 0 138074 800 6 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 88798 0 88854 800 6 la_data_out[100]
port 273 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 la_data_out[101]
port 274 nsew signal output
rlabel metal3 s 179755 123768 180555 123888 6 la_data_out[102]
port 275 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 102598 181899 102654 182699 6 la_data_out[104]
port 277 nsew signal output
rlabel metal3 s 0 165928 800 166048 6 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 la_data_out[107]
port 280 nsew signal output
rlabel metal3 s 179755 1368 180555 1488 6 la_data_out[108]
port 281 nsew signal output
rlabel metal3 s 0 150968 800 151088 6 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 54298 181899 54354 182699 6 la_data_out[10]
port 283 nsew signal output
rlabel metal3 s 0 95888 800 96008 6 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 34058 181899 34114 182699 6 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 103978 0 104034 800 6 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 144458 181899 144514 182699 6 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 114098 181899 114154 182699 6 la_data_out[114]
port 288 nsew signal output
rlabel metal3 s 0 97248 800 97368 6 la_data_out[115]
port 289 nsew signal output
rlabel metal3 s 0 99968 800 100088 6 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 48318 181899 48374 182699 6 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 43718 181899 43774 182699 6 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 179418 181899 179474 182699 6 la_data_out[119]
port 293 nsew signal output
rlabel metal3 s 179755 136008 180555 136128 6 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 la_data_out[120]
port 295 nsew signal output
rlabel metal3 s 0 173408 800 173528 6 la_data_out[121]
port 296 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 176658 181899 176714 182699 6 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 173438 0 173494 800 6 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 60278 0 60334 800 6 la_data_out[125]
port 300 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 la_data_out[126]
port 301 nsew signal output
rlabel metal3 s 0 167288 800 167408 6 la_data_out[127]
port 302 nsew signal output
rlabel metal3 s 179755 102688 180555 102808 6 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 160098 0 160154 800 6 la_data_out[13]
port 304 nsew signal output
rlabel metal3 s 179755 78888 180555 79008 6 la_data_out[14]
port 305 nsew signal output
rlabel metal3 s 0 126488 800 126608 6 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 175278 0 175334 800 6 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 61658 181899 61714 182699 6 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 124678 0 124734 800 6 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 133878 181899 133934 182699 6 la_data_out[21]
port 313 nsew signal output
rlabel metal3 s 179755 131928 180555 132048 6 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 72238 181899 72294 182699 6 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 66718 181899 66774 182699 6 la_data_out[24]
port 316 nsew signal output
rlabel metal3 s 179755 163208 180555 163328 6 la_data_out[25]
port 317 nsew signal output
rlabel metal3 s 179755 10888 180555 11008 6 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 129278 0 129334 800 6 la_data_out[27]
port 319 nsew signal output
rlabel metal3 s 179755 48968 180555 49088 6 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 la_data_out[2]
port 322 nsew signal output
rlabel metal3 s 179755 82968 180555 83088 6 la_data_out[30]
port 323 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 la_data_out[31]
port 324 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 36358 181899 36414 182699 6 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 la_data_out[34]
port 327 nsew signal output
rlabel metal3 s 179755 87048 180555 87168 6 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 174358 0 174414 800 6 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 151358 0 151414 800 6 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 172978 181899 173034 182699 6 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 la_data_out[39]
port 332 nsew signal output
rlabel metal3 s 0 153688 800 153808 6 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 119158 0 119214 800 6 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 la_data_out[41]
port 335 nsew signal output
rlabel metal3 s 179755 97248 180555 97368 6 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 145838 0 145894 800 6 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 165618 0 165674 800 6 la_data_out[45]
port 339 nsew signal output
rlabel metal3 s 179755 39448 180555 39568 6 la_data_out[46]
port 340 nsew signal output
rlabel metal3 s 179755 23808 180555 23928 6 la_data_out[47]
port 341 nsew signal output
rlabel metal3 s 179755 8168 180555 8288 6 la_data_out[48]
port 342 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 la_data_out[49]
port 343 nsew signal output
rlabel metal3 s 179755 105408 180555 105528 6 la_data_out[4]
port 344 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 127438 181899 127494 182699 6 la_data_out[51]
port 346 nsew signal output
rlabel metal3 s 179755 91128 180555 91248 6 la_data_out[52]
port 347 nsew signal output
rlabel metal3 s 179755 176808 180555 176928 6 la_data_out[53]
port 348 nsew signal output
rlabel metal3 s 179755 180888 180555 181008 6 la_data_out[54]
port 349 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 152278 0 152334 800 6 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 77758 181899 77814 182699 6 la_data_out[58]
port 353 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 155958 181899 156014 182699 6 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 155958 0 156014 800 6 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 la_data_out[61]
port 357 nsew signal output
rlabel metal3 s 0 73448 800 73568 6 la_data_out[62]
port 358 nsew signal output
rlabel metal3 s 179755 50328 180555 50448 6 la_data_out[63]
port 359 nsew signal output
rlabel metal3 s 179755 63248 180555 63368 6 la_data_out[64]
port 360 nsew signal output
rlabel metal3 s 179755 27888 180555 28008 6 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 99838 181899 99894 182699 6 la_data_out[66]
port 362 nsew signal output
rlabel metal3 s 179755 35368 180555 35488 6 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 98918 181899 98974 182699 6 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 la_data_out[69]
port 365 nsew signal output
rlabel metal3 s 0 155048 800 155168 6 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 52458 181899 52514 182699 6 la_data_out[70]
port 367 nsew signal output
rlabel metal3 s 179755 164568 180555 164688 6 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 172058 181899 172114 182699 6 la_data_out[72]
port 369 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 la_data_out[73]
port 370 nsew signal output
rlabel metal3 s 0 122408 800 122528 6 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 la_data_out[77]
port 374 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 104438 181899 104494 182699 6 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 175738 181899 175794 182699 6 la_data_out[7]
port 377 nsew signal output
rlabel metal3 s 179755 121048 180555 121168 6 la_data_out[80]
port 378 nsew signal output
rlabel metal3 s 179755 31968 180555 32088 6 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 86498 181899 86554 182699 6 la_data_out[82]
port 380 nsew signal output
rlabel metal3 s 0 55088 800 55208 6 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 148598 0 148654 800 6 la_data_out[85]
port 383 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 la_data_out[86]
port 384 nsew signal output
rlabel metal3 s 179755 70048 180555 70168 6 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 163318 181899 163374 182699 6 la_data_out[88]
port 386 nsew signal output
rlabel metal3 s 0 123768 800 123888 6 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 125598 181899 125654 182699 6 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 28538 181899 28594 182699 6 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 25778 181899 25834 182699 6 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 124678 181899 124734 182699 6 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 139858 181899 139914 182699 6 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 2318 0 2374 800 6 la_data_out[94]
port 393 nsew signal output
rlabel metal3 s 179755 61888 180555 62008 6 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 57978 181899 58034 182699 6 la_data_out[96]
port 395 nsew signal output
rlabel metal3 s 0 98608 800 98728 6 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 103058 0 103114 800 6 la_data_out[98]
port 397 nsew signal output
rlabel metal3 s 179755 133288 180555 133408 6 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 96158 0 96214 800 6 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 la_oenb[100]
port 401 nsew signal input
rlabel metal3 s 179755 6808 180555 6928 6 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 44638 181899 44694 182699 6 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_oenb[104]
port 405 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 la_oenb[105]
port 406 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 la_oenb[106]
port 407 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 106278 181899 106334 182699 6 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 128358 0 128414 800 6 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 51538 181899 51594 182699 6 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 69478 181899 69534 182699 6 la_oenb[110]
port 412 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 la_oenb[111]
port 413 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 144918 0 144974 800 6 la_oenb[113]
port 415 nsew signal input
rlabel metal3 s 179755 171368 180555 171488 6 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_oenb[115]
port 417 nsew signal input
rlabel metal3 s 0 57808 800 57928 6 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 56138 181899 56194 182699 6 la_oenb[117]
port 419 nsew signal input
rlabel metal3 s 179755 148928 180555 149048 6 la_oenb[118]
port 420 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 162398 181899 162454 182699 6 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 150438 0 150494 800 6 la_oenb[120]
port 423 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 la_oenb[121]
port 424 nsew signal input
rlabel metal3 s 179755 126488 180555 126608 6 la_oenb[122]
port 425 nsew signal input
rlabel metal3 s 179755 18368 180555 18488 6 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 7838 181899 7894 182699 6 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 la_oenb[127]
port 430 nsew signal input
rlabel metal3 s 179755 147568 180555 147688 6 la_oenb[12]
port 431 nsew signal input
rlabel metal3 s 179755 122408 180555 122528 6 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 147218 181899 147274 182699 6 la_oenb[14]
port 433 nsew signal input
rlabel metal3 s 179755 125128 180555 125248 6 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 22098 181899 22154 182699 6 la_oenb[17]
port 436 nsew signal input
rlabel metal3 s 179755 114928 180555 115048 6 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_oenb[19]
port 438 nsew signal input
rlabel metal3 s 0 180208 800 180328 6 la_oenb[1]
port 439 nsew signal input
rlabel metal3 s 179755 95208 180555 95328 6 la_oenb[20]
port 440 nsew signal input
rlabel metal3 s 0 156408 800 156528 6 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 94318 181899 94374 182699 6 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 67638 181899 67694 182699 6 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 140778 181899 140834 182699 6 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 16118 181899 16174 182699 6 la_oenb[27]
port 447 nsew signal input
rlabel metal3 s 179755 14288 180555 14408 6 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_oenb[29]
port 449 nsew signal input
rlabel metal3 s 179755 98608 180555 98728 6 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 la_oenb[31]
port 452 nsew signal input
rlabel metal3 s 179755 72768 180555 72888 6 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 92938 181899 92994 182699 6 la_oenb[33]
port 454 nsew signal input
rlabel metal3 s 179755 57808 180555 57928 6 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 178958 0 179014 800 6 la_oenb[37]
port 458 nsew signal input
rlabel metal3 s 179755 158448 180555 158568 6 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 la_oenb[39]
port 460 nsew signal input
rlabel metal3 s 0 142128 800 142248 6 la_oenb[3]
port 461 nsew signal input
rlabel metal3 s 0 125128 800 125248 6 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 112258 181899 112314 182699 6 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_oenb[42]
port 464 nsew signal input
rlabel metal3 s 179755 77528 180555 77648 6 la_oenb[43]
port 465 nsew signal input
rlabel metal3 s 0 161848 800 161968 6 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 146758 0 146814 800 6 la_oenb[45]
port 467 nsew signal input
rlabel metal3 s 179755 68688 180555 68808 6 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 170218 181899 170274 182699 6 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 73158 181899 73214 182699 6 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 478 0 534 800 6 la_oenb[4]
port 472 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 1858 181899 1914 182699 6 la_oenb[51]
port 474 nsew signal input
rlabel metal3 s 179755 38088 180555 38208 6 la_oenb[52]
port 475 nsew signal input
rlabel metal3 s 179755 88408 180555 88528 6 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_oenb[54]
port 477 nsew signal input
rlabel metal3 s 0 136688 800 136808 6 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 41878 181899 41934 182699 6 la_oenb[56]
port 479 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 153198 0 153254 800 6 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 95238 181899 95294 182699 6 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 122838 181899 122894 182699 6 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 123758 0 123814 800 6 la_oenb[60]
port 484 nsew signal input
rlabel metal3 s 179755 56448 180555 56568 6 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 la_oenb[62]
port 486 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 la_oenb[63]
port 487 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 la_oenb[64]
port 488 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 11518 181899 11574 182699 6 la_oenb[66]
port 490 nsew signal input
rlabel metal3 s 179755 22448 180555 22568 6 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 103518 181899 103574 182699 6 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 140778 0 140834 800 6 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 129278 181899 129334 182699 6 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 50158 181899 50214 182699 6 la_oenb[71]
port 496 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 80978 181899 81034 182699 6 la_oenb[74]
port 499 nsew signal input
rlabel metal3 s 0 170008 800 170128 6 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 18878 181899 18934 182699 6 la_oenb[76]
port 501 nsew signal input
rlabel metal3 s 179755 5448 180555 5568 6 la_oenb[77]
port 502 nsew signal input
rlabel metal3 s 0 178848 800 178968 6 la_oenb[78]
port 503 nsew signal input
rlabel metal3 s 179755 43528 180555 43648 6 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_oenb[7]
port 505 nsew signal input
rlabel metal3 s 179755 151648 180555 151768 6 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 136638 181899 136694 182699 6 la_oenb[81]
port 507 nsew signal input
rlabel metal3 s 0 119688 800 119808 6 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 136178 0 136234 800 6 la_oenb[83]
port 509 nsew signal input
rlabel metal3 s 0 105408 800 105528 6 la_oenb[84]
port 510 nsew signal input
rlabel metal3 s 179755 84328 180555 84448 6 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 154118 181899 154174 182699 6 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 75918 181899 75974 182699 6 la_oenb[87]
port 513 nsew signal input
rlabel metal3 s 179755 172728 180555 172848 6 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_oenb[89]
port 515 nsew signal input
rlabel metal3 s 179755 137368 180555 137488 6 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 115938 181899 115994 182699 6 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 177578 181899 177634 182699 6 la_oenb[93]
port 520 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 la_oenb[94]
port 521 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 la_oenb[96]
port 523 nsew signal input
rlabel metal3 s 179755 150288 180555 150408 6 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 91098 181899 91154 182699 6 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 150898 181899 150954 182699 6 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 user_clock2
port 528 nsew signal input
rlabel metal2 s 26698 181899 26754 182699 6 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 132038 181899 132094 182699 6 user_irq[2]
port 531 nsew signal output
rlabel metal2 s 87418 181899 87474 182699 6 wb_clk_i
port 532 nsew signal input
rlabel metal3 s 179755 4088 180555 4208 6 wb_rst_i
port 533 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 wbs_ack_o
port 534 nsew signal output
rlabel metal2 s 85578 181899 85634 182699 6 wbs_adr_i[0]
port 535 nsew signal input
rlabel metal3 s 179755 53048 180555 53168 6 wbs_adr_i[10]
port 536 nsew signal input
rlabel metal2 s 177118 0 177174 800 6 wbs_adr_i[11]
port 537 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 wbs_adr_i[12]
port 538 nsew signal input
rlabel metal3 s 0 177488 800 177608 6 wbs_adr_i[13]
port 539 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 wbs_adr_i[14]
port 540 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 wbs_adr_i[15]
port 541 nsew signal input
rlabel metal3 s 179755 142128 180555 142248 6 wbs_adr_i[16]
port 542 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 wbs_adr_i[17]
port 543 nsew signal input
rlabel metal3 s 179755 12928 180555 13048 6 wbs_adr_i[18]
port 544 nsew signal input
rlabel metal2 s 108578 181899 108634 182699 6 wbs_adr_i[19]
port 545 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_adr_i[1]
port 546 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 wbs_adr_i[20]
port 547 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_adr_i[21]
port 548 nsew signal input
rlabel metal2 s 130658 0 130714 800 6 wbs_adr_i[22]
port 549 nsew signal input
rlabel metal2 s 74078 181899 74134 182699 6 wbs_adr_i[23]
port 550 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_adr_i[24]
port 551 nsew signal input
rlabel metal2 s 167458 0 167514 800 6 wbs_adr_i[25]
port 552 nsew signal input
rlabel metal3 s 0 140768 800 140888 6 wbs_adr_i[26]
port 553 nsew signal input
rlabel metal2 s 116858 181899 116914 182699 6 wbs_adr_i[27]
port 554 nsew signal input
rlabel metal2 s 9678 181899 9734 182699 6 wbs_adr_i[28]
port 555 nsew signal input
rlabel metal3 s 179755 179528 180555 179648 6 wbs_adr_i[29]
port 556 nsew signal input
rlabel metal2 s 23018 181899 23074 182699 6 wbs_adr_i[2]
port 557 nsew signal input
rlabel metal2 s 71318 181899 71374 182699 6 wbs_adr_i[30]
port 558 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_adr_i[31]
port 559 nsew signal input
rlabel metal3 s 179755 101328 180555 101448 6 wbs_adr_i[3]
port 560 nsew signal input
rlabel metal2 s 38198 181899 38254 182699 6 wbs_adr_i[4]
port 561 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 wbs_adr_i[5]
port 562 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 wbs_adr_i[6]
port 563 nsew signal input
rlabel metal2 s 159178 0 159234 800 6 wbs_adr_i[7]
port 564 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 wbs_adr_i[8]
port 565 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 wbs_adr_i[9]
port 566 nsew signal input
rlabel metal2 s 88338 181899 88394 182699 6 wbs_cyc_i
port 567 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 wbs_dat_i[0]
port 568 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 wbs_dat_i[10]
port 569 nsew signal input
rlabel metal3 s 0 129888 800 130008 6 wbs_dat_i[11]
port 570 nsew signal input
rlabel metal2 s 148138 181899 148194 182699 6 wbs_dat_i[12]
port 571 nsew signal input
rlabel metal3 s 179755 153008 180555 153128 6 wbs_dat_i[13]
port 572 nsew signal input
rlabel metal3 s 179755 55088 180555 55208 6 wbs_dat_i[14]
port 573 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 wbs_dat_i[15]
port 574 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 wbs_dat_i[16]
port 575 nsew signal input
rlabel metal2 s 121918 0 121974 800 6 wbs_dat_i[17]
port 576 nsew signal input
rlabel metal3 s 0 135328 800 135448 6 wbs_dat_i[18]
port 577 nsew signal input
rlabel metal2 s 123758 181899 123814 182699 6 wbs_dat_i[19]
port 578 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 wbs_dat_i[1]
port 579 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 wbs_dat_i[20]
port 580 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_dat_i[21]
port 581 nsew signal input
rlabel metal2 s 166538 181899 166594 182699 6 wbs_dat_i[22]
port 582 nsew signal input
rlabel metal2 s 127438 0 127494 800 6 wbs_dat_i[23]
port 583 nsew signal input
rlabel metal2 s 17958 181899 18014 182699 6 wbs_dat_i[24]
port 584 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 wbs_dat_i[25]
port 585 nsew signal input
rlabel metal3 s 179755 21088 180555 21208 6 wbs_dat_i[26]
port 586 nsew signal input
rlabel metal3 s 179755 59168 180555 59288 6 wbs_dat_i[27]
port 587 nsew signal input
rlabel metal2 s 58898 181899 58954 182699 6 wbs_dat_i[28]
port 588 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 wbs_dat_i[29]
port 589 nsew signal input
rlabel metal3 s 179755 170008 180555 170128 6 wbs_dat_i[2]
port 590 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 wbs_dat_i[30]
port 591 nsew signal input
rlabel metal2 s 45558 181899 45614 182699 6 wbs_dat_i[31]
port 592 nsew signal input
rlabel metal2 s 117778 181899 117834 182699 6 wbs_dat_i[3]
port 593 nsew signal input
rlabel metal3 s 0 159128 800 159248 6 wbs_dat_i[4]
port 594 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_i[5]
port 595 nsew signal input
rlabel metal2 s 142618 181899 142674 182699 6 wbs_dat_i[6]
port 596 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_i[7]
port 597 nsew signal input
rlabel metal2 s 113178 181899 113234 182699 6 wbs_dat_i[8]
port 598 nsew signal input
rlabel metal3 s 0 164568 800 164688 6 wbs_dat_i[9]
port 599 nsew signal input
rlabel metal2 s 5538 181899 5594 182699 6 wbs_dat_o[0]
port 600 nsew signal output
rlabel metal3 s 179755 144848 180555 144968 6 wbs_dat_o[10]
port 601 nsew signal output
rlabel metal2 s 116398 0 116454 800 6 wbs_dat_o[11]
port 602 nsew signal output
rlabel metal2 s 168378 0 168434 800 6 wbs_dat_o[12]
port 603 nsew signal output
rlabel metal2 s 32678 0 32734 800 6 wbs_dat_o[13]
port 604 nsew signal output
rlabel metal3 s 0 133968 800 134088 6 wbs_dat_o[14]
port 605 nsew signal output
rlabel metal2 s 171138 0 171194 800 6 wbs_dat_o[15]
port 606 nsew signal output
rlabel metal2 s 138938 181899 138994 182699 6 wbs_dat_o[16]
port 607 nsew signal output
rlabel metal2 s 2778 181899 2834 182699 6 wbs_dat_o[17]
port 608 nsew signal output
rlabel metal3 s 179755 89768 180555 89888 6 wbs_dat_o[18]
port 609 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 wbs_dat_o[19]
port 610 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 wbs_dat_o[1]
port 611 nsew signal output
rlabel metal2 s 74998 181899 75054 182699 6 wbs_dat_o[20]
port 612 nsew signal output
rlabel metal2 s 40958 181899 41014 182699 6 wbs_dat_o[21]
port 613 nsew signal output
rlabel metal2 s 133418 0 133474 800 6 wbs_dat_o[22]
port 614 nsew signal output
rlabel metal2 s 8758 181899 8814 182699 6 wbs_dat_o[23]
port 615 nsew signal output
rlabel metal2 s 115018 181899 115074 182699 6 wbs_dat_o[24]
port 616 nsew signal output
rlabel metal3 s 179755 119688 180555 119808 6 wbs_dat_o[25]
port 617 nsew signal output
rlabel metal2 s 126518 181899 126574 182699 6 wbs_dat_o[26]
port 618 nsew signal output
rlabel metal2 s 149058 181899 149114 182699 6 wbs_dat_o[27]
port 619 nsew signal output
rlabel metal3 s 179755 47608 180555 47728 6 wbs_dat_o[28]
port 620 nsew signal output
rlabel metal2 s 27618 181899 27674 182699 6 wbs_dat_o[29]
port 621 nsew signal output
rlabel metal3 s 0 111528 800 111648 6 wbs_dat_o[2]
port 622 nsew signal output
rlabel metal2 s 138018 181899 138074 182699 6 wbs_dat_o[30]
port 623 nsew signal output
rlabel metal2 s 49238 181899 49294 182699 6 wbs_dat_o[31]
port 624 nsew signal output
rlabel metal3 s 0 112888 800 113008 6 wbs_dat_o[3]
port 625 nsew signal output
rlabel metal2 s 31298 181899 31354 182699 6 wbs_dat_o[4]
port 626 nsew signal output
rlabel metal2 s 107198 181899 107254 182699 6 wbs_dat_o[5]
port 627 nsew signal output
rlabel metal2 s 80058 0 80114 800 6 wbs_dat_o[6]
port 628 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_o[7]
port 629 nsew signal output
rlabel metal3 s 179755 127848 180555 127968 6 wbs_dat_o[8]
port 630 nsew signal output
rlabel metal3 s 179755 129208 180555 129328 6 wbs_dat_o[9]
port 631 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 wbs_sel_i[0]
port 632 nsew signal input
rlabel metal2 s 17038 181899 17094 182699 6 wbs_sel_i[1]
port 633 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 wbs_sel_i[2]
port 634 nsew signal input
rlabel metal2 s 33138 181899 33194 182699 6 wbs_sel_i[3]
port 635 nsew signal input
rlabel metal2 s 120998 0 121054 800 6 wbs_stb_i
port 636 nsew signal input
rlabel metal2 s 101678 181899 101734 182699 6 wbs_we_i
port 637 nsew signal input
rlabel metal4 s 144804 -1864 145404 184104 6 vccd1
port 638 nsew power bidirectional
rlabel metal4 s 108804 -1864 109404 184104 6 vccd1
port 639 nsew power bidirectional
rlabel metal4 s 72804 -1864 73404 184104 6 vccd1
port 640 nsew power bidirectional
rlabel metal4 s 36804 -1864 37404 184104 6 vccd1
port 641 nsew power bidirectional
rlabel metal4 s 804 -1864 1404 184104 6 vccd1
port 642 nsew power bidirectional
rlabel metal4 s 181900 -924 182500 183164 6 vccd1
port 643 nsew power bidirectional
rlabel metal4 s -1996 -924 -1396 183164 4 vccd1
port 644 nsew power bidirectional
rlabel metal5 s -1996 182564 182500 183164 6 vccd1
port 645 nsew power bidirectional
rlabel metal5 s -2936 145828 183440 146428 6 vccd1
port 646 nsew power bidirectional
rlabel metal5 s -2936 109828 183440 110428 6 vccd1
port 647 nsew power bidirectional
rlabel metal5 s -2936 73828 183440 74428 6 vccd1
port 648 nsew power bidirectional
rlabel metal5 s -2936 37828 183440 38428 6 vccd1
port 649 nsew power bidirectional
rlabel metal5 s -2936 1828 183440 2428 6 vccd1
port 650 nsew power bidirectional
rlabel metal5 s -1996 -924 182500 -324 8 vccd1
port 651 nsew power bidirectional
rlabel metal4 s 182840 -1864 183440 184104 6 vssd1
port 652 nsew ground bidirectional
rlabel metal4 s 162804 -1864 163404 184104 6 vssd1
port 653 nsew ground bidirectional
rlabel metal4 s 126804 -1864 127404 184104 6 vssd1
port 654 nsew ground bidirectional
rlabel metal4 s 90804 -1864 91404 184104 6 vssd1
port 655 nsew ground bidirectional
rlabel metal4 s 54804 -1864 55404 184104 6 vssd1
port 656 nsew ground bidirectional
rlabel metal4 s 18804 -1864 19404 184104 6 vssd1
port 657 nsew ground bidirectional
rlabel metal4 s -2936 -1864 -2336 184104 4 vssd1
port 658 nsew ground bidirectional
rlabel metal5 s -2936 183504 183440 184104 6 vssd1
port 659 nsew ground bidirectional
rlabel metal5 s -2936 163828 183440 164428 6 vssd1
port 660 nsew ground bidirectional
rlabel metal5 s -2936 127828 183440 128428 6 vssd1
port 661 nsew ground bidirectional
rlabel metal5 s -2936 91828 183440 92428 6 vssd1
port 662 nsew ground bidirectional
rlabel metal5 s -2936 55828 183440 56428 6 vssd1
port 663 nsew ground bidirectional
rlabel metal5 s -2936 19828 183440 20428 6 vssd1
port 664 nsew ground bidirectional
rlabel metal5 s -2936 -1864 183440 -1264 8 vssd1
port 665 nsew ground bidirectional
rlabel metal4 s 148404 -3744 149004 185984 6 vccd2
port 666 nsew power bidirectional
rlabel metal4 s 112404 -3744 113004 185984 6 vccd2
port 667 nsew power bidirectional
rlabel metal4 s 76404 -3744 77004 185984 6 vccd2
port 668 nsew power bidirectional
rlabel metal4 s 40404 -3744 41004 185984 6 vccd2
port 669 nsew power bidirectional
rlabel metal4 s 4404 -3744 5004 185984 6 vccd2
port 670 nsew power bidirectional
rlabel metal4 s 183780 -2804 184380 185044 6 vccd2
port 671 nsew power bidirectional
rlabel metal4 s -3876 -2804 -3276 185044 4 vccd2
port 672 nsew power bidirectional
rlabel metal5 s -3876 184444 184380 185044 6 vccd2
port 673 nsew power bidirectional
rlabel metal5 s -4816 149476 185320 150076 6 vccd2
port 674 nsew power bidirectional
rlabel metal5 s -4816 113476 185320 114076 6 vccd2
port 675 nsew power bidirectional
rlabel metal5 s -4816 77476 185320 78076 6 vccd2
port 676 nsew power bidirectional
rlabel metal5 s -4816 41476 185320 42076 6 vccd2
port 677 nsew power bidirectional
rlabel metal5 s -4816 5476 185320 6076 6 vccd2
port 678 nsew power bidirectional
rlabel metal5 s -3876 -2804 184380 -2204 8 vccd2
port 679 nsew power bidirectional
rlabel metal4 s 184720 -3744 185320 185984 6 vssd2
port 680 nsew ground bidirectional
rlabel metal4 s 166404 -3744 167004 185984 6 vssd2
port 681 nsew ground bidirectional
rlabel metal4 s 130404 -3744 131004 185984 6 vssd2
port 682 nsew ground bidirectional
rlabel metal4 s 94404 -3744 95004 185984 6 vssd2
port 683 nsew ground bidirectional
rlabel metal4 s 58404 -3744 59004 185984 6 vssd2
port 684 nsew ground bidirectional
rlabel metal4 s 22404 -3744 23004 185984 6 vssd2
port 685 nsew ground bidirectional
rlabel metal4 s -4816 -3744 -4216 185984 4 vssd2
port 686 nsew ground bidirectional
rlabel metal5 s -4816 185384 185320 185984 6 vssd2
port 687 nsew ground bidirectional
rlabel metal5 s -4816 167476 185320 168076 6 vssd2
port 688 nsew ground bidirectional
rlabel metal5 s -4816 131476 185320 132076 6 vssd2
port 689 nsew ground bidirectional
rlabel metal5 s -4816 95476 185320 96076 6 vssd2
port 690 nsew ground bidirectional
rlabel metal5 s -4816 59476 185320 60076 6 vssd2
port 691 nsew ground bidirectional
rlabel metal5 s -4816 23476 185320 24076 6 vssd2
port 692 nsew ground bidirectional
rlabel metal5 s -4816 -3744 185320 -3144 8 vssd2
port 693 nsew ground bidirectional
rlabel metal4 s 152004 -5624 152604 187864 6 vdda1
port 694 nsew power bidirectional
rlabel metal4 s 116004 -5624 116604 187864 6 vdda1
port 695 nsew power bidirectional
rlabel metal4 s 80004 -5624 80604 187864 6 vdda1
port 696 nsew power bidirectional
rlabel metal4 s 44004 -5624 44604 187864 6 vdda1
port 697 nsew power bidirectional
rlabel metal4 s 8004 -5624 8604 187864 6 vdda1
port 698 nsew power bidirectional
rlabel metal4 s 185660 -4684 186260 186924 6 vdda1
port 699 nsew power bidirectional
rlabel metal4 s -5756 -4684 -5156 186924 4 vdda1
port 700 nsew power bidirectional
rlabel metal5 s -5756 186324 186260 186924 6 vdda1
port 701 nsew power bidirectional
rlabel metal5 s -6696 153076 187200 153676 6 vdda1
port 702 nsew power bidirectional
rlabel metal5 s -6696 117076 187200 117676 6 vdda1
port 703 nsew power bidirectional
rlabel metal5 s -6696 81076 187200 81676 6 vdda1
port 704 nsew power bidirectional
rlabel metal5 s -6696 45076 187200 45676 6 vdda1
port 705 nsew power bidirectional
rlabel metal5 s -6696 9076 187200 9676 6 vdda1
port 706 nsew power bidirectional
rlabel metal5 s -5756 -4684 186260 -4084 8 vdda1
port 707 nsew power bidirectional
rlabel metal4 s 186600 -5624 187200 187864 6 vssa1
port 708 nsew ground bidirectional
rlabel metal4 s 170004 -5624 170604 187864 6 vssa1
port 709 nsew ground bidirectional
rlabel metal4 s 134004 -5624 134604 187864 6 vssa1
port 710 nsew ground bidirectional
rlabel metal4 s 98004 -5624 98604 187864 6 vssa1
port 711 nsew ground bidirectional
rlabel metal4 s 62004 -5624 62604 187864 6 vssa1
port 712 nsew ground bidirectional
rlabel metal4 s 26004 -5624 26604 187864 6 vssa1
port 713 nsew ground bidirectional
rlabel metal4 s -6696 -5624 -6096 187864 4 vssa1
port 714 nsew ground bidirectional
rlabel metal5 s -6696 187264 187200 187864 6 vssa1
port 715 nsew ground bidirectional
rlabel metal5 s -6696 171076 187200 171676 6 vssa1
port 716 nsew ground bidirectional
rlabel metal5 s -6696 135076 187200 135676 6 vssa1
port 717 nsew ground bidirectional
rlabel metal5 s -6696 99076 187200 99676 6 vssa1
port 718 nsew ground bidirectional
rlabel metal5 s -6696 63076 187200 63676 6 vssa1
port 719 nsew ground bidirectional
rlabel metal5 s -6696 27076 187200 27676 6 vssa1
port 720 nsew ground bidirectional
rlabel metal5 s -6696 -5624 187200 -5024 8 vssa1
port 721 nsew ground bidirectional
rlabel metal4 s 155604 -7504 156204 189744 6 vdda2
port 722 nsew power bidirectional
rlabel metal4 s 119604 -7504 120204 189744 6 vdda2
port 723 nsew power bidirectional
rlabel metal4 s 83604 -7504 84204 189744 6 vdda2
port 724 nsew power bidirectional
rlabel metal4 s 47604 -7504 48204 189744 6 vdda2
port 725 nsew power bidirectional
rlabel metal4 s 11604 -7504 12204 189744 6 vdda2
port 726 nsew power bidirectional
rlabel metal4 s 187540 -6564 188140 188804 6 vdda2
port 727 nsew power bidirectional
rlabel metal4 s -7636 -6564 -7036 188804 4 vdda2
port 728 nsew power bidirectional
rlabel metal5 s -7636 188204 188140 188804 6 vdda2
port 729 nsew power bidirectional
rlabel metal5 s -8576 156676 189080 157276 6 vdda2
port 730 nsew power bidirectional
rlabel metal5 s -8576 120676 189080 121276 6 vdda2
port 731 nsew power bidirectional
rlabel metal5 s -8576 84676 189080 85276 6 vdda2
port 732 nsew power bidirectional
rlabel metal5 s -8576 48676 189080 49276 6 vdda2
port 733 nsew power bidirectional
rlabel metal5 s -8576 12676 189080 13276 6 vdda2
port 734 nsew power bidirectional
rlabel metal5 s -7636 -6564 188140 -5964 8 vdda2
port 735 nsew power bidirectional
rlabel metal4 s 188480 -7504 189080 189744 6 vssa2
port 736 nsew ground bidirectional
rlabel metal4 s 173604 -7504 174204 189744 6 vssa2
port 737 nsew ground bidirectional
rlabel metal4 s 137604 -7504 138204 189744 6 vssa2
port 738 nsew ground bidirectional
rlabel metal4 s 101604 -7504 102204 189744 6 vssa2
port 739 nsew ground bidirectional
rlabel metal4 s 65604 -7504 66204 189744 6 vssa2
port 740 nsew ground bidirectional
rlabel metal4 s 29604 -7504 30204 189744 6 vssa2
port 741 nsew ground bidirectional
rlabel metal4 s -8576 -7504 -7976 189744 4 vssa2
port 742 nsew ground bidirectional
rlabel metal5 s -8576 189144 189080 189744 6 vssa2
port 743 nsew ground bidirectional
rlabel metal5 s -8576 174676 189080 175276 6 vssa2
port 744 nsew ground bidirectional
rlabel metal5 s -8576 138676 189080 139276 6 vssa2
port 745 nsew ground bidirectional
rlabel metal5 s -8576 102676 189080 103276 6 vssa2
port 746 nsew ground bidirectional
rlabel metal5 s -8576 66676 189080 67276 6 vssa2
port 747 nsew ground bidirectional
rlabel metal5 s -8576 30676 189080 31276 6 vssa2
port 748 nsew ground bidirectional
rlabel metal5 s -8576 -7504 189080 -6904 8 vssa2
port 749 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180555 182699
string LEFview TRUE
string GDS_FILE /project/openlane/user_project_wrapper/runs/user_project_wrapper/results/magic/user_project_wrapper.gds
string GDS_END 72821766
string GDS_START 130
<< end >>

