magic
tech sky130A
magscale 1 2
timestamp 1622251967
<< obsli1 >>
rect 949 1717 178451 179367
<< obsm1 >>
rect 937 1708 179018 179568
<< metal2 >>
rect 938 181037 994 181837
rect 1858 181037 1914 181837
rect 2778 181037 2834 181837
rect 3698 181037 3754 181837
rect 4618 181037 4674 181837
rect 5538 181037 5594 181837
rect 6458 181037 6514 181837
rect 7378 181037 7434 181837
rect 8298 181037 8354 181837
rect 9218 181037 9274 181837
rect 10138 181037 10194 181837
rect 11058 181037 11114 181837
rect 12438 181037 12494 181837
rect 13358 181037 13414 181837
rect 14278 181037 14334 181837
rect 15198 181037 15254 181837
rect 16118 181037 16174 181837
rect 17038 181037 17094 181837
rect 17958 181037 18014 181837
rect 18878 181037 18934 181837
rect 19798 181037 19854 181837
rect 20718 181037 20774 181837
rect 21638 181037 21694 181837
rect 22558 181037 22614 181837
rect 23478 181037 23534 181837
rect 24398 181037 24454 181837
rect 25318 181037 25374 181837
rect 26238 181037 26294 181837
rect 27158 181037 27214 181837
rect 28078 181037 28134 181837
rect 29458 181037 29514 181837
rect 30378 181037 30434 181837
rect 31298 181037 31354 181837
rect 32218 181037 32274 181837
rect 33138 181037 33194 181837
rect 34058 181037 34114 181837
rect 34978 181037 35034 181837
rect 35898 181037 35954 181837
rect 36818 181037 36874 181837
rect 37738 181037 37794 181837
rect 38658 181037 38714 181837
rect 39578 181037 39634 181837
rect 40498 181037 40554 181837
rect 41418 181037 41474 181837
rect 42338 181037 42394 181837
rect 43258 181037 43314 181837
rect 44178 181037 44234 181837
rect 45558 181037 45614 181837
rect 46478 181037 46534 181837
rect 47398 181037 47454 181837
rect 48318 181037 48374 181837
rect 49238 181037 49294 181837
rect 50158 181037 50214 181837
rect 51078 181037 51134 181837
rect 51998 181037 52054 181837
rect 52918 181037 52974 181837
rect 53838 181037 53894 181837
rect 54758 181037 54814 181837
rect 55678 181037 55734 181837
rect 56598 181037 56654 181837
rect 57518 181037 57574 181837
rect 58438 181037 58494 181837
rect 59358 181037 59414 181837
rect 60278 181037 60334 181837
rect 61198 181037 61254 181837
rect 62578 181037 62634 181837
rect 63498 181037 63554 181837
rect 64418 181037 64474 181837
rect 65338 181037 65394 181837
rect 66258 181037 66314 181837
rect 67178 181037 67234 181837
rect 68098 181037 68154 181837
rect 69018 181037 69074 181837
rect 69938 181037 69994 181837
rect 70858 181037 70914 181837
rect 71778 181037 71834 181837
rect 72698 181037 72754 181837
rect 73618 181037 73674 181837
rect 74538 181037 74594 181837
rect 75458 181037 75514 181837
rect 76378 181037 76434 181837
rect 77298 181037 77354 181837
rect 78218 181037 78274 181837
rect 79598 181037 79654 181837
rect 80518 181037 80574 181837
rect 81438 181037 81494 181837
rect 82358 181037 82414 181837
rect 83278 181037 83334 181837
rect 84198 181037 84254 181837
rect 85118 181037 85174 181837
rect 86038 181037 86094 181837
rect 86958 181037 87014 181837
rect 87878 181037 87934 181837
rect 88798 181037 88854 181837
rect 89718 181037 89774 181837
rect 90638 181037 90694 181837
rect 91558 181037 91614 181837
rect 92478 181037 92534 181837
rect 93398 181037 93454 181837
rect 94318 181037 94374 181837
rect 95238 181037 95294 181837
rect 96618 181037 96674 181837
rect 97538 181037 97594 181837
rect 98458 181037 98514 181837
rect 99378 181037 99434 181837
rect 100298 181037 100354 181837
rect 101218 181037 101274 181837
rect 102138 181037 102194 181837
rect 103058 181037 103114 181837
rect 103978 181037 104034 181837
rect 104898 181037 104954 181837
rect 105818 181037 105874 181837
rect 106738 181037 106794 181837
rect 107658 181037 107714 181837
rect 108578 181037 108634 181837
rect 109498 181037 109554 181837
rect 110418 181037 110474 181837
rect 111338 181037 111394 181837
rect 112718 181037 112774 181837
rect 113638 181037 113694 181837
rect 114558 181037 114614 181837
rect 115478 181037 115534 181837
rect 116398 181037 116454 181837
rect 117318 181037 117374 181837
rect 118238 181037 118294 181837
rect 119158 181037 119214 181837
rect 120078 181037 120134 181837
rect 120998 181037 121054 181837
rect 121918 181037 121974 181837
rect 122838 181037 122894 181837
rect 123758 181037 123814 181837
rect 124678 181037 124734 181837
rect 125598 181037 125654 181837
rect 126518 181037 126574 181837
rect 127438 181037 127494 181837
rect 128358 181037 128414 181837
rect 129738 181037 129794 181837
rect 130658 181037 130714 181837
rect 131578 181037 131634 181837
rect 132498 181037 132554 181837
rect 133418 181037 133474 181837
rect 134338 181037 134394 181837
rect 135258 181037 135314 181837
rect 136178 181037 136234 181837
rect 137098 181037 137154 181837
rect 138018 181037 138074 181837
rect 138938 181037 138994 181837
rect 139858 181037 139914 181837
rect 140778 181037 140834 181837
rect 141698 181037 141754 181837
rect 142618 181037 142674 181837
rect 143538 181037 143594 181837
rect 144458 181037 144514 181837
rect 145378 181037 145434 181837
rect 146758 181037 146814 181837
rect 147678 181037 147734 181837
rect 148598 181037 148654 181837
rect 149518 181037 149574 181837
rect 150438 181037 150494 181837
rect 151358 181037 151414 181837
rect 152278 181037 152334 181837
rect 153198 181037 153254 181837
rect 154118 181037 154174 181837
rect 155038 181037 155094 181837
rect 155958 181037 156014 181837
rect 156878 181037 156934 181837
rect 157798 181037 157854 181837
rect 158718 181037 158774 181837
rect 159638 181037 159694 181837
rect 160558 181037 160614 181837
rect 161478 181037 161534 181837
rect 162858 181037 162914 181837
rect 163778 181037 163834 181837
rect 164698 181037 164754 181837
rect 165618 181037 165674 181837
rect 166538 181037 166594 181837
rect 167458 181037 167514 181837
rect 168378 181037 168434 181837
rect 169298 181037 169354 181837
rect 170218 181037 170274 181837
rect 171138 181037 171194 181837
rect 172058 181037 172114 181837
rect 172978 181037 173034 181837
rect 173898 181037 173954 181837
rect 174818 181037 174874 181837
rect 175738 181037 175794 181837
rect 176658 181037 176714 181837
rect 177578 181037 177634 181837
rect 178498 181037 178554 181837
rect 478 0 534 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 3238 0 3294 800
rect 4158 0 4214 800
rect 5078 0 5134 800
rect 5998 0 6054 800
rect 6918 0 6974 800
rect 7838 0 7894 800
rect 8758 0 8814 800
rect 9678 0 9734 800
rect 10598 0 10654 800
rect 11518 0 11574 800
rect 12438 0 12494 800
rect 13358 0 13414 800
rect 14278 0 14334 800
rect 15198 0 15254 800
rect 16118 0 16174 800
rect 17498 0 17554 800
rect 18418 0 18474 800
rect 19338 0 19394 800
rect 20258 0 20314 800
rect 21178 0 21234 800
rect 22098 0 22154 800
rect 23018 0 23074 800
rect 23938 0 23994 800
rect 24858 0 24914 800
rect 25778 0 25834 800
rect 26698 0 26754 800
rect 27618 0 27674 800
rect 28538 0 28594 800
rect 29458 0 29514 800
rect 30378 0 30434 800
rect 31298 0 31354 800
rect 32218 0 32274 800
rect 33138 0 33194 800
rect 34518 0 34574 800
rect 35438 0 35494 800
rect 36358 0 36414 800
rect 37278 0 37334 800
rect 38198 0 38254 800
rect 39118 0 39174 800
rect 40038 0 40094 800
rect 40958 0 41014 800
rect 41878 0 41934 800
rect 42798 0 42854 800
rect 43718 0 43774 800
rect 44638 0 44694 800
rect 45558 0 45614 800
rect 46478 0 46534 800
rect 47398 0 47454 800
rect 48318 0 48374 800
rect 49238 0 49294 800
rect 50158 0 50214 800
rect 51538 0 51594 800
rect 52458 0 52514 800
rect 53378 0 53434 800
rect 54298 0 54354 800
rect 55218 0 55274 800
rect 56138 0 56194 800
rect 57058 0 57114 800
rect 57978 0 58034 800
rect 58898 0 58954 800
rect 59818 0 59874 800
rect 60738 0 60794 800
rect 61658 0 61714 800
rect 62578 0 62634 800
rect 63498 0 63554 800
rect 64418 0 64474 800
rect 65338 0 65394 800
rect 66258 0 66314 800
rect 67638 0 67694 800
rect 68558 0 68614 800
rect 69478 0 69534 800
rect 70398 0 70454 800
rect 71318 0 71374 800
rect 72238 0 72294 800
rect 73158 0 73214 800
rect 74078 0 74134 800
rect 74998 0 75054 800
rect 75918 0 75974 800
rect 76838 0 76894 800
rect 77758 0 77814 800
rect 78678 0 78734 800
rect 79598 0 79654 800
rect 80518 0 80574 800
rect 81438 0 81494 800
rect 82358 0 82414 800
rect 83278 0 83334 800
rect 84658 0 84714 800
rect 85578 0 85634 800
rect 86498 0 86554 800
rect 87418 0 87474 800
rect 88338 0 88394 800
rect 89258 0 89314 800
rect 90178 0 90234 800
rect 91098 0 91154 800
rect 92018 0 92074 800
rect 92938 0 92994 800
rect 93858 0 93914 800
rect 94778 0 94834 800
rect 95698 0 95754 800
rect 96618 0 96674 800
rect 97538 0 97594 800
rect 98458 0 98514 800
rect 99378 0 99434 800
rect 100298 0 100354 800
rect 101678 0 101734 800
rect 102598 0 102654 800
rect 103518 0 103574 800
rect 104438 0 104494 800
rect 105358 0 105414 800
rect 106278 0 106334 800
rect 107198 0 107254 800
rect 108118 0 108174 800
rect 109038 0 109094 800
rect 109958 0 110014 800
rect 110878 0 110934 800
rect 111798 0 111854 800
rect 112718 0 112774 800
rect 113638 0 113694 800
rect 114558 0 114614 800
rect 115478 0 115534 800
rect 116398 0 116454 800
rect 117778 0 117834 800
rect 118698 0 118754 800
rect 119618 0 119674 800
rect 120538 0 120594 800
rect 121458 0 121514 800
rect 122378 0 122434 800
rect 123298 0 123354 800
rect 124218 0 124274 800
rect 125138 0 125194 800
rect 126058 0 126114 800
rect 126978 0 127034 800
rect 127898 0 127954 800
rect 128818 0 128874 800
rect 129738 0 129794 800
rect 130658 0 130714 800
rect 131578 0 131634 800
rect 132498 0 132554 800
rect 133418 0 133474 800
rect 134798 0 134854 800
rect 135718 0 135774 800
rect 136638 0 136694 800
rect 137558 0 137614 800
rect 138478 0 138534 800
rect 139398 0 139454 800
rect 140318 0 140374 800
rect 141238 0 141294 800
rect 142158 0 142214 800
rect 143078 0 143134 800
rect 143998 0 144054 800
rect 144918 0 144974 800
rect 145838 0 145894 800
rect 146758 0 146814 800
rect 147678 0 147734 800
rect 148598 0 148654 800
rect 149518 0 149574 800
rect 150438 0 150494 800
rect 151818 0 151874 800
rect 152738 0 152794 800
rect 153658 0 153714 800
rect 154578 0 154634 800
rect 155498 0 155554 800
rect 156418 0 156474 800
rect 157338 0 157394 800
rect 158258 0 158314 800
rect 159178 0 159234 800
rect 160098 0 160154 800
rect 161018 0 161074 800
rect 161938 0 161994 800
rect 162858 0 162914 800
rect 163778 0 163834 800
rect 164698 0 164754 800
rect 165618 0 165674 800
rect 166538 0 166594 800
rect 167918 0 167974 800
rect 168838 0 168894 800
rect 169758 0 169814 800
rect 170678 0 170734 800
rect 171598 0 171654 800
rect 172518 0 172574 800
rect 173438 0 173494 800
rect 174358 0 174414 800
rect 175278 0 175334 800
rect 176198 0 176254 800
rect 177118 0 177174 800
rect 178038 0 178094 800
rect 178958 0 179014 800
<< obsm2 >>
rect 1122 180981 1802 181037
rect 1970 180981 2722 181037
rect 2890 180981 3642 181037
rect 3810 180981 4562 181037
rect 4730 180981 5482 181037
rect 5650 180981 6402 181037
rect 6570 180981 7322 181037
rect 7490 180981 8242 181037
rect 8410 180981 9162 181037
rect 9330 180981 10082 181037
rect 10250 180981 11002 181037
rect 11170 180981 12382 181037
rect 12550 180981 13302 181037
rect 13470 180981 14222 181037
rect 14390 180981 15142 181037
rect 15310 180981 16062 181037
rect 16230 180981 16982 181037
rect 17150 180981 17902 181037
rect 18070 180981 18822 181037
rect 18990 180981 19742 181037
rect 19910 180981 20662 181037
rect 20830 180981 21582 181037
rect 21750 180981 22502 181037
rect 22670 180981 23422 181037
rect 23590 180981 24342 181037
rect 24510 180981 25262 181037
rect 25430 180981 26182 181037
rect 26350 180981 27102 181037
rect 27270 180981 28022 181037
rect 28190 180981 29402 181037
rect 29570 180981 30322 181037
rect 30490 180981 31242 181037
rect 31410 180981 32162 181037
rect 32330 180981 33082 181037
rect 33250 180981 34002 181037
rect 34170 180981 34922 181037
rect 35090 180981 35842 181037
rect 36010 180981 36762 181037
rect 36930 180981 37682 181037
rect 37850 180981 38602 181037
rect 38770 180981 39522 181037
rect 39690 180981 40442 181037
rect 40610 180981 41362 181037
rect 41530 180981 42282 181037
rect 42450 180981 43202 181037
rect 43370 180981 44122 181037
rect 44290 180981 45502 181037
rect 45670 180981 46422 181037
rect 46590 180981 47342 181037
rect 47510 180981 48262 181037
rect 48430 180981 49182 181037
rect 49350 180981 50102 181037
rect 50270 180981 51022 181037
rect 51190 180981 51942 181037
rect 52110 180981 52862 181037
rect 53030 180981 53782 181037
rect 53950 180981 54702 181037
rect 54870 180981 55622 181037
rect 55790 180981 56542 181037
rect 56710 180981 57462 181037
rect 57630 180981 58382 181037
rect 58550 180981 59302 181037
rect 59470 180981 60222 181037
rect 60390 180981 61142 181037
rect 61310 180981 62522 181037
rect 62690 180981 63442 181037
rect 63610 180981 64362 181037
rect 64530 180981 65282 181037
rect 65450 180981 66202 181037
rect 66370 180981 67122 181037
rect 67290 180981 68042 181037
rect 68210 180981 68962 181037
rect 69130 180981 69882 181037
rect 70050 180981 70802 181037
rect 70970 180981 71722 181037
rect 71890 180981 72642 181037
rect 72810 180981 73562 181037
rect 73730 180981 74482 181037
rect 74650 180981 75402 181037
rect 75570 180981 76322 181037
rect 76490 180981 77242 181037
rect 77410 180981 78162 181037
rect 78330 180981 79542 181037
rect 79710 180981 80462 181037
rect 80630 180981 81382 181037
rect 81550 180981 82302 181037
rect 82470 180981 83222 181037
rect 83390 180981 84142 181037
rect 84310 180981 85062 181037
rect 85230 180981 85982 181037
rect 86150 180981 86902 181037
rect 87070 180981 87822 181037
rect 87990 180981 88742 181037
rect 88910 180981 89662 181037
rect 89830 180981 90582 181037
rect 90750 180981 91502 181037
rect 91670 180981 92422 181037
rect 92590 180981 93342 181037
rect 93510 180981 94262 181037
rect 94430 180981 95182 181037
rect 95350 180981 96562 181037
rect 96730 180981 97482 181037
rect 97650 180981 98402 181037
rect 98570 180981 99322 181037
rect 99490 180981 100242 181037
rect 100410 180981 101162 181037
rect 101330 180981 102082 181037
rect 102250 180981 103002 181037
rect 103170 180981 103922 181037
rect 104090 180981 104842 181037
rect 105010 180981 105762 181037
rect 105930 180981 106682 181037
rect 106850 180981 107602 181037
rect 107770 180981 108522 181037
rect 108690 180981 109442 181037
rect 109610 180981 110362 181037
rect 110530 180981 111282 181037
rect 111450 180981 112662 181037
rect 112830 180981 113582 181037
rect 113750 180981 114502 181037
rect 114670 180981 115422 181037
rect 115590 180981 116342 181037
rect 116510 180981 117262 181037
rect 117430 180981 118182 181037
rect 118350 180981 119102 181037
rect 119270 180981 120022 181037
rect 120190 180981 120942 181037
rect 121110 180981 121862 181037
rect 122030 180981 122782 181037
rect 122950 180981 123702 181037
rect 123870 180981 124622 181037
rect 124790 180981 125542 181037
rect 125710 180981 126462 181037
rect 126630 180981 127382 181037
rect 127550 180981 128302 181037
rect 128470 180981 129682 181037
rect 129850 180981 130602 181037
rect 130770 180981 131522 181037
rect 131690 180981 132442 181037
rect 132610 180981 133362 181037
rect 133530 180981 134282 181037
rect 134450 180981 135202 181037
rect 135370 180981 136122 181037
rect 136290 180981 137042 181037
rect 137210 180981 137962 181037
rect 138130 180981 138882 181037
rect 139050 180981 139802 181037
rect 139970 180981 140722 181037
rect 140890 180981 141642 181037
rect 141810 180981 142562 181037
rect 142730 180981 143482 181037
rect 143650 180981 144402 181037
rect 144570 180981 145322 181037
rect 145490 180981 146702 181037
rect 146870 180981 147622 181037
rect 147790 180981 148542 181037
rect 148710 180981 149462 181037
rect 149630 180981 150382 181037
rect 150550 180981 151302 181037
rect 151470 180981 152222 181037
rect 152390 180981 153142 181037
rect 153310 180981 154062 181037
rect 154230 180981 154982 181037
rect 155150 180981 155902 181037
rect 156070 180981 156822 181037
rect 156990 180981 157742 181037
rect 157910 180981 158662 181037
rect 158830 180981 159582 181037
rect 159750 180981 160502 181037
rect 160670 180981 161422 181037
rect 161590 180981 162802 181037
rect 162970 180981 163722 181037
rect 163890 180981 164642 181037
rect 164810 180981 165562 181037
rect 165730 180981 166482 181037
rect 166650 180981 167402 181037
rect 167570 180981 168322 181037
rect 168490 180981 169242 181037
rect 169410 180981 170162 181037
rect 170330 180981 171082 181037
rect 171250 180981 172002 181037
rect 172170 180981 172922 181037
rect 173090 180981 173842 181037
rect 174010 180981 174762 181037
rect 174930 180981 175682 181037
rect 175850 180981 176602 181037
rect 176770 180981 177522 181037
rect 177690 180981 178442 181037
rect 178610 180981 179012 181037
rect 1122 856 179012 180981
rect 1122 800 1342 856
rect 1510 800 2262 856
rect 2430 800 3182 856
rect 3350 800 4102 856
rect 4270 800 5022 856
rect 5190 800 5942 856
rect 6110 800 6862 856
rect 7030 800 7782 856
rect 7950 800 8702 856
rect 8870 800 9622 856
rect 9790 800 10542 856
rect 10710 800 11462 856
rect 11630 800 12382 856
rect 12550 800 13302 856
rect 13470 800 14222 856
rect 14390 800 15142 856
rect 15310 800 16062 856
rect 16230 800 17442 856
rect 17610 800 18362 856
rect 18530 800 19282 856
rect 19450 800 20202 856
rect 20370 800 21122 856
rect 21290 800 22042 856
rect 22210 800 22962 856
rect 23130 800 23882 856
rect 24050 800 24802 856
rect 24970 800 25722 856
rect 25890 800 26642 856
rect 26810 800 27562 856
rect 27730 800 28482 856
rect 28650 800 29402 856
rect 29570 800 30322 856
rect 30490 800 31242 856
rect 31410 800 32162 856
rect 32330 800 33082 856
rect 33250 800 34462 856
rect 34630 800 35382 856
rect 35550 800 36302 856
rect 36470 800 37222 856
rect 37390 800 38142 856
rect 38310 800 39062 856
rect 39230 800 39982 856
rect 40150 800 40902 856
rect 41070 800 41822 856
rect 41990 800 42742 856
rect 42910 800 43662 856
rect 43830 800 44582 856
rect 44750 800 45502 856
rect 45670 800 46422 856
rect 46590 800 47342 856
rect 47510 800 48262 856
rect 48430 800 49182 856
rect 49350 800 50102 856
rect 50270 800 51482 856
rect 51650 800 52402 856
rect 52570 800 53322 856
rect 53490 800 54242 856
rect 54410 800 55162 856
rect 55330 800 56082 856
rect 56250 800 57002 856
rect 57170 800 57922 856
rect 58090 800 58842 856
rect 59010 800 59762 856
rect 59930 800 60682 856
rect 60850 800 61602 856
rect 61770 800 62522 856
rect 62690 800 63442 856
rect 63610 800 64362 856
rect 64530 800 65282 856
rect 65450 800 66202 856
rect 66370 800 67582 856
rect 67750 800 68502 856
rect 68670 800 69422 856
rect 69590 800 70342 856
rect 70510 800 71262 856
rect 71430 800 72182 856
rect 72350 800 73102 856
rect 73270 800 74022 856
rect 74190 800 74942 856
rect 75110 800 75862 856
rect 76030 800 76782 856
rect 76950 800 77702 856
rect 77870 800 78622 856
rect 78790 800 79542 856
rect 79710 800 80462 856
rect 80630 800 81382 856
rect 81550 800 82302 856
rect 82470 800 83222 856
rect 83390 800 84602 856
rect 84770 800 85522 856
rect 85690 800 86442 856
rect 86610 800 87362 856
rect 87530 800 88282 856
rect 88450 800 89202 856
rect 89370 800 90122 856
rect 90290 800 91042 856
rect 91210 800 91962 856
rect 92130 800 92882 856
rect 93050 800 93802 856
rect 93970 800 94722 856
rect 94890 800 95642 856
rect 95810 800 96562 856
rect 96730 800 97482 856
rect 97650 800 98402 856
rect 98570 800 99322 856
rect 99490 800 100242 856
rect 100410 800 101622 856
rect 101790 800 102542 856
rect 102710 800 103462 856
rect 103630 800 104382 856
rect 104550 800 105302 856
rect 105470 800 106222 856
rect 106390 800 107142 856
rect 107310 800 108062 856
rect 108230 800 108982 856
rect 109150 800 109902 856
rect 110070 800 110822 856
rect 110990 800 111742 856
rect 111910 800 112662 856
rect 112830 800 113582 856
rect 113750 800 114502 856
rect 114670 800 115422 856
rect 115590 800 116342 856
rect 116510 800 117722 856
rect 117890 800 118642 856
rect 118810 800 119562 856
rect 119730 800 120482 856
rect 120650 800 121402 856
rect 121570 800 122322 856
rect 122490 800 123242 856
rect 123410 800 124162 856
rect 124330 800 125082 856
rect 125250 800 126002 856
rect 126170 800 126922 856
rect 127090 800 127842 856
rect 128010 800 128762 856
rect 128930 800 129682 856
rect 129850 800 130602 856
rect 130770 800 131522 856
rect 131690 800 132442 856
rect 132610 800 133362 856
rect 133530 800 134742 856
rect 134910 800 135662 856
rect 135830 800 136582 856
rect 136750 800 137502 856
rect 137670 800 138422 856
rect 138590 800 139342 856
rect 139510 800 140262 856
rect 140430 800 141182 856
rect 141350 800 142102 856
rect 142270 800 143022 856
rect 143190 800 143942 856
rect 144110 800 144862 856
rect 145030 800 145782 856
rect 145950 800 146702 856
rect 146870 800 147622 856
rect 147790 800 148542 856
rect 148710 800 149462 856
rect 149630 800 150382 856
rect 150550 800 151762 856
rect 151930 800 152682 856
rect 152850 800 153602 856
rect 153770 800 154522 856
rect 154690 800 155442 856
rect 155610 800 156362 856
rect 156530 800 157282 856
rect 157450 800 158202 856
rect 158370 800 159122 856
rect 159290 800 160042 856
rect 160210 800 160962 856
rect 161130 800 161882 856
rect 162050 800 162802 856
rect 162970 800 163722 856
rect 163890 800 164642 856
rect 164810 800 165562 856
rect 165730 800 166482 856
rect 166650 800 167862 856
rect 168030 800 168782 856
rect 168950 800 169702 856
rect 169870 800 170622 856
rect 170790 800 171542 856
rect 171710 800 172462 856
rect 172630 800 173382 856
rect 173550 800 174302 856
rect 174470 800 175222 856
rect 175390 800 176142 856
rect 176310 800 177062 856
rect 177230 800 177982 856
rect 178150 800 178902 856
<< metal3 >>
rect 0 180888 800 181008
rect 178893 180208 179693 180328
rect 0 179528 800 179648
rect 178893 178848 179693 178968
rect 0 178168 800 178288
rect 178893 177488 179693 177608
rect 0 176808 800 176928
rect 178893 176128 179693 176248
rect 0 175448 800 175568
rect 178893 174768 179693 174888
rect 0 174088 800 174208
rect 178893 173408 179693 173528
rect 0 172048 800 172168
rect 178893 172048 179693 172168
rect 0 170688 800 170808
rect 178893 170688 179693 170808
rect 0 169328 800 169448
rect 178893 169328 179693 169448
rect 0 167968 800 168088
rect 178893 167968 179693 168088
rect 0 166608 800 166728
rect 178893 166608 179693 166728
rect 0 165248 800 165368
rect 178893 165248 179693 165368
rect 0 163888 800 164008
rect 178893 163888 179693 164008
rect 0 162528 800 162648
rect 178893 162528 179693 162648
rect 0 161168 800 161288
rect 178893 161168 179693 161288
rect 0 159808 800 159928
rect 178893 159808 179693 159928
rect 0 158448 800 158568
rect 178893 158448 179693 158568
rect 0 157088 800 157208
rect 178893 157088 179693 157208
rect 0 155728 800 155848
rect 178893 155048 179693 155168
rect 0 154368 800 154488
rect 178893 153688 179693 153808
rect 0 153008 800 153128
rect 178893 152328 179693 152448
rect 0 151648 800 151768
rect 178893 150968 179693 151088
rect 0 150288 800 150408
rect 178893 149608 179693 149728
rect 0 148248 800 148368
rect 178893 148248 179693 148368
rect 0 146888 800 147008
rect 178893 146888 179693 147008
rect 0 145528 800 145648
rect 178893 145528 179693 145648
rect 0 144168 800 144288
rect 178893 144168 179693 144288
rect 0 142808 800 142928
rect 178893 142808 179693 142928
rect 0 141448 800 141568
rect 178893 141448 179693 141568
rect 0 140088 800 140208
rect 178893 140088 179693 140208
rect 0 138728 800 138848
rect 178893 138728 179693 138848
rect 0 137368 800 137488
rect 178893 137368 179693 137488
rect 0 136008 800 136128
rect 178893 136008 179693 136128
rect 0 134648 800 134768
rect 178893 134648 179693 134768
rect 0 133288 800 133408
rect 178893 133288 179693 133408
rect 0 131928 800 132048
rect 178893 131248 179693 131368
rect 0 130568 800 130688
rect 178893 129888 179693 130008
rect 0 129208 800 129328
rect 178893 128528 179693 128648
rect 0 127848 800 127968
rect 178893 127168 179693 127288
rect 0 126488 800 126608
rect 178893 125808 179693 125928
rect 0 125128 800 125248
rect 178893 124448 179693 124568
rect 0 123088 800 123208
rect 178893 123088 179693 123208
rect 0 121728 800 121848
rect 178893 121728 179693 121848
rect 0 120368 800 120488
rect 178893 120368 179693 120488
rect 0 119008 800 119128
rect 178893 119008 179693 119128
rect 0 117648 800 117768
rect 178893 117648 179693 117768
rect 0 116288 800 116408
rect 178893 116288 179693 116408
rect 0 114928 800 115048
rect 178893 114928 179693 115048
rect 0 113568 800 113688
rect 178893 113568 179693 113688
rect 0 112208 800 112328
rect 178893 112208 179693 112328
rect 0 110848 800 110968
rect 178893 110848 179693 110968
rect 0 109488 800 109608
rect 178893 109488 179693 109608
rect 0 108128 800 108248
rect 178893 108128 179693 108248
rect 0 106768 800 106888
rect 178893 106088 179693 106208
rect 0 105408 800 105528
rect 178893 104728 179693 104848
rect 0 104048 800 104168
rect 178893 103368 179693 103488
rect 0 102688 800 102808
rect 178893 102008 179693 102128
rect 0 101328 800 101448
rect 178893 100648 179693 100768
rect 0 99968 800 100088
rect 178893 99288 179693 99408
rect 0 97928 800 98048
rect 178893 97928 179693 98048
rect 0 96568 800 96688
rect 178893 96568 179693 96688
rect 0 95208 800 95328
rect 178893 95208 179693 95328
rect 0 93848 800 93968
rect 178893 93848 179693 93968
rect 0 92488 800 92608
rect 178893 92488 179693 92608
rect 0 91128 800 91248
rect 178893 91128 179693 91248
rect 0 89768 800 89888
rect 178893 89768 179693 89888
rect 0 88408 800 88528
rect 178893 88408 179693 88528
rect 0 87048 800 87168
rect 178893 87048 179693 87168
rect 0 85688 800 85808
rect 178893 85688 179693 85808
rect 0 84328 800 84448
rect 178893 84328 179693 84448
rect 0 82968 800 83088
rect 178893 82968 179693 83088
rect 0 81608 800 81728
rect 178893 80928 179693 81048
rect 0 80248 800 80368
rect 178893 79568 179693 79688
rect 0 78888 800 79008
rect 178893 78208 179693 78328
rect 0 77528 800 77648
rect 178893 76848 179693 76968
rect 0 76168 800 76288
rect 178893 75488 179693 75608
rect 0 74128 800 74248
rect 178893 74128 179693 74248
rect 0 72768 800 72888
rect 178893 72768 179693 72888
rect 0 71408 800 71528
rect 178893 71408 179693 71528
rect 0 70048 800 70168
rect 178893 70048 179693 70168
rect 0 68688 800 68808
rect 178893 68688 179693 68808
rect 0 67328 800 67448
rect 178893 67328 179693 67448
rect 0 65968 800 66088
rect 178893 65968 179693 66088
rect 0 64608 800 64728
rect 178893 64608 179693 64728
rect 0 63248 800 63368
rect 178893 63248 179693 63368
rect 0 61888 800 62008
rect 178893 61888 179693 62008
rect 0 60528 800 60648
rect 178893 60528 179693 60648
rect 0 59168 800 59288
rect 178893 59168 179693 59288
rect 0 57808 800 57928
rect 178893 57128 179693 57248
rect 0 56448 800 56568
rect 178893 55768 179693 55888
rect 0 55088 800 55208
rect 178893 54408 179693 54528
rect 0 53728 800 53848
rect 178893 53048 179693 53168
rect 0 52368 800 52488
rect 178893 51688 179693 51808
rect 0 51008 800 51128
rect 178893 50328 179693 50448
rect 0 48968 800 49088
rect 178893 48968 179693 49088
rect 0 47608 800 47728
rect 178893 47608 179693 47728
rect 0 46248 800 46368
rect 178893 46248 179693 46368
rect 0 44888 800 45008
rect 178893 44888 179693 45008
rect 0 43528 800 43648
rect 178893 43528 179693 43648
rect 0 42168 800 42288
rect 178893 42168 179693 42288
rect 0 40808 800 40928
rect 178893 40808 179693 40928
rect 0 39448 800 39568
rect 178893 39448 179693 39568
rect 0 38088 800 38208
rect 178893 38088 179693 38208
rect 0 36728 800 36848
rect 178893 36728 179693 36848
rect 0 35368 800 35488
rect 178893 35368 179693 35488
rect 0 34008 800 34128
rect 178893 34008 179693 34128
rect 0 32648 800 32768
rect 178893 31968 179693 32088
rect 0 31288 800 31408
rect 178893 30608 179693 30728
rect 0 29928 800 30048
rect 178893 29248 179693 29368
rect 0 28568 800 28688
rect 178893 27888 179693 28008
rect 0 27208 800 27328
rect 178893 26528 179693 26648
rect 0 25848 800 25968
rect 178893 25168 179693 25288
rect 0 23808 800 23928
rect 178893 23808 179693 23928
rect 0 22448 800 22568
rect 178893 22448 179693 22568
rect 0 21088 800 21208
rect 178893 21088 179693 21208
rect 0 19728 800 19848
rect 178893 19728 179693 19848
rect 0 18368 800 18488
rect 178893 18368 179693 18488
rect 0 17008 800 17128
rect 178893 17008 179693 17128
rect 0 15648 800 15768
rect 178893 15648 179693 15768
rect 0 14288 800 14408
rect 178893 14288 179693 14408
rect 0 12928 800 13048
rect 178893 12928 179693 13048
rect 0 11568 800 11688
rect 178893 11568 179693 11688
rect 0 10208 800 10328
rect 178893 10208 179693 10328
rect 0 8848 800 8968
rect 178893 8848 179693 8968
rect 0 7488 800 7608
rect 178893 6808 179693 6928
rect 0 6128 800 6248
rect 178893 5448 179693 5568
rect 0 4768 800 4888
rect 178893 4088 179693 4208
rect 0 3408 800 3528
rect 178893 2728 179693 2848
rect 0 2048 800 2168
rect 178893 1368 179693 1488
<< obsm3 >>
rect 800 180128 178813 180301
rect 800 179728 178893 180128
rect 880 179448 178893 179728
rect 800 179048 178893 179448
rect 800 178768 178813 179048
rect 800 178368 178893 178768
rect 880 178088 178893 178368
rect 800 177688 178893 178088
rect 800 177408 178813 177688
rect 800 177008 178893 177408
rect 880 176728 178893 177008
rect 800 176328 178893 176728
rect 800 176048 178813 176328
rect 800 175648 178893 176048
rect 880 175368 178893 175648
rect 800 174968 178893 175368
rect 800 174688 178813 174968
rect 800 174288 178893 174688
rect 880 174008 178893 174288
rect 800 173608 178893 174008
rect 800 173328 178813 173608
rect 800 172248 178893 173328
rect 880 171968 178813 172248
rect 800 170888 178893 171968
rect 880 170608 178813 170888
rect 800 169528 178893 170608
rect 880 169248 178813 169528
rect 800 168168 178893 169248
rect 880 167888 178813 168168
rect 800 166808 178893 167888
rect 880 166528 178813 166808
rect 800 165448 178893 166528
rect 880 165168 178813 165448
rect 800 164088 178893 165168
rect 880 163808 178813 164088
rect 800 162728 178893 163808
rect 880 162448 178813 162728
rect 800 161368 178893 162448
rect 880 161088 178813 161368
rect 800 160008 178893 161088
rect 880 159728 178813 160008
rect 800 158648 178893 159728
rect 880 158368 178813 158648
rect 800 157288 178893 158368
rect 880 157008 178813 157288
rect 800 155928 178893 157008
rect 880 155648 178893 155928
rect 800 155248 178893 155648
rect 800 154968 178813 155248
rect 800 154568 178893 154968
rect 880 154288 178893 154568
rect 800 153888 178893 154288
rect 800 153608 178813 153888
rect 800 153208 178893 153608
rect 880 152928 178893 153208
rect 800 152528 178893 152928
rect 800 152248 178813 152528
rect 800 151848 178893 152248
rect 880 151568 178893 151848
rect 800 151168 178893 151568
rect 800 150888 178813 151168
rect 800 150488 178893 150888
rect 880 150208 178893 150488
rect 800 149808 178893 150208
rect 800 149528 178813 149808
rect 800 148448 178893 149528
rect 880 148168 178813 148448
rect 800 147088 178893 148168
rect 880 146808 178813 147088
rect 800 145728 178893 146808
rect 880 145448 178813 145728
rect 800 144368 178893 145448
rect 880 144088 178813 144368
rect 800 143008 178893 144088
rect 880 142728 178813 143008
rect 800 141648 178893 142728
rect 880 141368 178813 141648
rect 800 140288 178893 141368
rect 880 140008 178813 140288
rect 800 138928 178893 140008
rect 880 138648 178813 138928
rect 800 137568 178893 138648
rect 880 137288 178813 137568
rect 800 136208 178893 137288
rect 880 135928 178813 136208
rect 800 134848 178893 135928
rect 880 134568 178813 134848
rect 800 133488 178893 134568
rect 880 133208 178813 133488
rect 800 132128 178893 133208
rect 880 131848 178893 132128
rect 800 131448 178893 131848
rect 800 131168 178813 131448
rect 800 130768 178893 131168
rect 880 130488 178893 130768
rect 800 130088 178893 130488
rect 800 129808 178813 130088
rect 800 129408 178893 129808
rect 880 129128 178893 129408
rect 800 128728 178893 129128
rect 800 128448 178813 128728
rect 800 128048 178893 128448
rect 880 127768 178893 128048
rect 800 127368 178893 127768
rect 800 127088 178813 127368
rect 800 126688 178893 127088
rect 880 126408 178893 126688
rect 800 126008 178893 126408
rect 800 125728 178813 126008
rect 800 125328 178893 125728
rect 880 125048 178893 125328
rect 800 124648 178893 125048
rect 800 124368 178813 124648
rect 800 123288 178893 124368
rect 880 123008 178813 123288
rect 800 121928 178893 123008
rect 880 121648 178813 121928
rect 800 120568 178893 121648
rect 880 120288 178813 120568
rect 800 119208 178893 120288
rect 880 118928 178813 119208
rect 800 117848 178893 118928
rect 880 117568 178813 117848
rect 800 116488 178893 117568
rect 880 116208 178813 116488
rect 800 115128 178893 116208
rect 880 114848 178813 115128
rect 800 113768 178893 114848
rect 880 113488 178813 113768
rect 800 112408 178893 113488
rect 880 112128 178813 112408
rect 800 111048 178893 112128
rect 880 110768 178813 111048
rect 800 109688 178893 110768
rect 880 109408 178813 109688
rect 800 108328 178893 109408
rect 880 108048 178813 108328
rect 800 106968 178893 108048
rect 880 106688 178893 106968
rect 800 106288 178893 106688
rect 800 106008 178813 106288
rect 800 105608 178893 106008
rect 880 105328 178893 105608
rect 800 104928 178893 105328
rect 800 104648 178813 104928
rect 800 104248 178893 104648
rect 880 103968 178893 104248
rect 800 103568 178893 103968
rect 800 103288 178813 103568
rect 800 102888 178893 103288
rect 880 102608 178893 102888
rect 800 102208 178893 102608
rect 800 101928 178813 102208
rect 800 101528 178893 101928
rect 880 101248 178893 101528
rect 800 100848 178893 101248
rect 800 100568 178813 100848
rect 800 100168 178893 100568
rect 880 99888 178893 100168
rect 800 99488 178893 99888
rect 800 99208 178813 99488
rect 800 98128 178893 99208
rect 880 97848 178813 98128
rect 800 96768 178893 97848
rect 880 96488 178813 96768
rect 800 95408 178893 96488
rect 880 95128 178813 95408
rect 800 94048 178893 95128
rect 880 93768 178813 94048
rect 800 92688 178893 93768
rect 880 92408 178813 92688
rect 800 91328 178893 92408
rect 880 91048 178813 91328
rect 800 89968 178893 91048
rect 880 89688 178813 89968
rect 800 88608 178893 89688
rect 880 88328 178813 88608
rect 800 87248 178893 88328
rect 880 86968 178813 87248
rect 800 85888 178893 86968
rect 880 85608 178813 85888
rect 800 84528 178893 85608
rect 880 84248 178813 84528
rect 800 83168 178893 84248
rect 880 82888 178813 83168
rect 800 81808 178893 82888
rect 880 81528 178893 81808
rect 800 81128 178893 81528
rect 800 80848 178813 81128
rect 800 80448 178893 80848
rect 880 80168 178893 80448
rect 800 79768 178893 80168
rect 800 79488 178813 79768
rect 800 79088 178893 79488
rect 880 78808 178893 79088
rect 800 78408 178893 78808
rect 800 78128 178813 78408
rect 800 77728 178893 78128
rect 880 77448 178893 77728
rect 800 77048 178893 77448
rect 800 76768 178813 77048
rect 800 76368 178893 76768
rect 880 76088 178893 76368
rect 800 75688 178893 76088
rect 800 75408 178813 75688
rect 800 74328 178893 75408
rect 880 74048 178813 74328
rect 800 72968 178893 74048
rect 880 72688 178813 72968
rect 800 71608 178893 72688
rect 880 71328 178813 71608
rect 800 70248 178893 71328
rect 880 69968 178813 70248
rect 800 68888 178893 69968
rect 880 68608 178813 68888
rect 800 67528 178893 68608
rect 880 67248 178813 67528
rect 800 66168 178893 67248
rect 880 65888 178813 66168
rect 800 64808 178893 65888
rect 880 64528 178813 64808
rect 800 63448 178893 64528
rect 880 63168 178813 63448
rect 800 62088 178893 63168
rect 880 61808 178813 62088
rect 800 60728 178893 61808
rect 880 60448 178813 60728
rect 800 59368 178893 60448
rect 880 59088 178813 59368
rect 800 58008 178893 59088
rect 880 57728 178893 58008
rect 800 57328 178893 57728
rect 800 57048 178813 57328
rect 800 56648 178893 57048
rect 880 56368 178893 56648
rect 800 55968 178893 56368
rect 800 55688 178813 55968
rect 800 55288 178893 55688
rect 880 55008 178893 55288
rect 800 54608 178893 55008
rect 800 54328 178813 54608
rect 800 53928 178893 54328
rect 880 53648 178893 53928
rect 800 53248 178893 53648
rect 800 52968 178813 53248
rect 800 52568 178893 52968
rect 880 52288 178893 52568
rect 800 51888 178893 52288
rect 800 51608 178813 51888
rect 800 51208 178893 51608
rect 880 50928 178893 51208
rect 800 50528 178893 50928
rect 800 50248 178813 50528
rect 800 49168 178893 50248
rect 880 48888 178813 49168
rect 800 47808 178893 48888
rect 880 47528 178813 47808
rect 800 46448 178893 47528
rect 880 46168 178813 46448
rect 800 45088 178893 46168
rect 880 44808 178813 45088
rect 800 43728 178893 44808
rect 880 43448 178813 43728
rect 800 42368 178893 43448
rect 880 42088 178813 42368
rect 800 41008 178893 42088
rect 880 40728 178813 41008
rect 800 39648 178893 40728
rect 880 39368 178813 39648
rect 800 38288 178893 39368
rect 880 38008 178813 38288
rect 800 36928 178893 38008
rect 880 36648 178813 36928
rect 800 35568 178893 36648
rect 880 35288 178813 35568
rect 800 34208 178893 35288
rect 880 33928 178813 34208
rect 800 32848 178893 33928
rect 880 32568 178893 32848
rect 800 32168 178893 32568
rect 800 31888 178813 32168
rect 800 31488 178893 31888
rect 880 31208 178893 31488
rect 800 30808 178893 31208
rect 800 30528 178813 30808
rect 800 30128 178893 30528
rect 880 29848 178893 30128
rect 800 29448 178893 29848
rect 800 29168 178813 29448
rect 800 28768 178893 29168
rect 880 28488 178893 28768
rect 800 28088 178893 28488
rect 800 27808 178813 28088
rect 800 27408 178893 27808
rect 880 27128 178893 27408
rect 800 26728 178893 27128
rect 800 26448 178813 26728
rect 800 26048 178893 26448
rect 880 25768 178893 26048
rect 800 25368 178893 25768
rect 800 25088 178813 25368
rect 800 24008 178893 25088
rect 880 23728 178813 24008
rect 800 22648 178893 23728
rect 880 22368 178813 22648
rect 800 21288 178893 22368
rect 880 21008 178813 21288
rect 800 19928 178893 21008
rect 880 19648 178813 19928
rect 800 18568 178893 19648
rect 880 18288 178813 18568
rect 800 17208 178893 18288
rect 880 16928 178813 17208
rect 800 15848 178893 16928
rect 880 15568 178813 15848
rect 800 14488 178893 15568
rect 880 14208 178813 14488
rect 800 13128 178893 14208
rect 880 12848 178813 13128
rect 800 11768 178893 12848
rect 880 11488 178813 11768
rect 800 10408 178893 11488
rect 880 10128 178813 10408
rect 800 9048 178893 10128
rect 880 8768 178813 9048
rect 800 7688 178893 8768
rect 880 7408 178893 7688
rect 800 7008 178893 7408
rect 800 6728 178813 7008
rect 800 6328 178893 6728
rect 880 6048 178893 6328
rect 800 5648 178893 6048
rect 800 5368 178813 5648
rect 800 4968 178893 5368
rect 880 4688 178893 4968
rect 800 4288 178893 4688
rect 800 4008 178813 4288
rect 800 3608 178893 4008
rect 880 3328 178893 3608
rect 800 2928 178893 3328
rect 800 2648 178813 2928
rect 800 2248 178893 2648
rect 880 1968 178893 2248
rect 800 1568 178893 1968
rect 800 1395 178813 1568
<< metal4 >>
rect -8576 -7504 -7976 189200
rect -7636 -6564 -7036 188260
rect -6696 -5624 -6096 187320
rect -5756 -4684 -5156 186380
rect -4816 -3744 -4216 185440
rect -3876 -2804 -3276 184500
rect -2936 -1864 -2336 183560
rect -1996 -924 -1396 182620
rect 804 -1864 1404 183560
rect 4404 -3744 5004 185440
rect 8004 -5624 8604 187320
rect 11604 -7504 12204 189200
rect 18804 -1864 19404 183560
rect 22404 -3744 23004 185440
rect 26004 -5624 26604 187320
rect 29604 -7504 30204 189200
rect 36804 -1864 37404 183560
rect 40404 -3744 41004 185440
rect 44004 -5624 44604 187320
rect 47604 -7504 48204 189200
rect 54804 -1864 55404 183560
rect 58404 -3744 59004 185440
rect 62004 -5624 62604 187320
rect 65604 -7504 66204 189200
rect 72804 -1864 73404 183560
rect 76404 -3744 77004 185440
rect 80004 -5624 80604 187320
rect 83604 -7504 84204 189200
rect 90804 -1864 91404 183560
rect 94404 -3744 95004 185440
rect 98004 -5624 98604 187320
rect 101604 -7504 102204 189200
rect 108804 -1864 109404 183560
rect 112404 -3744 113004 185440
rect 116004 -5624 116604 187320
rect 119604 -7504 120204 189200
rect 126804 -1864 127404 183560
rect 130404 -3744 131004 185440
rect 134004 -5624 134604 187320
rect 137604 -7504 138204 189200
rect 144804 -1864 145404 183560
rect 148404 -3744 149004 185440
rect 152004 -5624 152604 187320
rect 155604 -7504 156204 189200
rect 162804 -1864 163404 183560
rect 166404 -3744 167004 185440
rect 170004 -5624 170604 187320
rect 173604 -7504 174204 189200
rect 181072 -924 181672 182620
rect 182012 -1864 182612 183560
rect 182952 -2804 183552 184500
rect 183892 -3744 184492 185440
rect 184832 -4684 185432 186380
rect 185772 -5624 186372 187320
rect 186712 -6564 187312 188260
rect 187652 -7504 188252 189200
<< obsm4 >>
rect 3371 3027 4324 177989
rect 5084 3027 7924 177989
rect 8684 3027 11524 177989
rect 12284 3027 18724 177989
rect 19484 3027 22324 177989
rect 23084 3027 25924 177989
rect 26684 3027 29524 177989
rect 30284 3027 36724 177989
rect 37484 3027 40324 177989
rect 41084 3027 43924 177989
rect 44684 3027 47524 177989
rect 48284 3027 54724 177989
rect 55484 3027 58324 177989
rect 59084 3027 61924 177989
rect 62684 3027 65524 177989
rect 66284 3027 72724 177989
rect 73484 3027 76324 177989
rect 77084 3027 79924 177989
rect 80684 3027 83524 177989
rect 84284 3027 90724 177989
rect 91484 3027 94324 177989
rect 95084 3027 97924 177989
rect 98684 3027 101524 177989
rect 102284 3027 108724 177989
rect 109484 3027 112324 177989
rect 113084 3027 115924 177989
rect 116684 3027 119524 177989
rect 120284 3027 126724 177989
rect 127484 3027 130324 177989
rect 131084 3027 133924 177989
rect 134684 3027 137524 177989
rect 138284 3027 144724 177989
rect 145484 3027 148324 177989
rect 149084 3027 151924 177989
rect 152684 3027 155524 177989
rect 156284 3027 162724 177989
rect 163484 3027 165357 177989
<< metal5 >>
rect -8576 188600 188252 189200
rect -7636 187660 187312 188260
rect -6696 186720 186372 187320
rect -5756 185780 185432 186380
rect -4816 184840 184492 185440
rect -3876 183900 183552 184500
rect -2936 182960 182612 183560
rect -1996 182020 181672 182620
rect -8576 174676 188252 175276
rect -6696 171076 186372 171676
rect -4816 167476 184492 168076
rect -2936 163828 182612 164428
rect -8576 156676 188252 157276
rect -6696 153076 186372 153676
rect -4816 149476 184492 150076
rect -2936 145828 182612 146428
rect -8576 138676 188252 139276
rect -6696 135076 186372 135676
rect -4816 131476 184492 132076
rect -2936 127828 182612 128428
rect -8576 120676 188252 121276
rect -6696 117076 186372 117676
rect -4816 113476 184492 114076
rect -2936 109828 182612 110428
rect -8576 102676 188252 103276
rect -6696 99076 186372 99676
rect -4816 95476 184492 96076
rect -2936 91828 182612 92428
rect -8576 84676 188252 85276
rect -6696 81076 186372 81676
rect -4816 77476 184492 78076
rect -2936 73828 182612 74428
rect -8576 66676 188252 67276
rect -6696 63076 186372 63676
rect -4816 59476 184492 60076
rect -2936 55828 182612 56428
rect -8576 48676 188252 49276
rect -6696 45076 186372 45676
rect -4816 41476 184492 42076
rect -2936 37828 182612 38428
rect -8576 30676 188252 31276
rect -6696 27076 186372 27676
rect -4816 23476 184492 24076
rect -2936 19828 182612 20428
rect -8576 12676 188252 13276
rect -6696 9076 186372 9676
rect -4816 5476 184492 6076
rect -2936 1828 182612 2428
rect -1996 -924 181672 -324
rect -2936 -1864 182612 -1264
rect -3876 -2804 183552 -2204
rect -4816 -3744 184492 -3144
rect -5756 -4684 185432 -4084
rect -6696 -5624 186372 -5024
rect -7636 -6564 187312 -5964
rect -8576 -7504 188252 -6904
<< obsm5 >>
rect -8576 189200 -7976 189202
rect 29604 189200 30204 189202
rect 65604 189200 66204 189202
rect 101604 189200 102204 189202
rect 137604 189200 138204 189202
rect 173604 189200 174204 189202
rect 187652 189200 188252 189202
rect -8576 188598 -7976 188600
rect 29604 188598 30204 188600
rect 65604 188598 66204 188600
rect 101604 188598 102204 188600
rect 137604 188598 138204 188600
rect 173604 188598 174204 188600
rect 187652 188598 188252 188600
rect -7636 188260 -7036 188262
rect 11604 188260 12204 188262
rect 47604 188260 48204 188262
rect 83604 188260 84204 188262
rect 119604 188260 120204 188262
rect 155604 188260 156204 188262
rect 186712 188260 187312 188262
rect -7636 187658 -7036 187660
rect 11604 187658 12204 187660
rect 47604 187658 48204 187660
rect 83604 187658 84204 187660
rect 119604 187658 120204 187660
rect 155604 187658 156204 187660
rect 186712 187658 187312 187660
rect -6696 187320 -6096 187322
rect 26004 187320 26604 187322
rect 62004 187320 62604 187322
rect 98004 187320 98604 187322
rect 134004 187320 134604 187322
rect 170004 187320 170604 187322
rect 185772 187320 186372 187322
rect -6696 186718 -6096 186720
rect 26004 186718 26604 186720
rect 62004 186718 62604 186720
rect 98004 186718 98604 186720
rect 134004 186718 134604 186720
rect 170004 186718 170604 186720
rect 185772 186718 186372 186720
rect -5756 186380 -5156 186382
rect 8004 186380 8604 186382
rect 44004 186380 44604 186382
rect 80004 186380 80604 186382
rect 116004 186380 116604 186382
rect 152004 186380 152604 186382
rect 184832 186380 185432 186382
rect -5756 185778 -5156 185780
rect 8004 185778 8604 185780
rect 44004 185778 44604 185780
rect 80004 185778 80604 185780
rect 116004 185778 116604 185780
rect 152004 185778 152604 185780
rect 184832 185778 185432 185780
rect -4816 185440 -4216 185442
rect 22404 185440 23004 185442
rect 58404 185440 59004 185442
rect 94404 185440 95004 185442
rect 130404 185440 131004 185442
rect 166404 185440 167004 185442
rect 183892 185440 184492 185442
rect -4816 184838 -4216 184840
rect 22404 184838 23004 184840
rect 58404 184838 59004 184840
rect 94404 184838 95004 184840
rect 130404 184838 131004 184840
rect 166404 184838 167004 184840
rect 183892 184838 184492 184840
rect -3876 184500 -3276 184502
rect 4404 184500 5004 184502
rect 40404 184500 41004 184502
rect 76404 184500 77004 184502
rect 112404 184500 113004 184502
rect 148404 184500 149004 184502
rect 182952 184500 183552 184502
rect -3876 183898 -3276 183900
rect 4404 183898 5004 183900
rect 40404 183898 41004 183900
rect 76404 183898 77004 183900
rect 112404 183898 113004 183900
rect 148404 183898 149004 183900
rect 182952 183898 183552 183900
rect -2936 183560 -2336 183562
rect 18804 183560 19404 183562
rect 54804 183560 55404 183562
rect 90804 183560 91404 183562
rect 126804 183560 127404 183562
rect 162804 183560 163404 183562
rect 182012 183560 182612 183562
rect -2936 182958 -2336 182960
rect 18804 182958 19404 182960
rect 54804 182958 55404 182960
rect 90804 182958 91404 182960
rect 126804 182958 127404 182960
rect 162804 182958 163404 182960
rect 182012 182958 182612 182960
rect -1996 182620 -1396 182622
rect 804 182620 1404 182622
rect 36804 182620 37404 182622
rect 72804 182620 73404 182622
rect 108804 182620 109404 182622
rect 144804 182620 145404 182622
rect 181072 182620 181672 182622
rect -1996 182018 -1396 182020
rect 804 182018 1404 182020
rect 36804 182018 37404 182020
rect 72804 182018 73404 182020
rect 108804 182018 109404 182020
rect 144804 182018 145404 182020
rect 181072 182018 181672 182020
rect 0 175596 179693 181700
rect -8576 175276 -7976 175278
rect 187652 175276 188252 175278
rect -8576 174674 -7976 174676
rect 187652 174674 188252 174676
rect 0 171996 179693 174356
rect -6696 171676 -6096 171678
rect 185772 171676 186372 171678
rect -6696 171074 -6096 171076
rect 185772 171074 186372 171076
rect 0 168396 179693 170756
rect -4816 168076 -4216 168078
rect 183892 168076 184492 168078
rect -4816 167474 -4216 167476
rect 183892 167474 184492 167476
rect 0 164748 179693 167156
rect -2936 164428 -2336 164430
rect 182012 164428 182612 164430
rect -2936 163826 -2336 163828
rect 182012 163826 182612 163828
rect 0 157596 179693 163508
rect -7636 157276 -7036 157278
rect 186712 157276 187312 157278
rect -7636 156674 -7036 156676
rect 186712 156674 187312 156676
rect 0 153996 179693 156356
rect -5756 153676 -5156 153678
rect 184832 153676 185432 153678
rect -5756 153074 -5156 153076
rect 184832 153074 185432 153076
rect 0 150396 179693 152756
rect -3876 150076 -3276 150078
rect 182952 150076 183552 150078
rect -3876 149474 -3276 149476
rect 182952 149474 183552 149476
rect 0 146748 179693 149156
rect -1996 146428 -1396 146430
rect 181072 146428 181672 146430
rect -1996 145826 -1396 145828
rect 181072 145826 181672 145828
rect 0 139596 179693 145508
rect -8576 139276 -7976 139278
rect 187652 139276 188252 139278
rect -8576 138674 -7976 138676
rect 187652 138674 188252 138676
rect 0 135996 179693 138356
rect -6696 135676 -6096 135678
rect 185772 135676 186372 135678
rect -6696 135074 -6096 135076
rect 185772 135074 186372 135076
rect 0 132396 179693 134756
rect -4816 132076 -4216 132078
rect 183892 132076 184492 132078
rect -4816 131474 -4216 131476
rect 183892 131474 184492 131476
rect 0 128748 179693 131156
rect -2936 128428 -2336 128430
rect 182012 128428 182612 128430
rect -2936 127826 -2336 127828
rect 182012 127826 182612 127828
rect 0 121596 179693 127508
rect -7636 121276 -7036 121278
rect 186712 121276 187312 121278
rect -7636 120674 -7036 120676
rect 186712 120674 187312 120676
rect 0 117996 179693 120356
rect -5756 117676 -5156 117678
rect 184832 117676 185432 117678
rect -5756 117074 -5156 117076
rect 184832 117074 185432 117076
rect 0 114396 179693 116756
rect -3876 114076 -3276 114078
rect 182952 114076 183552 114078
rect -3876 113474 -3276 113476
rect 182952 113474 183552 113476
rect 0 110748 179693 113156
rect -1996 110428 -1396 110430
rect 181072 110428 181672 110430
rect -1996 109826 -1396 109828
rect 181072 109826 181672 109828
rect 0 103596 179693 109508
rect -8576 103276 -7976 103278
rect 187652 103276 188252 103278
rect -8576 102674 -7976 102676
rect 187652 102674 188252 102676
rect 0 99996 179693 102356
rect -6696 99676 -6096 99678
rect 185772 99676 186372 99678
rect -6696 99074 -6096 99076
rect 185772 99074 186372 99076
rect 0 96396 179693 98756
rect -4816 96076 -4216 96078
rect 183892 96076 184492 96078
rect -4816 95474 -4216 95476
rect 183892 95474 184492 95476
rect 0 92748 179693 95156
rect -2936 92428 -2336 92430
rect 182012 92428 182612 92430
rect -2936 91826 -2336 91828
rect 182012 91826 182612 91828
rect 0 85596 179693 91508
rect -7636 85276 -7036 85278
rect 186712 85276 187312 85278
rect -7636 84674 -7036 84676
rect 186712 84674 187312 84676
rect 0 81996 179693 84356
rect -5756 81676 -5156 81678
rect 184832 81676 185432 81678
rect -5756 81074 -5156 81076
rect 184832 81074 185432 81076
rect 0 78396 179693 80756
rect -3876 78076 -3276 78078
rect 182952 78076 183552 78078
rect -3876 77474 -3276 77476
rect 182952 77474 183552 77476
rect 0 74748 179693 77156
rect -1996 74428 -1396 74430
rect 181072 74428 181672 74430
rect -1996 73826 -1396 73828
rect 181072 73826 181672 73828
rect 0 67596 179693 73508
rect -8576 67276 -7976 67278
rect 187652 67276 188252 67278
rect -8576 66674 -7976 66676
rect 187652 66674 188252 66676
rect 0 63996 179693 66356
rect -6696 63676 -6096 63678
rect 185772 63676 186372 63678
rect -6696 63074 -6096 63076
rect 185772 63074 186372 63076
rect 0 60396 179693 62756
rect -4816 60076 -4216 60078
rect 183892 60076 184492 60078
rect -4816 59474 -4216 59476
rect 183892 59474 184492 59476
rect 0 56748 179693 59156
rect -2936 56428 -2336 56430
rect 182012 56428 182612 56430
rect -2936 55826 -2336 55828
rect 182012 55826 182612 55828
rect 0 49596 179693 55508
rect -7636 49276 -7036 49278
rect 186712 49276 187312 49278
rect -7636 48674 -7036 48676
rect 186712 48674 187312 48676
rect 0 45996 179693 48356
rect -5756 45676 -5156 45678
rect 184832 45676 185432 45678
rect -5756 45074 -5156 45076
rect 184832 45074 185432 45076
rect 0 42396 179693 44756
rect -3876 42076 -3276 42078
rect 182952 42076 183552 42078
rect -3876 41474 -3276 41476
rect 182952 41474 183552 41476
rect 0 38748 179693 41156
rect -1996 38428 -1396 38430
rect 181072 38428 181672 38430
rect -1996 37826 -1396 37828
rect 181072 37826 181672 37828
rect 0 31596 179693 37508
rect -8576 31276 -7976 31278
rect 187652 31276 188252 31278
rect -8576 30674 -7976 30676
rect 187652 30674 188252 30676
rect 0 27996 179693 30356
rect -6696 27676 -6096 27678
rect 185772 27676 186372 27678
rect -6696 27074 -6096 27076
rect 185772 27074 186372 27076
rect 0 24396 179693 26756
rect -4816 24076 -4216 24078
rect 183892 24076 184492 24078
rect -4816 23474 -4216 23476
rect 183892 23474 184492 23476
rect 0 20748 179693 23156
rect -2936 20428 -2336 20430
rect 182012 20428 182612 20430
rect -2936 19826 -2336 19828
rect 182012 19826 182612 19828
rect 0 13596 179693 19508
rect -7636 13276 -7036 13278
rect 186712 13276 187312 13278
rect -7636 12674 -7036 12676
rect 186712 12674 187312 12676
rect 0 9996 179693 12356
rect -5756 9676 -5156 9678
rect 184832 9676 185432 9678
rect -5756 9074 -5156 9076
rect 184832 9074 185432 9076
rect 0 6396 179693 8756
rect -3876 6076 -3276 6078
rect 182952 6076 183552 6078
rect -3876 5474 -3276 5476
rect 182952 5474 183552 5476
rect 0 2748 179693 5156
rect -1996 2428 -1396 2430
rect 181072 2428 181672 2430
rect -1996 1826 -1396 1828
rect 181072 1826 181672 1828
rect 0 0 179693 1508
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 181072 -324 181672 -322
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 181072 -926 181672 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 182012 -1264 182612 -1262
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 182012 -1866 182612 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 182952 -2204 183552 -2202
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 182952 -2806 183552 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 183892 -3144 184492 -3142
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 183892 -3746 184492 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 184832 -4084 185432 -4082
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 184832 -4686 185432 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 185772 -5024 186372 -5022
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 185772 -5626 186372 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 186712 -5964 187312 -5962
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 186712 -6566 187312 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 187652 -6904 188252 -6902
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 187652 -7506 188252 -7504
<< labels >>
rlabel metal2 s 4618 181037 4674 181837 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 178893 140088 179693 140208 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 139398 0 139454 800 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal3 s 0 174088 800 174208 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal3 s 178893 142808 179693 142928 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 160098 0 160154 800 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal3 s 0 130568 800 130688 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 8758 0 8814 800 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 122378 0 122434 800 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal2 s 96618 0 96674 800 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 108578 181037 108634 181837 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal2 s 168838 0 168894 800 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 0 2048 800 2168 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal2 s 106278 0 106334 800 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 178893 74128 179693 74248 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 118238 181037 118294 181837 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal2 s 109958 0 110014 800 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal2 s 134338 181037 134394 181837 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal2 s 10598 0 10654 800 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 0 59168 800 59288 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 178893 117648 179693 117768 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 0 78888 800 79008 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 178893 167968 179693 168088 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal2 s 113638 0 113694 800 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 0 175448 800 175568 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal2 s 51538 0 51594 800 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal2 s 85578 0 85634 800 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 145378 181037 145434 181837 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal3 s 178893 93848 179693 93968 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal2 s 161938 0 161994 800 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 io_in[10]
port 31 nsew signal input
rlabel metal2 s 167458 181037 167514 181837 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 io_in[12]
port 33 nsew signal input
rlabel metal2 s 62578 181037 62634 181837 6 io_in[13]
port 34 nsew signal input
rlabel metal2 s 32218 181037 32274 181837 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 io_in[15]
port 36 nsew signal input
rlabel metal3 s 0 114928 800 115048 6 io_in[16]
port 37 nsew signal input
rlabel metal3 s 178893 106088 179693 106208 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 160558 181037 160614 181837 6 io_in[18]
port 39 nsew signal input
rlabel metal3 s 178893 2728 179693 2848 6 io_in[19]
port 40 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 104898 181037 104954 181837 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 110418 181037 110474 181837 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 68098 181037 68154 181837 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s 0 113568 800 113688 6 io_in[24]
port 46 nsew signal input
rlabel metal3 s 178893 85688 179693 85808 6 io_in[25]
port 47 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 io_in[26]
port 48 nsew signal input
rlabel metal2 s 46478 181037 46534 181837 6 io_in[27]
port 49 nsew signal input
rlabel metal2 s 47398 181037 47454 181837 6 io_in[28]
port 50 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 io_in[29]
port 51 nsew signal input
rlabel metal2 s 149518 181037 149574 181837 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s 178893 15648 179693 15768 6 io_in[30]
port 53 nsew signal input
rlabel metal3 s 178893 10208 179693 10328 6 io_in[31]
port 54 nsew signal input
rlabel metal2 s 14278 181037 14334 181837 6 io_in[32]
port 55 nsew signal input
rlabel metal3 s 0 180888 800 181008 6 io_in[33]
port 56 nsew signal input
rlabel metal3 s 178893 134648 179693 134768 6 io_in[34]
port 57 nsew signal input
rlabel metal2 s 175278 0 175334 800 6 io_in[35]
port 58 nsew signal input
rlabel metal2 s 84198 181037 84254 181837 6 io_in[36]
port 59 nsew signal input
rlabel metal2 s 23478 181037 23534 181837 6 io_in[37]
port 60 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 io_in[3]
port 61 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 178893 29248 179693 29368 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 0 151648 800 151768 6 io_in[6]
port 64 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 io_in[7]
port 65 nsew signal input
rlabel metal2 s 168378 181037 168434 181837 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 178893 161168 179693 161288 6 io_in[9]
port 67 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 io_oeb[0]
port 68 nsew signal output
rlabel metal2 s 165618 0 165674 800 6 io_oeb[10]
port 69 nsew signal output
rlabel metal2 s 148598 0 148654 800 6 io_oeb[11]
port 70 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 io_oeb[12]
port 71 nsew signal output
rlabel metal2 s 59358 181037 59414 181837 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 178893 103368 179693 103488 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 156878 181037 156934 181837 6 io_oeb[15]
port 74 nsew signal output
rlabel metal3 s 178893 40808 179693 40928 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 164698 181037 164754 181837 6 io_oeb[18]
port 77 nsew signal output
rlabel metal3 s 178893 67328 179693 67448 6 io_oeb[19]
port 78 nsew signal output
rlabel metal2 s 131578 0 131634 800 6 io_oeb[1]
port 79 nsew signal output
rlabel metal3 s 178893 109488 179693 109608 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 15198 181037 15254 181837 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 156418 0 156474 800 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s 178893 30608 179693 30728 6 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s 0 170688 800 170808 6 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 io_oeb[26]
port 86 nsew signal output
rlabel metal2 s 81438 181037 81494 181837 6 io_oeb[27]
port 87 nsew signal output
rlabel metal2 s 36818 181037 36874 181837 6 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 io_oeb[29]
port 89 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s 0 137368 800 137488 6 io_oeb[30]
port 91 nsew signal output
rlabel metal2 s 37278 0 37334 800 6 io_oeb[31]
port 92 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s 178893 25168 179693 25288 6 io_oeb[33]
port 94 nsew signal output
rlabel metal2 s 52918 181037 52974 181837 6 io_oeb[34]
port 95 nsew signal output
rlabel metal2 s 73158 0 73214 800 6 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 io_oeb[36]
port 97 nsew signal output
rlabel metal2 s 24398 181037 24454 181837 6 io_oeb[37]
port 98 nsew signal output
rlabel metal2 s 178958 0 179014 800 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 io_oeb[4]
port 100 nsew signal output
rlabel metal2 s 154578 0 154634 800 6 io_oeb[5]
port 101 nsew signal output
rlabel metal2 s 63498 0 63554 800 6 io_oeb[6]
port 102 nsew signal output
rlabel metal2 s 38658 181037 38714 181837 6 io_oeb[7]
port 103 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 io_oeb[8]
port 104 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 io_oeb[9]
port 105 nsew signal output
rlabel metal2 s 82358 181037 82414 181837 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 io_out[10]
port 107 nsew signal output
rlabel metal2 s 89258 0 89314 800 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 178893 110848 179693 110968 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 0 108128 800 108248 6 io_out[13]
port 110 nsew signal output
rlabel metal2 s 105358 0 105414 800 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 157798 181037 157854 181837 6 io_out[15]
port 112 nsew signal output
rlabel metal3 s 178893 173408 179693 173528 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 10138 181037 10194 181837 6 io_out[17]
port 114 nsew signal output
rlabel metal3 s 178893 26528 179693 26648 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 0 157088 800 157208 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 120998 181037 121054 181837 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 79598 181037 79654 181837 6 io_out[21]
port 119 nsew signal output
rlabel metal3 s 0 131928 800 132048 6 io_out[22]
port 120 nsew signal output
rlabel metal3 s 0 71408 800 71528 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s 178893 155048 179693 155168 6 io_out[24]
port 122 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 io_out[25]
port 123 nsew signal output
rlabel metal2 s 76838 0 76894 800 6 io_out[26]
port 124 nsew signal output
rlabel metal2 s 163778 181037 163834 181837 6 io_out[27]
port 125 nsew signal output
rlabel metal2 s 153658 0 153714 800 6 io_out[28]
port 126 nsew signal output
rlabel metal2 s 108118 0 108174 800 6 io_out[29]
port 127 nsew signal output
rlabel metal2 s 126058 0 126114 800 6 io_out[2]
port 128 nsew signal output
rlabel metal2 s 63498 181037 63554 181837 6 io_out[30]
port 129 nsew signal output
rlabel metal3 s 178893 108128 179693 108248 6 io_out[31]
port 130 nsew signal output
rlabel metal3 s 0 142808 800 142928 6 io_out[32]
port 131 nsew signal output
rlabel metal2 s 69938 181037 69994 181837 6 io_out[33]
port 132 nsew signal output
rlabel metal2 s 3698 181037 3754 181837 6 io_out[34]
port 133 nsew signal output
rlabel metal3 s 178893 80928 179693 81048 6 io_out[35]
port 134 nsew signal output
rlabel metal2 s 12438 181037 12494 181837 6 io_out[36]
port 135 nsew signal output
rlabel metal3 s 0 102688 800 102808 6 io_out[37]
port 136 nsew signal output
rlabel metal2 s 173898 181037 173954 181837 6 io_out[3]
port 137 nsew signal output
rlabel metal2 s 140778 181037 140834 181837 6 io_out[4]
port 138 nsew signal output
rlabel metal2 s 170218 181037 170274 181837 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 0 104048 800 104168 6 io_out[6]
port 140 nsew signal output
rlabel metal2 s 158718 181037 158774 181837 6 io_out[7]
port 141 nsew signal output
rlabel metal2 s 162858 0 162914 800 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 0 101328 800 101448 6 io_out[9]
port 143 nsew signal output
rlabel metal3 s 0 148248 800 148368 6 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_data_in[100]
port 145 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 la_data_in[101]
port 146 nsew signal input
rlabel metal3 s 178893 46248 179693 46368 6 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 132498 181037 132554 181837 6 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 la_data_in[104]
port 149 nsew signal input
rlabel metal3 s 0 127848 800 127968 6 la_data_in[105]
port 150 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 la_data_in[106]
port 151 nsew signal input
rlabel metal3 s 178893 138728 179693 138848 6 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_data_in[109]
port 154 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 la_data_in[10]
port 155 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 la_data_in[110]
port 156 nsew signal input
rlabel metal3 s 0 138728 800 138848 6 la_data_in[111]
port 157 nsew signal input
rlabel metal3 s 0 144168 800 144288 6 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 163778 0 163834 800 6 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 96618 181037 96674 181837 6 la_data_in[114]
port 160 nsew signal input
rlabel metal3 s 178893 42168 179693 42288 6 la_data_in[115]
port 161 nsew signal input
rlabel metal3 s 178893 113568 179693 113688 6 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 la_data_in[118]
port 164 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 la_data_in[119]
port 165 nsew signal input
rlabel metal3 s 178893 71408 179693 71528 6 la_data_in[11]
port 166 nsew signal input
rlabel metal3 s 0 56448 800 56568 6 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 142618 181037 142674 181837 6 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 54758 181037 54814 181837 6 la_data_in[124]
port 171 nsew signal input
rlabel metal3 s 178893 19728 179693 19848 6 la_data_in[125]
port 172 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 19798 181037 19854 181837 6 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 78218 181037 78274 181837 6 la_data_in[12]
port 175 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 la_data_in[13]
port 176 nsew signal input
rlabel metal3 s 178893 174768 179693 174888 6 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 la_data_in[15]
port 178 nsew signal input
rlabel metal3 s 0 146888 800 147008 6 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 938 181037 994 181837 6 la_data_in[17]
port 180 nsew signal input
rlabel metal3 s 0 145528 800 145648 6 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 13358 181037 13414 181837 6 la_data_in[19]
port 182 nsew signal input
rlabel metal3 s 178893 75488 179693 75608 6 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 130658 181037 130714 181837 6 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 109498 181037 109554 181837 6 la_data_in[21]
port 185 nsew signal input
rlabel metal3 s 178893 79568 179693 79688 6 la_data_in[22]
port 186 nsew signal input
rlabel metal3 s 178893 165248 179693 165368 6 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 120078 181037 120134 181837 6 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_data_in[27]
port 191 nsew signal input
rlabel metal3 s 178893 34008 179693 34128 6 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 95238 181037 95294 181837 6 la_data_in[2]
port 194 nsew signal input
rlabel metal3 s 178893 60528 179693 60648 6 la_data_in[30]
port 195 nsew signal input
rlabel metal3 s 178893 17008 179693 17128 6 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 34978 181037 35034 181837 6 la_data_in[32]
port 197 nsew signal input
rlabel metal3 s 178893 166608 179693 166728 6 la_data_in[33]
port 198 nsew signal input
rlabel metal3 s 178893 65968 179693 66088 6 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 144458 181037 144514 181837 6 la_data_in[35]
port 200 nsew signal input
rlabel metal3 s 178893 36728 179693 36848 6 la_data_in[36]
port 201 nsew signal input
rlabel metal3 s 0 117648 800 117768 6 la_data_in[37]
port 202 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 172978 181037 173034 181837 6 la_data_in[39]
port 204 nsew signal input
rlabel metal3 s 178893 44888 179693 45008 6 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 152278 181037 152334 181837 6 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_data_in[41]
port 207 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 56598 181037 56654 181837 6 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 127438 181037 127494 181837 6 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 89718 181037 89774 181837 6 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 42338 181037 42394 181837 6 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 30378 181037 30434 181837 6 la_data_in[47]
port 213 nsew signal input
rlabel metal3 s 178893 153688 179693 153808 6 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 6458 181037 6514 181837 6 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_data_in[4]
port 216 nsew signal input
rlabel metal3 s 178893 112208 179693 112328 6 la_data_in[50]
port 217 nsew signal input
rlabel metal3 s 0 162528 800 162648 6 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 83278 181037 83334 181837 6 la_data_in[52]
port 219 nsew signal input
rlabel metal3 s 178893 129888 179693 130008 6 la_data_in[53]
port 220 nsew signal input
rlabel metal3 s 178893 157088 179693 157208 6 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 60278 181037 60334 181837 6 la_data_in[55]
port 222 nsew signal input
rlabel metal3 s 0 120368 800 120488 6 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 64418 181037 64474 181837 6 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 169758 0 169814 800 6 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 166538 181037 166594 181837 6 la_data_in[59]
port 226 nsew signal input
rlabel metal3 s 178893 64608 179693 64728 6 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 159638 181037 159694 181837 6 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 88798 181037 88854 181837 6 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 155958 181037 156014 181837 6 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 76378 181037 76434 181837 6 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 91558 181037 91614 181837 6 la_data_in[65]
port 233 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 la_data_in[67]
port 235 nsew signal input
rlabel metal3 s 178893 51688 179693 51808 6 la_data_in[68]
port 236 nsew signal input
rlabel metal3 s 178893 177488 179693 177608 6 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 la_data_in[6]
port 238 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 la_data_in[70]
port 239 nsew signal input
rlabel metal3 s 178893 145528 179693 145648 6 la_data_in[71]
port 240 nsew signal input
rlabel metal3 s 178893 159808 179693 159928 6 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 119158 181037 119214 181837 6 la_data_in[73]
port 242 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 la_data_in[74]
port 243 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 39578 181037 39634 181837 6 la_data_in[78]
port 247 nsew signal input
rlabel metal3 s 178893 92488 179693 92608 6 la_data_in[79]
port 248 nsew signal input
rlabel metal3 s 0 93848 800 93968 6 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 20718 181037 20774 181837 6 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 154118 181037 154174 181837 6 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 177578 181037 177634 181837 6 la_data_in[84]
port 254 nsew signal input
rlabel metal3 s 0 159808 800 159928 6 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 100298 181037 100354 181837 6 la_data_in[86]
port 256 nsew signal input
rlabel metal3 s 0 116288 800 116408 6 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 29458 181037 29514 181837 6 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 97538 181037 97594 181837 6 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 la_data_in[8]
port 260 nsew signal input
rlabel metal3 s 178893 116288 179693 116408 6 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 135258 181037 135314 181837 6 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 65338 181037 65394 181837 6 la_data_in[93]
port 264 nsew signal input
rlabel metal3 s 0 167968 800 168088 6 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 146758 0 146814 800 6 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 177118 0 177174 800 6 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 129738 181037 129794 181837 6 la_data_in[98]
port 269 nsew signal input
rlabel metal3 s 178893 99288 179693 99408 6 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 151358 181037 151414 181837 6 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 88338 0 88394 800 6 la_data_out[100]
port 273 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 la_data_out[101]
port 274 nsew signal output
rlabel metal3 s 178893 123088 179693 123208 6 la_data_out[102]
port 275 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 102138 181037 102194 181837 6 la_data_out[104]
port 277 nsew signal output
rlabel metal3 s 0 165248 800 165368 6 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 125138 0 125194 800 6 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 72238 0 72294 800 6 la_data_out[107]
port 280 nsew signal output
rlabel metal3 s 178893 1368 179693 1488 6 la_data_out[108]
port 281 nsew signal output
rlabel metal3 s 0 150288 800 150408 6 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 53838 181037 53894 181837 6 la_data_out[10]
port 283 nsew signal output
rlabel metal3 s 0 95208 800 95328 6 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 34058 181037 34114 181837 6 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 103518 0 103574 800 6 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 143538 181037 143594 181837 6 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 113638 181037 113694 181837 6 la_data_out[114]
port 288 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 la_data_out[115]
port 289 nsew signal output
rlabel metal3 s 0 99968 800 100088 6 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 48318 181037 48374 181837 6 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 43258 181037 43314 181837 6 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 178498 181037 178554 181837 6 la_data_out[119]
port 293 nsew signal output
rlabel metal3 s 178893 136008 179693 136128 6 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 la_data_out[120]
port 295 nsew signal output
rlabel metal3 s 0 172048 800 172168 6 la_data_out[121]
port 296 nsew signal output
rlabel metal3 s 0 67328 800 67448 6 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 175738 181037 175794 181837 6 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 172518 0 172574 800 6 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 la_data_out[125]
port 300 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 la_data_out[126]
port 301 nsew signal output
rlabel metal3 s 0 166608 800 166728 6 la_data_out[127]
port 302 nsew signal output
rlabel metal3 s 178893 102008 179693 102128 6 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 159178 0 159234 800 6 la_data_out[13]
port 304 nsew signal output
rlabel metal3 s 178893 78208 179693 78328 6 la_data_out[14]
port 305 nsew signal output
rlabel metal3 s 0 126488 800 126608 6 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 174358 0 174414 800 6 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 61198 181037 61254 181837 6 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 124218 0 124274 800 6 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 133418 181037 133474 181837 6 la_data_out[21]
port 313 nsew signal output
rlabel metal3 s 178893 131248 179693 131368 6 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 71778 181037 71834 181837 6 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 66258 181037 66314 181837 6 la_data_out[24]
port 316 nsew signal output
rlabel metal3 s 178893 162528 179693 162648 6 la_data_out[25]
port 317 nsew signal output
rlabel metal3 s 178893 11568 179693 11688 6 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 128818 0 128874 800 6 la_data_out[27]
port 319 nsew signal output
rlabel metal3 s 178893 48968 179693 49088 6 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 la_data_out[2]
port 322 nsew signal output
rlabel metal3 s 178893 82968 179693 83088 6 la_data_out[30]
port 323 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 la_data_out[31]
port 324 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 35898 181037 35954 181837 6 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 la_data_out[34]
port 327 nsew signal output
rlabel metal3 s 178893 87048 179693 87168 6 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 173438 0 173494 800 6 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 150438 0 150494 800 6 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 172058 181037 172114 181837 6 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 la_data_out[39]
port 332 nsew signal output
rlabel metal3 s 0 153008 800 153128 6 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 118698 0 118754 800 6 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 la_data_out[41]
port 335 nsew signal output
rlabel metal3 s 178893 96568 179693 96688 6 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 164698 0 164754 800 6 la_data_out[45]
port 339 nsew signal output
rlabel metal3 s 178893 39448 179693 39568 6 la_data_out[46]
port 340 nsew signal output
rlabel metal3 s 178893 23808 179693 23928 6 la_data_out[47]
port 341 nsew signal output
rlabel metal3 s 178893 8848 179693 8968 6 la_data_out[48]
port 342 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 la_data_out[49]
port 343 nsew signal output
rlabel metal3 s 178893 104728 179693 104848 6 la_data_out[4]
port 344 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 126518 181037 126574 181837 6 la_data_out[51]
port 346 nsew signal output
rlabel metal3 s 178893 91128 179693 91248 6 la_data_out[52]
port 347 nsew signal output
rlabel metal3 s 178893 176128 179693 176248 6 la_data_out[53]
port 348 nsew signal output
rlabel metal3 s 178893 180208 179693 180328 6 la_data_out[54]
port 349 nsew signal output
rlabel metal3 s 0 65968 800 66088 6 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 151818 0 151874 800 6 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 78678 0 78734 800 6 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 77298 181037 77354 181837 6 la_data_out[58]
port 353 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 155038 181037 155094 181837 6 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 155498 0 155554 800 6 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 la_data_out[61]
port 357 nsew signal output
rlabel metal3 s 0 72768 800 72888 6 la_data_out[62]
port 358 nsew signal output
rlabel metal3 s 178893 50328 179693 50448 6 la_data_out[63]
port 359 nsew signal output
rlabel metal3 s 178893 63248 179693 63368 6 la_data_out[64]
port 360 nsew signal output
rlabel metal3 s 178893 27888 179693 28008 6 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 99378 181037 99434 181837 6 la_data_out[66]
port 362 nsew signal output
rlabel metal3 s 178893 35368 179693 35488 6 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 98458 181037 98514 181837 6 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 la_data_out[69]
port 365 nsew signal output
rlabel metal3 s 0 154368 800 154488 6 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 51998 181037 52054 181837 6 la_data_out[70]
port 367 nsew signal output
rlabel metal3 s 178893 163888 179693 164008 6 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 171138 181037 171194 181837 6 la_data_out[72]
port 369 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 la_data_out[73]
port 370 nsew signal output
rlabel metal3 s 0 121728 800 121848 6 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 91098 0 91154 800 6 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 la_data_out[77]
port 374 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 103978 181037 104034 181837 6 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 174818 181037 174874 181837 6 la_data_out[7]
port 377 nsew signal output
rlabel metal3 s 178893 120368 179693 120488 6 la_data_out[80]
port 378 nsew signal output
rlabel metal3 s 178893 31968 179693 32088 6 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 86038 181037 86094 181837 6 la_data_out[82]
port 380 nsew signal output
rlabel metal3 s 0 55088 800 55208 6 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 92938 0 92994 800 6 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 147678 0 147734 800 6 la_data_out[85]
port 383 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 la_data_out[86]
port 384 nsew signal output
rlabel metal3 s 178893 70048 179693 70168 6 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 162858 181037 162914 181837 6 la_data_out[88]
port 386 nsew signal output
rlabel metal3 s 0 123088 800 123208 6 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 124678 181037 124734 181837 6 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 28078 181037 28134 181837 6 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 25318 181037 25374 181837 6 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 123758 181037 123814 181837 6 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 138938 181037 138994 181837 6 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 2318 0 2374 800 6 la_data_out[94]
port 393 nsew signal output
rlabel metal3 s 178893 61888 179693 62008 6 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 57518 181037 57574 181837 6 la_data_out[96]
port 395 nsew signal output
rlabel metal3 s 0 97928 800 98048 6 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 102598 0 102654 800 6 la_data_out[98]
port 397 nsew signal output
rlabel metal3 s 178893 133288 179693 133408 6 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 95698 0 95754 800 6 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 la_oenb[100]
port 401 nsew signal input
rlabel metal3 s 178893 6808 179693 6928 6 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 44178 181037 44234 181837 6 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 la_oenb[104]
port 405 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 la_oenb[105]
port 406 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 la_oenb[106]
port 407 nsew signal input
rlabel metal3 s 0 92488 800 92608 6 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 105818 181037 105874 181837 6 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 51078 181037 51134 181837 6 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 69018 181037 69074 181837 6 la_oenb[110]
port 412 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 la_oenb[111]
port 413 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 143998 0 144054 800 6 la_oenb[113]
port 415 nsew signal input
rlabel metal3 s 178893 170688 179693 170808 6 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 la_oenb[115]
port 417 nsew signal input
rlabel metal3 s 0 57808 800 57928 6 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 55678 181037 55734 181837 6 la_oenb[117]
port 419 nsew signal input
rlabel metal3 s 178893 148248 179693 148368 6 la_oenb[118]
port 420 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 161478 181037 161534 181837 6 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 la_oenb[120]
port 423 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 la_oenb[121]
port 424 nsew signal input
rlabel metal3 s 178893 125808 179693 125928 6 la_oenb[122]
port 425 nsew signal input
rlabel metal3 s 178893 18368 179693 18488 6 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 171598 0 171654 800 6 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 7378 181037 7434 181837 6 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 la_oenb[127]
port 430 nsew signal input
rlabel metal3 s 178893 146888 179693 147008 6 la_oenb[12]
port 431 nsew signal input
rlabel metal3 s 178893 121728 179693 121848 6 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 146758 181037 146814 181837 6 la_oenb[14]
port 433 nsew signal input
rlabel metal3 s 178893 124448 179693 124568 6 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 21638 181037 21694 181837 6 la_oenb[17]
port 436 nsew signal input
rlabel metal3 s 178893 114928 179693 115048 6 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 157338 0 157394 800 6 la_oenb[19]
port 438 nsew signal input
rlabel metal3 s 0 179528 800 179648 6 la_oenb[1]
port 439 nsew signal input
rlabel metal3 s 178893 95208 179693 95328 6 la_oenb[20]
port 440 nsew signal input
rlabel metal3 s 0 155728 800 155848 6 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 93398 181037 93454 181837 6 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 67178 181037 67234 181837 6 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 139858 181037 139914 181837 6 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 16118 181037 16174 181837 6 la_oenb[27]
port 447 nsew signal input
rlabel metal3 s 178893 14288 179693 14408 6 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 la_oenb[29]
port 449 nsew signal input
rlabel metal3 s 178893 97928 179693 98048 6 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 la_oenb[31]
port 452 nsew signal input
rlabel metal3 s 178893 72768 179693 72888 6 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 92478 181037 92534 181837 6 la_oenb[33]
port 454 nsew signal input
rlabel metal3 s 178893 57128 179693 57248 6 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 178038 0 178094 800 6 la_oenb[37]
port 458 nsew signal input
rlabel metal3 s 178893 158448 179693 158568 6 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_oenb[39]
port 460 nsew signal input
rlabel metal3 s 0 141448 800 141568 6 la_oenb[3]
port 461 nsew signal input
rlabel metal3 s 0 125128 800 125248 6 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 111338 181037 111394 181837 6 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_oenb[42]
port 464 nsew signal input
rlabel metal3 s 178893 76848 179693 76968 6 la_oenb[43]
port 465 nsew signal input
rlabel metal3 s 0 161168 800 161288 6 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 la_oenb[45]
port 467 nsew signal input
rlabel metal3 s 178893 68688 179693 68808 6 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 169298 181037 169354 181837 6 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 72698 181037 72754 181837 6 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 478 0 534 800 6 la_oenb[4]
port 472 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 1858 181037 1914 181837 6 la_oenb[51]
port 474 nsew signal input
rlabel metal3 s 178893 38088 179693 38208 6 la_oenb[52]
port 475 nsew signal input
rlabel metal3 s 178893 88408 179693 88528 6 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_oenb[54]
port 477 nsew signal input
rlabel metal3 s 0 136008 800 136128 6 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 41418 181037 41474 181837 6 la_oenb[56]
port 479 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 152738 0 152794 800 6 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 94318 181037 94374 181837 6 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 121918 181037 121974 181837 6 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 123298 0 123354 800 6 la_oenb[60]
port 484 nsew signal input
rlabel metal3 s 178893 55768 179693 55888 6 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 la_oenb[62]
port 486 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 la_oenb[63]
port 487 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 la_oenb[64]
port 488 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 11058 181037 11114 181837 6 la_oenb[66]
port 490 nsew signal input
rlabel metal3 s 178893 22448 179693 22568 6 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 103058 181037 103114 181837 6 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 140318 0 140374 800 6 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 128358 181037 128414 181837 6 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 50158 181037 50214 181837 6 la_oenb[71]
port 496 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 134798 0 134854 800 6 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 80518 181037 80574 181837 6 la_oenb[74]
port 499 nsew signal input
rlabel metal3 s 0 169328 800 169448 6 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 18878 181037 18934 181837 6 la_oenb[76]
port 501 nsew signal input
rlabel metal3 s 178893 5448 179693 5568 6 la_oenb[77]
port 502 nsew signal input
rlabel metal3 s 0 178168 800 178288 6 la_oenb[78]
port 503 nsew signal input
rlabel metal3 s 178893 43528 179693 43648 6 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_oenb[7]
port 505 nsew signal input
rlabel metal3 s 178893 150968 179693 151088 6 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 136178 181037 136234 181837 6 la_oenb[81]
port 507 nsew signal input
rlabel metal3 s 0 119008 800 119128 6 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 135718 0 135774 800 6 la_oenb[83]
port 509 nsew signal input
rlabel metal3 s 0 105408 800 105528 6 la_oenb[84]
port 510 nsew signal input
rlabel metal3 s 178893 84328 179693 84448 6 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 153198 181037 153254 181837 6 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 75458 181037 75514 181837 6 la_oenb[87]
port 513 nsew signal input
rlabel metal3 s 178893 172048 179693 172168 6 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_oenb[89]
port 515 nsew signal input
rlabel metal3 s 178893 137368 179693 137488 6 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 115478 181037 115534 181837 6 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 176658 181037 176714 181837 6 la_oenb[93]
port 520 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 la_oenb[94]
port 521 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 la_oenb[96]
port 523 nsew signal input
rlabel metal3 s 178893 149608 179693 149728 6 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 90638 181037 90694 181837 6 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 150438 181037 150494 181837 6 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 user_clock2
port 528 nsew signal input
rlabel metal2 s 26238 181037 26294 181837 6 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 131578 181037 131634 181837 6 user_irq[2]
port 531 nsew signal output
rlabel metal2 s 86958 181037 87014 181837 6 wb_clk_i
port 532 nsew signal input
rlabel metal3 s 178893 4088 179693 4208 6 wb_rst_i
port 533 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 wbs_ack_o
port 534 nsew signal output
rlabel metal2 s 85118 181037 85174 181837 6 wbs_adr_i[0]
port 535 nsew signal input
rlabel metal3 s 178893 53048 179693 53168 6 wbs_adr_i[10]
port 536 nsew signal input
rlabel metal2 s 176198 0 176254 800 6 wbs_adr_i[11]
port 537 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 wbs_adr_i[12]
port 538 nsew signal input
rlabel metal3 s 0 176808 800 176928 6 wbs_adr_i[13]
port 539 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 wbs_adr_i[14]
port 540 nsew signal input
rlabel metal3 s 0 106768 800 106888 6 wbs_adr_i[15]
port 541 nsew signal input
rlabel metal3 s 178893 141448 179693 141568 6 wbs_adr_i[16]
port 542 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 wbs_adr_i[17]
port 543 nsew signal input
rlabel metal3 s 178893 12928 179693 13048 6 wbs_adr_i[18]
port 544 nsew signal input
rlabel metal2 s 107658 181037 107714 181837 6 wbs_adr_i[19]
port 545 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_adr_i[1]
port 546 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 wbs_adr_i[20]
port 547 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_adr_i[21]
port 548 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 wbs_adr_i[22]
port 549 nsew signal input
rlabel metal2 s 73618 181037 73674 181837 6 wbs_adr_i[23]
port 550 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_adr_i[24]
port 551 nsew signal input
rlabel metal2 s 166538 0 166594 800 6 wbs_adr_i[25]
port 552 nsew signal input
rlabel metal3 s 0 140088 800 140208 6 wbs_adr_i[26]
port 553 nsew signal input
rlabel metal2 s 116398 181037 116454 181837 6 wbs_adr_i[27]
port 554 nsew signal input
rlabel metal2 s 9218 181037 9274 181837 6 wbs_adr_i[28]
port 555 nsew signal input
rlabel metal3 s 178893 178848 179693 178968 6 wbs_adr_i[29]
port 556 nsew signal input
rlabel metal2 s 22558 181037 22614 181837 6 wbs_adr_i[2]
port 557 nsew signal input
rlabel metal2 s 70858 181037 70914 181837 6 wbs_adr_i[30]
port 558 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_adr_i[31]
port 559 nsew signal input
rlabel metal3 s 178893 100648 179693 100768 6 wbs_adr_i[3]
port 560 nsew signal input
rlabel metal2 s 37738 181037 37794 181837 6 wbs_adr_i[4]
port 561 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 wbs_adr_i[5]
port 562 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 wbs_adr_i[6]
port 563 nsew signal input
rlabel metal2 s 158258 0 158314 800 6 wbs_adr_i[7]
port 564 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 wbs_adr_i[8]
port 565 nsew signal input
rlabel metal3 s 0 109488 800 109608 6 wbs_adr_i[9]
port 566 nsew signal input
rlabel metal2 s 87878 181037 87934 181837 6 wbs_cyc_i
port 567 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 wbs_dat_i[0]
port 568 nsew signal input
rlabel metal2 s 130658 0 130714 800 6 wbs_dat_i[10]
port 569 nsew signal input
rlabel metal3 s 0 129208 800 129328 6 wbs_dat_i[11]
port 570 nsew signal input
rlabel metal2 s 147678 181037 147734 181837 6 wbs_dat_i[12]
port 571 nsew signal input
rlabel metal3 s 178893 152328 179693 152448 6 wbs_dat_i[13]
port 572 nsew signal input
rlabel metal3 s 178893 54408 179693 54528 6 wbs_dat_i[14]
port 573 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 wbs_dat_i[15]
port 574 nsew signal input
rlabel metal3 s 0 70048 800 70168 6 wbs_dat_i[16]
port 575 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 wbs_dat_i[17]
port 576 nsew signal input
rlabel metal3 s 0 134648 800 134768 6 wbs_dat_i[18]
port 577 nsew signal input
rlabel metal2 s 122838 181037 122894 181837 6 wbs_dat_i[19]
port 578 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 wbs_dat_i[1]
port 579 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 wbs_dat_i[20]
port 580 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_dat_i[21]
port 581 nsew signal input
rlabel metal2 s 165618 181037 165674 181837 6 wbs_dat_i[22]
port 582 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 wbs_dat_i[23]
port 583 nsew signal input
rlabel metal2 s 17958 181037 18014 181837 6 wbs_dat_i[24]
port 584 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 wbs_dat_i[25]
port 585 nsew signal input
rlabel metal3 s 178893 21088 179693 21208 6 wbs_dat_i[26]
port 586 nsew signal input
rlabel metal3 s 178893 59168 179693 59288 6 wbs_dat_i[27]
port 587 nsew signal input
rlabel metal2 s 58438 181037 58494 181837 6 wbs_dat_i[28]
port 588 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 wbs_dat_i[29]
port 589 nsew signal input
rlabel metal3 s 178893 169328 179693 169448 6 wbs_dat_i[2]
port 590 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 wbs_dat_i[30]
port 591 nsew signal input
rlabel metal2 s 45558 181037 45614 181837 6 wbs_dat_i[31]
port 592 nsew signal input
rlabel metal2 s 117318 181037 117374 181837 6 wbs_dat_i[3]
port 593 nsew signal input
rlabel metal3 s 0 158448 800 158568 6 wbs_dat_i[4]
port 594 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_i[5]
port 595 nsew signal input
rlabel metal2 s 141698 181037 141754 181837 6 wbs_dat_i[6]
port 596 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_i[7]
port 597 nsew signal input
rlabel metal2 s 112718 181037 112774 181837 6 wbs_dat_i[8]
port 598 nsew signal input
rlabel metal3 s 0 163888 800 164008 6 wbs_dat_i[9]
port 599 nsew signal input
rlabel metal2 s 5538 181037 5594 181837 6 wbs_dat_o[0]
port 600 nsew signal output
rlabel metal3 s 178893 144168 179693 144288 6 wbs_dat_o[10]
port 601 nsew signal output
rlabel metal2 s 115478 0 115534 800 6 wbs_dat_o[11]
port 602 nsew signal output
rlabel metal2 s 167918 0 167974 800 6 wbs_dat_o[12]
port 603 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_o[13]
port 604 nsew signal output
rlabel metal3 s 0 133288 800 133408 6 wbs_dat_o[14]
port 605 nsew signal output
rlabel metal2 s 170678 0 170734 800 6 wbs_dat_o[15]
port 606 nsew signal output
rlabel metal2 s 138018 181037 138074 181837 6 wbs_dat_o[16]
port 607 nsew signal output
rlabel metal2 s 2778 181037 2834 181837 6 wbs_dat_o[17]
port 608 nsew signal output
rlabel metal3 s 178893 89768 179693 89888 6 wbs_dat_o[18]
port 609 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 wbs_dat_o[19]
port 610 nsew signal output
rlabel metal2 s 93858 0 93914 800 6 wbs_dat_o[1]
port 611 nsew signal output
rlabel metal2 s 74538 181037 74594 181837 6 wbs_dat_o[20]
port 612 nsew signal output
rlabel metal2 s 40498 181037 40554 181837 6 wbs_dat_o[21]
port 613 nsew signal output
rlabel metal2 s 132498 0 132554 800 6 wbs_dat_o[22]
port 614 nsew signal output
rlabel metal2 s 8298 181037 8354 181837 6 wbs_dat_o[23]
port 615 nsew signal output
rlabel metal2 s 114558 181037 114614 181837 6 wbs_dat_o[24]
port 616 nsew signal output
rlabel metal3 s 178893 119008 179693 119128 6 wbs_dat_o[25]
port 617 nsew signal output
rlabel metal2 s 125598 181037 125654 181837 6 wbs_dat_o[26]
port 618 nsew signal output
rlabel metal2 s 148598 181037 148654 181837 6 wbs_dat_o[27]
port 619 nsew signal output
rlabel metal3 s 178893 47608 179693 47728 6 wbs_dat_o[28]
port 620 nsew signal output
rlabel metal2 s 27158 181037 27214 181837 6 wbs_dat_o[29]
port 621 nsew signal output
rlabel metal3 s 0 110848 800 110968 6 wbs_dat_o[2]
port 622 nsew signal output
rlabel metal2 s 137098 181037 137154 181837 6 wbs_dat_o[30]
port 623 nsew signal output
rlabel metal2 s 49238 181037 49294 181837 6 wbs_dat_o[31]
port 624 nsew signal output
rlabel metal3 s 0 112208 800 112328 6 wbs_dat_o[3]
port 625 nsew signal output
rlabel metal2 s 31298 181037 31354 181837 6 wbs_dat_o[4]
port 626 nsew signal output
rlabel metal2 s 106738 181037 106794 181837 6 wbs_dat_o[5]
port 627 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 wbs_dat_o[6]
port 628 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_o[7]
port 629 nsew signal output
rlabel metal3 s 178893 127168 179693 127288 6 wbs_dat_o[8]
port 630 nsew signal output
rlabel metal3 s 178893 128528 179693 128648 6 wbs_dat_o[9]
port 631 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 wbs_sel_i[0]
port 632 nsew signal input
rlabel metal2 s 17038 181037 17094 181837 6 wbs_sel_i[1]
port 633 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 wbs_sel_i[2]
port 634 nsew signal input
rlabel metal2 s 33138 181037 33194 181837 6 wbs_sel_i[3]
port 635 nsew signal input
rlabel metal2 s 120538 0 120594 800 6 wbs_stb_i
port 636 nsew signal input
rlabel metal2 s 101218 181037 101274 181837 6 wbs_we_i
port 637 nsew signal input
rlabel metal4 s 144804 -1864 145404 183560 6 vccd1
port 638 nsew power bidirectional
rlabel metal4 s 108804 -1864 109404 183560 6 vccd1
port 639 nsew power bidirectional
rlabel metal4 s 72804 -1864 73404 183560 6 vccd1
port 640 nsew power bidirectional
rlabel metal4 s 36804 -1864 37404 183560 6 vccd1
port 641 nsew power bidirectional
rlabel metal4 s 804 -1864 1404 183560 6 vccd1
port 642 nsew power bidirectional
rlabel metal4 s 181072 -924 181672 182620 6 vccd1
port 643 nsew power bidirectional
rlabel metal4 s -1996 -924 -1396 182620 4 vccd1
port 644 nsew power bidirectional
rlabel metal5 s -1996 182020 181672 182620 6 vccd1
port 645 nsew power bidirectional
rlabel metal5 s -2936 145828 182612 146428 6 vccd1
port 646 nsew power bidirectional
rlabel metal5 s -2936 109828 182612 110428 6 vccd1
port 647 nsew power bidirectional
rlabel metal5 s -2936 73828 182612 74428 6 vccd1
port 648 nsew power bidirectional
rlabel metal5 s -2936 37828 182612 38428 6 vccd1
port 649 nsew power bidirectional
rlabel metal5 s -2936 1828 182612 2428 6 vccd1
port 650 nsew power bidirectional
rlabel metal5 s -1996 -924 181672 -324 8 vccd1
port 651 nsew power bidirectional
rlabel metal4 s 182012 -1864 182612 183560 6 vssd1
port 652 nsew ground bidirectional
rlabel metal4 s 162804 -1864 163404 183560 6 vssd1
port 653 nsew ground bidirectional
rlabel metal4 s 126804 -1864 127404 183560 6 vssd1
port 654 nsew ground bidirectional
rlabel metal4 s 90804 -1864 91404 183560 6 vssd1
port 655 nsew ground bidirectional
rlabel metal4 s 54804 -1864 55404 183560 6 vssd1
port 656 nsew ground bidirectional
rlabel metal4 s 18804 -1864 19404 183560 6 vssd1
port 657 nsew ground bidirectional
rlabel metal4 s -2936 -1864 -2336 183560 4 vssd1
port 658 nsew ground bidirectional
rlabel metal5 s -2936 182960 182612 183560 6 vssd1
port 659 nsew ground bidirectional
rlabel metal5 s -2936 163828 182612 164428 6 vssd1
port 660 nsew ground bidirectional
rlabel metal5 s -2936 127828 182612 128428 6 vssd1
port 661 nsew ground bidirectional
rlabel metal5 s -2936 91828 182612 92428 6 vssd1
port 662 nsew ground bidirectional
rlabel metal5 s -2936 55828 182612 56428 6 vssd1
port 663 nsew ground bidirectional
rlabel metal5 s -2936 19828 182612 20428 6 vssd1
port 664 nsew ground bidirectional
rlabel metal5 s -2936 -1864 182612 -1264 8 vssd1
port 665 nsew ground bidirectional
rlabel metal4 s 148404 -3744 149004 185440 6 vccd2
port 666 nsew power bidirectional
rlabel metal4 s 112404 -3744 113004 185440 6 vccd2
port 667 nsew power bidirectional
rlabel metal4 s 76404 -3744 77004 185440 6 vccd2
port 668 nsew power bidirectional
rlabel metal4 s 40404 -3744 41004 185440 6 vccd2
port 669 nsew power bidirectional
rlabel metal4 s 4404 -3744 5004 185440 6 vccd2
port 670 nsew power bidirectional
rlabel metal4 s 182952 -2804 183552 184500 6 vccd2
port 671 nsew power bidirectional
rlabel metal4 s -3876 -2804 -3276 184500 4 vccd2
port 672 nsew power bidirectional
rlabel metal5 s -3876 183900 183552 184500 6 vccd2
port 673 nsew power bidirectional
rlabel metal5 s -4816 149476 184492 150076 6 vccd2
port 674 nsew power bidirectional
rlabel metal5 s -4816 113476 184492 114076 6 vccd2
port 675 nsew power bidirectional
rlabel metal5 s -4816 77476 184492 78076 6 vccd2
port 676 nsew power bidirectional
rlabel metal5 s -4816 41476 184492 42076 6 vccd2
port 677 nsew power bidirectional
rlabel metal5 s -4816 5476 184492 6076 6 vccd2
port 678 nsew power bidirectional
rlabel metal5 s -3876 -2804 183552 -2204 8 vccd2
port 679 nsew power bidirectional
rlabel metal4 s 183892 -3744 184492 185440 6 vssd2
port 680 nsew ground bidirectional
rlabel metal4 s 166404 -3744 167004 185440 6 vssd2
port 681 nsew ground bidirectional
rlabel metal4 s 130404 -3744 131004 185440 6 vssd2
port 682 nsew ground bidirectional
rlabel metal4 s 94404 -3744 95004 185440 6 vssd2
port 683 nsew ground bidirectional
rlabel metal4 s 58404 -3744 59004 185440 6 vssd2
port 684 nsew ground bidirectional
rlabel metal4 s 22404 -3744 23004 185440 6 vssd2
port 685 nsew ground bidirectional
rlabel metal4 s -4816 -3744 -4216 185440 4 vssd2
port 686 nsew ground bidirectional
rlabel metal5 s -4816 184840 184492 185440 6 vssd2
port 687 nsew ground bidirectional
rlabel metal5 s -4816 167476 184492 168076 6 vssd2
port 688 nsew ground bidirectional
rlabel metal5 s -4816 131476 184492 132076 6 vssd2
port 689 nsew ground bidirectional
rlabel metal5 s -4816 95476 184492 96076 6 vssd2
port 690 nsew ground bidirectional
rlabel metal5 s -4816 59476 184492 60076 6 vssd2
port 691 nsew ground bidirectional
rlabel metal5 s -4816 23476 184492 24076 6 vssd2
port 692 nsew ground bidirectional
rlabel metal5 s -4816 -3744 184492 -3144 8 vssd2
port 693 nsew ground bidirectional
rlabel metal4 s 152004 -5624 152604 187320 6 vdda1
port 694 nsew power bidirectional
rlabel metal4 s 116004 -5624 116604 187320 6 vdda1
port 695 nsew power bidirectional
rlabel metal4 s 80004 -5624 80604 187320 6 vdda1
port 696 nsew power bidirectional
rlabel metal4 s 44004 -5624 44604 187320 6 vdda1
port 697 nsew power bidirectional
rlabel metal4 s 8004 -5624 8604 187320 6 vdda1
port 698 nsew power bidirectional
rlabel metal4 s 184832 -4684 185432 186380 6 vdda1
port 699 nsew power bidirectional
rlabel metal4 s -5756 -4684 -5156 186380 4 vdda1
port 700 nsew power bidirectional
rlabel metal5 s -5756 185780 185432 186380 6 vdda1
port 701 nsew power bidirectional
rlabel metal5 s -6696 153076 186372 153676 6 vdda1
port 702 nsew power bidirectional
rlabel metal5 s -6696 117076 186372 117676 6 vdda1
port 703 nsew power bidirectional
rlabel metal5 s -6696 81076 186372 81676 6 vdda1
port 704 nsew power bidirectional
rlabel metal5 s -6696 45076 186372 45676 6 vdda1
port 705 nsew power bidirectional
rlabel metal5 s -6696 9076 186372 9676 6 vdda1
port 706 nsew power bidirectional
rlabel metal5 s -5756 -4684 185432 -4084 8 vdda1
port 707 nsew power bidirectional
rlabel metal4 s 185772 -5624 186372 187320 6 vssa1
port 708 nsew ground bidirectional
rlabel metal4 s 170004 -5624 170604 187320 6 vssa1
port 709 nsew ground bidirectional
rlabel metal4 s 134004 -5624 134604 187320 6 vssa1
port 710 nsew ground bidirectional
rlabel metal4 s 98004 -5624 98604 187320 6 vssa1
port 711 nsew ground bidirectional
rlabel metal4 s 62004 -5624 62604 187320 6 vssa1
port 712 nsew ground bidirectional
rlabel metal4 s 26004 -5624 26604 187320 6 vssa1
port 713 nsew ground bidirectional
rlabel metal4 s -6696 -5624 -6096 187320 4 vssa1
port 714 nsew ground bidirectional
rlabel metal5 s -6696 186720 186372 187320 6 vssa1
port 715 nsew ground bidirectional
rlabel metal5 s -6696 171076 186372 171676 6 vssa1
port 716 nsew ground bidirectional
rlabel metal5 s -6696 135076 186372 135676 6 vssa1
port 717 nsew ground bidirectional
rlabel metal5 s -6696 99076 186372 99676 6 vssa1
port 718 nsew ground bidirectional
rlabel metal5 s -6696 63076 186372 63676 6 vssa1
port 719 nsew ground bidirectional
rlabel metal5 s -6696 27076 186372 27676 6 vssa1
port 720 nsew ground bidirectional
rlabel metal5 s -6696 -5624 186372 -5024 8 vssa1
port 721 nsew ground bidirectional
rlabel metal4 s 155604 -7504 156204 189200 6 vdda2
port 722 nsew power bidirectional
rlabel metal4 s 119604 -7504 120204 189200 6 vdda2
port 723 nsew power bidirectional
rlabel metal4 s 83604 -7504 84204 189200 6 vdda2
port 724 nsew power bidirectional
rlabel metal4 s 47604 -7504 48204 189200 6 vdda2
port 725 nsew power bidirectional
rlabel metal4 s 11604 -7504 12204 189200 6 vdda2
port 726 nsew power bidirectional
rlabel metal4 s 186712 -6564 187312 188260 6 vdda2
port 727 nsew power bidirectional
rlabel metal4 s -7636 -6564 -7036 188260 4 vdda2
port 728 nsew power bidirectional
rlabel metal5 s -7636 187660 187312 188260 6 vdda2
port 729 nsew power bidirectional
rlabel metal5 s -8576 156676 188252 157276 6 vdda2
port 730 nsew power bidirectional
rlabel metal5 s -8576 120676 188252 121276 6 vdda2
port 731 nsew power bidirectional
rlabel metal5 s -8576 84676 188252 85276 6 vdda2
port 732 nsew power bidirectional
rlabel metal5 s -8576 48676 188252 49276 6 vdda2
port 733 nsew power bidirectional
rlabel metal5 s -8576 12676 188252 13276 6 vdda2
port 734 nsew power bidirectional
rlabel metal5 s -7636 -6564 187312 -5964 8 vdda2
port 735 nsew power bidirectional
rlabel metal4 s 187652 -7504 188252 189200 6 vssa2
port 736 nsew ground bidirectional
rlabel metal4 s 173604 -7504 174204 189200 6 vssa2
port 737 nsew ground bidirectional
rlabel metal4 s 137604 -7504 138204 189200 6 vssa2
port 738 nsew ground bidirectional
rlabel metal4 s 101604 -7504 102204 189200 6 vssa2
port 739 nsew ground bidirectional
rlabel metal4 s 65604 -7504 66204 189200 6 vssa2
port 740 nsew ground bidirectional
rlabel metal4 s 29604 -7504 30204 189200 6 vssa2
port 741 nsew ground bidirectional
rlabel metal4 s -8576 -7504 -7976 189200 4 vssa2
port 742 nsew ground bidirectional
rlabel metal5 s -8576 188600 188252 189200 6 vssa2
port 743 nsew ground bidirectional
rlabel metal5 s -8576 174676 188252 175276 6 vssa2
port 744 nsew ground bidirectional
rlabel metal5 s -8576 138676 188252 139276 6 vssa2
port 745 nsew ground bidirectional
rlabel metal5 s -8576 102676 188252 103276 6 vssa2
port 746 nsew ground bidirectional
rlabel metal5 s -8576 66676 188252 67276 6 vssa2
port 747 nsew ground bidirectional
rlabel metal5 s -8576 30676 188252 31276 6 vssa2
port 748 nsew ground bidirectional
rlabel metal5 s -8576 -7504 188252 -6904 8 vssa2
port 749 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 179693 181837
string LEFview TRUE
string GDS_FILE /project/openlane/user_project_wrapper/runs/user_project_wrapper/results/magic/user_project_wrapper.gds
string GDS_END 72477894
string GDS_START 130
<< end >>

