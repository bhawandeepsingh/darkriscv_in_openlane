module user_project_wrapper (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    vccd1,
    vssd1,
    vccd2,
    vssd2,
    vdda1,
    vssa1,
    vdda2,
    vssa2,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input vccd1;
 input vssd1;
 input vccd2;
 input vssd2;
 input vdda1;
 input vssa1;
 input vdda2;
 input vssa2;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 sky130_fd_sc_hd__inv_2 _11370_ (.A(\design_top.DATAO[14] ),
    .Y(_10587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11371_ (.A(_10587_),
    .X(_10588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11372_ (.A(_10588_),
    .X(_10589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11373_ (.A(\design_top.DACK[0] ),
    .Y(_01982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11374_ (.A(\design_top.core0.FLUSH[1] ),
    .Y(_10590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11375_ (.A(\design_top.core0.FLUSH[0] ),
    .Y(_10591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _11376_ (.A(_10590_),
    .B(_10591_),
    .C(\design_top.core0.XLCC ),
    .X(_10592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11377_ (.A(_10592_),
    .X(io_out[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11378_ (.A1(_01982_),
    .A2(\design_top.DACK[1] ),
    .B1(io_out[12]),
    .Y(_10593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11379_ (.A(_10593_),
    .Y(_10594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11380_ (.A(\design_top.core0.FLUSH[1] ),
    .B(\design_top.core0.FLUSH[0] ),
    .X(_10595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11381_ (.A(_10595_),
    .Y(_02661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _11382_ (.A(\design_top.core0.XSCC ),
    .B(_02661_),
    .Y(_10596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11383_ (.A(\design_top.core0.SIMM[30] ),
    .Y(_02690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11384_ (.A(_02689_),
    .X(_10597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11385_ (.A(_10597_),
    .Y(_10598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11386_ (.A1(\design_top.core0.SIMM[30] ),
    .A2(_10597_),
    .B1(_02690_),
    .B2(_10598_),
    .X(_10599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11387_ (.A(\design_top.core0.SIMM[29] ),
    .X(_10600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11388_ (.A(\design_top.core0.SIMM[29] ),
    .B(_02695_),
    .Y(_10601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _11389_ (.A1(_10600_),
    .A2(_02695_),
    .B1(_10601_),
    .Y(_10602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11390_ (.A(_10602_),
    .Y(_10603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11391_ (.A(\design_top.core0.SIMM[28] ),
    .Y(_02702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11392_ (.A(_02701_),
    .Y(_10604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11393_ (.A(\design_top.core0.SIMM[28] ),
    .X(_10605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11394_ (.A(_02701_),
    .X(_10606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11395_ (.A1(_02702_),
    .A2(_10604_),
    .B1(_10605_),
    .B2(_10606_),
    .X(_10607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11396_ (.A(_10607_),
    .Y(_10608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11397_ (.A(\design_top.core0.SIMM[25] ),
    .Y(_02720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11398_ (.A(_02719_),
    .Y(_10609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11399_ (.A(_02719_),
    .X(_10610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11400_ (.A1(_02720_),
    .A2(_10609_),
    .B1(\design_top.core0.SIMM[25] ),
    .B2(_10610_),
    .X(_10611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11401_ (.A(_10611_),
    .Y(_10612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11402_ (.A(\design_top.core0.SIMM[24] ),
    .Y(_02726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11403_ (.A(_02725_),
    .Y(_10613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11404_ (.A1(_02726_),
    .A2(_10613_),
    .B1(\design_top.core0.SIMM[24] ),
    .B2(_02725_),
    .X(_10614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11405_ (.A(_10614_),
    .Y(_10615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11406_ (.A(\design_top.core0.SIMM[27] ),
    .Y(_10616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11407_ (.A(_02707_),
    .Y(_10617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11408_ (.A1(\design_top.core0.SIMM[27] ),
    .A2(_02707_),
    .B1(_10616_),
    .B2(_10617_),
    .X(_10618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11409_ (.A(_02713_),
    .X(_10619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11410_ (.A(\design_top.core0.SIMM[26] ),
    .Y(_10620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11411_ (.A(_02713_),
    .Y(_10621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11412_ (.A1(\design_top.core0.SIMM[26] ),
    .A2(_10619_),
    .B1(_10620_),
    .B2(_10621_),
    .X(_10622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11413_ (.A(_10618_),
    .B(_10622_),
    .X(_10623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11414_ (.A(\design_top.core0.SIMM[20] ),
    .Y(_02750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11415_ (.A(_02749_),
    .Y(_10624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11416_ (.A(\design_top.core0.SIMM[20] ),
    .X(_10625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11417_ (.A1(_02750_),
    .A2(_10624_),
    .B1(_10625_),
    .B2(_02749_),
    .X(_10626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11418_ (.A(_10626_),
    .Y(_10627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11419_ (.A(\design_top.core0.SIMM[21] ),
    .Y(_02744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11420_ (.A(_02743_),
    .Y(_10628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11421_ (.A(_02743_),
    .X(_10629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11422_ (.A1(_02744_),
    .A2(_10628_),
    .B1(\design_top.core0.SIMM[21] ),
    .B2(_10629_),
    .X(_10630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11423_ (.A(_10630_),
    .Y(_10631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11424_ (.A(\design_top.core0.SIMM[22] ),
    .Y(_10632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11425_ (.A(_02737_),
    .Y(_10633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11426_ (.A(\design_top.core0.SIMM[22] ),
    .X(_10634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11427_ (.A(_02737_),
    .X(_10635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11428_ (.A1(_10632_),
    .A2(_10633_),
    .B1(_10634_),
    .B2(_10635_),
    .X(_10636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11429_ (.A(_10636_),
    .Y(_10637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11430_ (.A(_02731_),
    .X(_10638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11431_ (.A(\design_top.core0.SIMM[23] ),
    .B(_02731_),
    .Y(_10639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _11432_ (.A1(\design_top.core0.SIMM[23] ),
    .A2(_10638_),
    .B1(_10639_),
    .Y(_10640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11433_ (.A(_10640_),
    .Y(_10641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11434_ (.A(_10627_),
    .B(_10631_),
    .C(_10637_),
    .D(_10641_),
    .X(_10642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11435_ (.A(\design_top.core0.SIMM[18] ),
    .Y(_10643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11436_ (.A(_02761_),
    .Y(_10644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11437_ (.A1(_10643_),
    .A2(_10644_),
    .B1(\design_top.core0.SIMM[18] ),
    .B2(_02761_),
    .X(_10645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11438_ (.A(_10645_),
    .Y(_10646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11439_ (.A(\design_top.core0.SIMM[19] ),
    .B(_02755_),
    .Y(_10647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _11440_ (.A1(\design_top.core0.SIMM[19] ),
    .A2(_02755_),
    .B1(_10647_),
    .Y(_10648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11441_ (.A(_10648_),
    .Y(_10649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11442_ (.A(_02767_),
    .X(_10650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11443_ (.A1(\design_top.core0.SIMM[16] ),
    .A2(_02773_),
    .B1(\design_top.core0.SIMM[17] ),
    .B2(_10650_),
    .X(_10651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11444_ (.A1(\design_top.core0.SIMM[17] ),
    .A2(_10650_),
    .B1(_10651_),
    .Y(_10652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11445_ (.A(_10643_),
    .X(_02762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11446_ (.A(\design_top.core0.SIMM[19] ),
    .X(_10653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11447_ (.A(_10653_),
    .Y(_02756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11448_ (.A(_02755_),
    .Y(_10654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _11449_ (.A1(_02762_),
    .A2(_10644_),
    .A3(_10647_),
    .B1(_02756_),
    .B2(_10654_),
    .X(_10655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _11450_ (.A1(_10646_),
    .A2(_10649_),
    .A3(_10652_),
    .B1(_10655_),
    .X(_10656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11451_ (.A(_02779_),
    .X(_10657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11452_ (.A(\design_top.core0.SIMM[15] ),
    .B(_02779_),
    .Y(_10658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _11453_ (.A1(\design_top.core0.SIMM[15] ),
    .A2(_10657_),
    .B1(_10658_),
    .Y(_10659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11454_ (.A(_10659_),
    .Y(_10660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11455_ (.A(\design_top.core0.SIMM[14] ),
    .Y(_10661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11456_ (.A(_02785_),
    .Y(_10662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11457_ (.A(\design_top.core0.SIMM[14] ),
    .X(_10663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11458_ (.A(_02785_),
    .X(_10664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11459_ (.A1(_10661_),
    .A2(_10662_),
    .B1(_10663_),
    .B2(_10664_),
    .X(_10665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11460_ (.A(_10665_),
    .Y(_10666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11461_ (.A(\design_top.core0.SIMM[13] ),
    .Y(_02792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11462_ (.A(_02791_),
    .Y(_10667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11463_ (.A1(_02792_),
    .A2(_10667_),
    .B1(\design_top.core0.SIMM[13] ),
    .B2(_02791_),
    .X(_10668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11464_ (.A(_10668_),
    .Y(_10669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11465_ (.A(\design_top.core0.SIMM[12] ),
    .Y(_02798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11466_ (.A(_02797_),
    .Y(_10670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11467_ (.A(\design_top.core0.SIMM[12] ),
    .X(_10671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11468_ (.A(_02797_),
    .X(_10672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11469_ (.A1(_02798_),
    .A2(_10670_),
    .B1(_10671_),
    .B2(_10672_),
    .X(_10673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11470_ (.A(_10673_),
    .Y(_10674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11471_ (.A(_10660_),
    .B(_10666_),
    .C(_10669_),
    .D(_10674_),
    .X(_10675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11472_ (.A(_02803_),
    .X(_10676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11473_ (.A(\design_top.core0.SIMM[11] ),
    .B(_02803_),
    .Y(_10677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _11474_ (.A1(\design_top.core0.SIMM[11] ),
    .A2(_10676_),
    .B1(_10677_),
    .Y(_10678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11475_ (.A(_10678_),
    .Y(_10679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11476_ (.A(\design_top.core0.SIMM[10] ),
    .Y(_10680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11477_ (.A(_02809_),
    .Y(_10681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11478_ (.A(_02809_),
    .X(_10682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11479_ (.A1(_10680_),
    .A2(_10681_),
    .B1(\design_top.core0.SIMM[10] ),
    .B2(_10682_),
    .X(_10683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11480_ (.A(_10683_),
    .Y(_10684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11481_ (.A(_02821_),
    .X(_10685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11482_ (.A1(\design_top.core0.SIMM[9] ),
    .A2(_02815_),
    .B1(\design_top.core0.SIMM[8] ),
    .B2(_10685_),
    .X(_10686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11483_ (.A1(\design_top.core0.SIMM[9] ),
    .A2(_02815_),
    .B1(_10686_),
    .Y(_10687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11484_ (.A(_10680_),
    .X(_02810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11485_ (.A(_10681_),
    .X(_03049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11486_ (.A(\design_top.core0.SIMM[11] ),
    .X(_10688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11487_ (.A(_10688_),
    .Y(_02804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11488_ (.A(_10676_),
    .Y(_00803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _11489_ (.A1(_02810_),
    .A2(_03049_),
    .A3(_10677_),
    .B1(_02804_),
    .B2(_00803_),
    .X(_10689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _11490_ (.A1(_10679_),
    .A2(_10684_),
    .A3(_10687_),
    .B1(_10689_),
    .X(_10690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11491_ (.A(_02839_),
    .X(_10691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11492_ (.A(\design_top.core0.SIMM[5] ),
    .Y(_02840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11493_ (.A(_02839_),
    .Y(_00811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11494_ (.A1(\design_top.core0.SIMM[5] ),
    .A2(_10691_),
    .B1(_02840_),
    .B2(_00811_),
    .X(_10692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11495_ (.A(_02845_),
    .X(_10693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11496_ (.A(\design_top.core0.SIMM[4] ),
    .Y(_02846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11497_ (.A(_10693_),
    .Y(_10694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11498_ (.A1(\design_top.core0.SIMM[4] ),
    .A2(_10693_),
    .B1(_02846_),
    .B2(_10694_),
    .X(_10695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11499_ (.A(_02833_),
    .X(_10696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11500_ (.A(\design_top.core0.SIMM[6] ),
    .Y(_02834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11501_ (.A(_02833_),
    .Y(_10697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11502_ (.A1(\design_top.core0.SIMM[6] ),
    .A2(_10696_),
    .B1(_02834_),
    .B2(_10697_),
    .X(_10698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11503_ (.A(\design_top.core0.SIMM[7] ),
    .Y(_02828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11504_ (.A(_02827_),
    .Y(_10699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11505_ (.A1(\design_top.core0.SIMM[7] ),
    .A2(_02827_),
    .B1(_02828_),
    .B2(_10699_),
    .X(_10700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11506_ (.A(_10698_),
    .B(_10700_),
    .X(_10701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11507_ (.A(\design_top.core0.SIMM[3] ),
    .X(_10702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11508_ (.A(\design_top.core0.SIMM[3] ),
    .B(_02659_),
    .Y(_10703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _11509_ (.A1(_10702_),
    .A2(_02659_),
    .B1(_10703_),
    .X(_10704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11510_ (.A(\design_top.core0.SIMM[2] ),
    .Y(_02627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11511_ (.A(_02634_),
    .Y(_10705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11512_ (.A(\design_top.core0.SIMM[2] ),
    .X(_10706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11513_ (.A1(_02627_),
    .A2(_10705_),
    .B1(_10706_),
    .B2(_02634_),
    .X(_10707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11514_ (.A(_10707_),
    .Y(_10708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11515_ (.A(\design_top.core0.SIMM[1] ),
    .X(_10709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11516_ (.A(\design_top.core0.SIMM[0] ),
    .Y(_10710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11517_ (.A(_02650_),
    .Y(_10711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11518_ (.A(_10710_),
    .B(_10711_),
    .Y(_10712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11519_ (.A(\design_top.core0.SIMM[1] ),
    .Y(_02642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11520_ (.A(_02641_),
    .Y(_10713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11521_ (.A1(_02642_),
    .A2(_10713_),
    .B1(\design_top.core0.SIMM[1] ),
    .B2(_02641_),
    .X(_10714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11522_ (.A1(_10709_),
    .A2(_02641_),
    .B1(_10712_),
    .B2(_10714_),
    .X(_10715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11523_ (.A(_10715_),
    .Y(_10716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11524_ (.A(\design_top.core0.SIMM[3] ),
    .Y(_02652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11525_ (.A(_02659_),
    .Y(_10717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _11526_ (.A1(_02627_),
    .A2(_10705_),
    .A3(_10703_),
    .B1(_02652_),
    .B2(_10717_),
    .X(_10718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _11527_ (.A1(_10704_),
    .A2(_10708_),
    .A3(_10716_),
    .B1(_10718_),
    .X(_10719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11528_ (.A1(\design_top.core0.SIMM[5] ),
    .A2(_02839_),
    .B1(\design_top.core0.SIMM[4] ),
    .B2(_02845_),
    .X(_10720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11529_ (.A1(\design_top.core0.SIMM[5] ),
    .A2(_02839_),
    .B1(_10720_),
    .Y(_10721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _11530_ (.A1(_02828_),
    .A2(_10699_),
    .B1(_02834_),
    .C1(_10697_),
    .X(_10722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11531_ (.A1(_02828_),
    .A2(_10699_),
    .B1(_10701_),
    .B2(_10721_),
    .C1(_10722_),
    .X(_10723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o41a_2 _11532_ (.A1(_10692_),
    .A2(_10695_),
    .A3(_10701_),
    .A4(_10719_),
    .B1(_10723_),
    .X(_10724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11533_ (.A(\design_top.core0.SIMM[9] ),
    .Y(_02816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11534_ (.A(_02815_),
    .Y(_00805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11535_ (.A1(_02816_),
    .A2(_00805_),
    .B1(\design_top.core0.SIMM[9] ),
    .B2(_02815_),
    .X(_10725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11536_ (.A(_10725_),
    .Y(_10726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11537_ (.A(\design_top.core0.SIMM[8] ),
    .Y(_02822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11538_ (.A(_02821_),
    .Y(_10727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11539_ (.A1(_02822_),
    .A2(_10727_),
    .B1(\design_top.core0.SIMM[8] ),
    .B2(_02821_),
    .X(_10728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11540_ (.A(_10728_),
    .Y(_10729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11541_ (.A(_10679_),
    .B(_10684_),
    .C(_10726_),
    .D(_10729_),
    .X(_10730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11542_ (.A(_10675_),
    .B(_10730_),
    .X(_10731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11543_ (.A1(\design_top.core0.SIMM[13] ),
    .A2(_02791_),
    .B1(_10671_),
    .B2(_10672_),
    .X(_10732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11544_ (.A1(\design_top.core0.SIMM[13] ),
    .A2(_02791_),
    .B1(_10732_),
    .Y(_10733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11545_ (.A(_10661_),
    .X(_02786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11546_ (.A(_10662_),
    .X(_10734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11547_ (.A(\design_top.core0.SIMM[15] ),
    .X(_10735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11548_ (.A(_10735_),
    .Y(_02780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11549_ (.A(_10657_),
    .Y(_10736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _11550_ (.A1(_02786_),
    .A2(_10734_),
    .A3(_10658_),
    .B1(_02780_),
    .B2(_10736_),
    .X(_10737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _11551_ (.A1(_10660_),
    .A2(_10666_),
    .A3(_10733_),
    .B1(_10737_),
    .X(_10738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11552_ (.A1(_10675_),
    .A2(_10690_),
    .B1(_10724_),
    .B2(_10731_),
    .C1(_10738_),
    .X(_10739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11553_ (.A(\design_top.core0.SIMM[16] ),
    .Y(_02774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11554_ (.A(_02773_),
    .Y(_10740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11555_ (.A1(_02774_),
    .A2(_10740_),
    .B1(\design_top.core0.SIMM[16] ),
    .B2(_02773_),
    .X(_10741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11556_ (.A(_10741_),
    .Y(_10742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11557_ (.A(\design_top.core0.SIMM[17] ),
    .Y(_02768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11558_ (.A(_02767_),
    .Y(_10743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11559_ (.A1(_02768_),
    .A2(_10743_),
    .B1(\design_top.core0.SIMM[17] ),
    .B2(_10650_),
    .X(_10744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11560_ (.A(_10744_),
    .Y(_10745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11561_ (.A(_10742_),
    .B(_10745_),
    .C(_10646_),
    .D(_10649_),
    .X(_10746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11562_ (.A(_10746_),
    .B(_10642_),
    .X(_10747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11563_ (.A1(_10625_),
    .A2(_02749_),
    .B1(\design_top.core0.SIMM[21] ),
    .B2(_10629_),
    .X(_10748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11564_ (.A1(\design_top.core0.SIMM[21] ),
    .A2(_10629_),
    .B1(_10748_),
    .Y(_10749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11565_ (.A(_10632_),
    .X(_02738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11566_ (.A(\design_top.core0.SIMM[23] ),
    .X(_10750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11567_ (.A(_10750_),
    .Y(_02732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11568_ (.A(_10638_),
    .Y(_02939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _11569_ (.A1(_02738_),
    .A2(_10633_),
    .A3(_10639_),
    .B1(_02732_),
    .B2(_02939_),
    .X(_10751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _11570_ (.A1(_10637_),
    .A2(_10641_),
    .A3(_10749_),
    .B1(_10751_),
    .X(_10752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11571_ (.A1(_10642_),
    .A2(_10656_),
    .B1(_10739_),
    .B2(_10747_),
    .C1(_10752_),
    .X(_10753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11572_ (.A(_10616_),
    .X(_02708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11573_ (.A1(\design_top.core0.SIMM[25] ),
    .A2(_10610_),
    .B1(\design_top.core0.SIMM[24] ),
    .B2(_02725_),
    .X(_10754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _11574_ (.A1(\design_top.core0.SIMM[25] ),
    .A2(_10610_),
    .B1(_10754_),
    .Y(_10755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11575_ (.A(_10621_),
    .X(_10756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _11576_ (.A1(_10616_),
    .A2(_10617_),
    .B1(_10620_),
    .C1(_10756_),
    .X(_10757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11577_ (.A1(_02708_),
    .A2(_10617_),
    .B1(_10623_),
    .B2(_10755_),
    .C1(_10757_),
    .X(_10758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o41a_2 _11578_ (.A1(_10612_),
    .A2(_10615_),
    .A3(_10623_),
    .A4(_10753_),
    .B1(_10758_),
    .X(_10759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11579_ (.A(\design_top.core0.SIMM[29] ),
    .Y(_02696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11580_ (.A(_02695_),
    .Y(_10760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _11581_ (.A1(_02702_),
    .A2(_10604_),
    .A3(_10601_),
    .B1(_02696_),
    .B2(_10760_),
    .X(_10761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _11582_ (.A1(_10603_),
    .A2(_10608_),
    .A3(_10759_),
    .B1(_10761_),
    .X(_10762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _11583_ (.A1(_02690_),
    .A2(_10598_),
    .B1(_10599_),
    .B2(_10762_),
    .Y(_10763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11584_ (.A(_02684_),
    .Y(_10764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11585_ (.A(\design_top.core0.SIMM[31] ),
    .Y(_00780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11586_ (.A1(\design_top.core0.SIMM[31] ),
    .A2(_10764_),
    .B1(_00780_),
    .B2(_02684_),
    .X(_10765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11587_ (.A1_N(_10763_),
    .A2_N(_10765_),
    .B1(_10763_),
    .B2(_10765_),
    .X(\design_top.DADDR[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11588_ (.A(_10594_),
    .B(_10596_),
    .C(\design_top.DADDR[31] ),
    .X(_10766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11589_ (.A(_02857_),
    .B(_10766_),
    .X(_10767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11590_ (.A(_10767_),
    .X(_10768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11591_ (.A(_10768_),
    .X(_10769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _11592_ (.A1_N(_10719_),
    .A2_N(_10695_),
    .B1(_10719_),
    .B2(_10695_),
    .X(_01837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11593_ (.A(_10705_),
    .X(_10770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11594_ (.A1(_02627_),
    .A2(_10770_),
    .B1(_10716_),
    .B2(_10708_),
    .X(_10771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11595_ (.A1_N(_10704_),
    .A2_N(_10771_),
    .B1(_10704_),
    .B2(_10771_),
    .X(_10772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11596_ (.A(_10772_),
    .Y(_10773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11597_ (.A(_01837_),
    .B(_10773_),
    .X(_10774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11598_ (.A1(_10716_),
    .A2(_10708_),
    .B1(_10715_),
    .B2(_10707_),
    .X(_10775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11599_ (.A(_10774_),
    .B(_10775_),
    .X(_10776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11600_ (.A(_10694_),
    .X(_03097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11601_ (.A1(_02846_),
    .A2(_03097_),
    .B1(_10719_),
    .B2(_10695_),
    .X(_10777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11602_ (.A1_N(_10692_),
    .A2_N(_10777_),
    .B1(_10692_),
    .B2(_10777_),
    .X(_10778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11603_ (.A(_10778_),
    .Y(_03199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11604_ (.A(_10697_),
    .X(_03081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _11605_ (.A1(_10692_),
    .A2(_10695_),
    .A3(_10719_),
    .B1(_10721_),
    .X(_10779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11606_ (.A1(_02834_),
    .A2(_03081_),
    .B1(_10698_),
    .B2(_10779_),
    .X(_10780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11607_ (.A1_N(_10700_),
    .A2_N(_10780_),
    .B1(_10700_),
    .B2(_10780_),
    .X(_02862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11608_ (.A(_02862_),
    .Y(_01847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11609_ (.A1_N(_10698_),
    .A2_N(_10779_),
    .B1(_10698_),
    .B2(_10779_),
    .X(_02861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11610_ (.A(_02861_),
    .Y(_03216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11611_ (.A(_01847_),
    .B(_03216_),
    .X(_10781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11612_ (.A(_03199_),
    .B(_10781_),
    .X(_10782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11613_ (.A(_10782_),
    .X(_10783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11614_ (.A(_10776_),
    .B(_10783_),
    .X(_10784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11615_ (.A(_10769_),
    .B(_10784_),
    .X(_10785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11616_ (.A(_10785_),
    .X(_10786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11617_ (.A(wbs_adr_i[3]),
    .X(_10787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11618_ (.A(wbs_adr_i[2]),
    .X(_10788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11619_ (.A(wbs_adr_i[1]),
    .X(_10789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11620_ (.A(wbs_adr_i[0]),
    .X(_10790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11621_ (.A(_10787_),
    .B(_10788_),
    .C(_10789_),
    .D(_10790_),
    .X(_10791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11622_ (.A(_10791_),
    .X(_10792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11623_ (.A(_10792_),
    .X(_10793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11624_ (.A(\design_top.XRES ),
    .Y(_10794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11625_ (.A(_10794_),
    .X(_10795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11626_ (.A(wbs_we_i),
    .Y(_10796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _11627_ (.A(_10795_),
    .B(_10796_),
    .C_N(wbs_sel_i[0]),
    .X(_10797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11628_ (.A(_10797_),
    .X(_10798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11629_ (.A(_10798_),
    .X(_10799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11630_ (.A1(_10793_),
    .A2(_10799_),
    .B1(_10785_),
    .X(_10800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11631_ (.A(_10800_),
    .X(_10801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11632_ (.A1_N(_10589_),
    .A2_N(_10786_),
    .B1(\design_top.MEM[0][14] ),
    .B2(_10801_),
    .X(_07430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11633_ (.A(\design_top.DATAO[13] ),
    .Y(_10802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11634_ (.A(_10802_),
    .X(_10803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11635_ (.A(_10803_),
    .X(_10804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11636_ (.A1_N(_10804_),
    .A2_N(_10786_),
    .B1(\design_top.MEM[0][13] ),
    .B2(_10801_),
    .X(_07429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11637_ (.A(\design_top.DATAO[12] ),
    .Y(_10805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11638_ (.A(_10805_),
    .X(_10806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11639_ (.A(_10806_),
    .X(_10807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11640_ (.A1_N(_10807_),
    .A2_N(_10786_),
    .B1(\design_top.MEM[0][12] ),
    .B2(_10801_),
    .X(_07428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11641_ (.A(\design_top.DATAO[11] ),
    .Y(_10808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11642_ (.A(_10808_),
    .X(_10809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11643_ (.A(_10809_),
    .X(_10810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11644_ (.A1_N(_10810_),
    .A2_N(_10786_),
    .B1(\design_top.MEM[0][11] ),
    .B2(_10801_),
    .X(_07427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11645_ (.A(\design_top.DATAO[10] ),
    .Y(_10811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11646_ (.A(_10811_),
    .X(_10812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11647_ (.A(_10812_),
    .X(_10813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11648_ (.A1_N(_10813_),
    .A2_N(_10786_),
    .B1(\design_top.MEM[0][10] ),
    .B2(_10801_),
    .X(_07426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11649_ (.A(\design_top.DATAO[9] ),
    .Y(_10814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11650_ (.A(_10814_),
    .X(_10815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11651_ (.A(_10815_),
    .X(_10816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11652_ (.A1_N(_10816_),
    .A2_N(_10785_),
    .B1(\design_top.MEM[0][9] ),
    .B2(_10800_),
    .X(_07425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11653_ (.A(\design_top.DATAO[8] ),
    .Y(_10817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11654_ (.A(_10817_),
    .X(_10818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11655_ (.A(_10818_),
    .X(_10819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11656_ (.A1_N(_10819_),
    .A2_N(_10785_),
    .B1(\design_top.MEM[0][8] ),
    .B2(_10800_),
    .X(_07424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11657_ (.A(_10775_),
    .X(\design_top.DADDR[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11658_ (.A(\design_top.DATAO[31] ),
    .Y(_10820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11659_ (.A(_10714_),
    .Y(_10821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11660_ (.A(_10710_),
    .X(_02643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11661_ (.A(_10711_),
    .X(_10822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _11662_ (.A1(_02643_),
    .A2(_10822_),
    .B1(_10712_),
    .Y(_10823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11663_ (.A(_10823_),
    .Y(_10824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11664_ (.A(_10821_),
    .B(_10824_),
    .X(_10825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11665_ (.A(_10820_),
    .B(_10825_),
    .X(_10826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11666_ (.A(_10773_),
    .X(\design_top.DADDR[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11667_ (.A(\design_top.DADDR[31] ),
    .Y(_10827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11668_ (.A(_10596_),
    .B(_10827_),
    .X(_10828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11669_ (.A(\design_top.DADDR[2] ),
    .B(_10826_),
    .C(\design_top.DADDR[3] ),
    .D(_10828_),
    .X(_10829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11670_ (.A(_10829_),
    .Y(_10830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11671_ (.A(\design_top.IRES[7] ),
    .Y(_10831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11672_ (.A(_10831_),
    .X(_10832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11673_ (.A(_10832_),
    .X(_10833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11674_ (.A1(\design_top.IREQ[7] ),
    .A2(_10829_),
    .B1(\design_top.IACK[7] ),
    .B2(_10830_),
    .C1(_10833_),
    .X(_07423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11675_ (.A(\design_top.IOMUX[3][11] ),
    .B(\design_top.IOMUX[3][10] ),
    .C(\design_top.IOMUX[3][9] ),
    .D(\design_top.IOMUX[3][8] ),
    .X(_10834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11676_ (.A(\design_top.IOMUX[3][15] ),
    .B(\design_top.IOMUX[3][14] ),
    .C(\design_top.IOMUX[3][13] ),
    .D(\design_top.IOMUX[3][12] ),
    .X(_10835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11677_ (.A(\design_top.IOMUX[3][3] ),
    .B(\design_top.IOMUX[3][2] ),
    .C(\design_top.IOMUX[3][1] ),
    .D(\design_top.IOMUX[3][0] ),
    .X(_10836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11678_ (.A(\design_top.IOMUX[3][7] ),
    .B(\design_top.IOMUX[3][6] ),
    .C(\design_top.IOMUX[3][5] ),
    .D(\design_top.IOMUX[3][4] ),
    .X(_10837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11679_ (.A(_10834_),
    .B(_10835_),
    .C(_10836_),
    .D(_10837_),
    .X(_10838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11680_ (.A(\design_top.IOMUX[3][27] ),
    .B(\design_top.IOMUX[3][26] ),
    .C(\design_top.IOMUX[3][25] ),
    .D(\design_top.IOMUX[3][24] ),
    .X(_10839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11681_ (.A(\design_top.IOMUX[3][31] ),
    .B(\design_top.IOMUX[3][30] ),
    .C(\design_top.IOMUX[3][29] ),
    .D(\design_top.IOMUX[3][28] ),
    .X(_10840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11682_ (.A(\design_top.IOMUX[3][19] ),
    .B(\design_top.IOMUX[3][18] ),
    .C(\design_top.IOMUX[3][17] ),
    .D(\design_top.IOMUX[3][16] ),
    .X(_10841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11683_ (.A(\design_top.IOMUX[3][23] ),
    .B(\design_top.IOMUX[3][22] ),
    .C(\design_top.IOMUX[3][21] ),
    .D(\design_top.IOMUX[3][20] ),
    .X(_10842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11684_ (.A(_10839_),
    .B(_10840_),
    .C(_10841_),
    .D(_10842_),
    .X(_10843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11685_ (.A(_10838_),
    .B(_10843_),
    .Y(_10844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11686_ (.A(\design_top.TIMER[31] ),
    .B(\design_top.TIMER[30] ),
    .X(_10845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11687_ (.A(\design_top.TIMER[19] ),
    .B(\design_top.TIMER[18] ),
    .X(_10846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11688_ (.A(\design_top.TIMER[1] ),
    .B(\design_top.TIMER[0] ),
    .X(_10847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11689_ (.A(\design_top.TIMER[2] ),
    .B(_10847_),
    .X(_10848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11690_ (.A(\design_top.TIMER[3] ),
    .B(_10848_),
    .X(_10849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11691_ (.A(\design_top.TIMER[4] ),
    .B(_10849_),
    .X(_10850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11692_ (.A(\design_top.TIMER[5] ),
    .B(_10850_),
    .X(_10851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11693_ (.A(\design_top.TIMER[6] ),
    .B(_10851_),
    .X(_10852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11694_ (.A(\design_top.TIMER[7] ),
    .B(_10852_),
    .X(_10853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11695_ (.A(\design_top.TIMER[8] ),
    .B(_10853_),
    .X(_10854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11696_ (.A(\design_top.TIMER[9] ),
    .B(_10854_),
    .X(_10855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11697_ (.A(\design_top.TIMER[10] ),
    .B(_10855_),
    .X(_10856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11698_ (.A(\design_top.TIMER[11] ),
    .B(_10856_),
    .X(_10857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11699_ (.A(\design_top.TIMER[12] ),
    .B(_10857_),
    .X(_10858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11700_ (.A(\design_top.TIMER[13] ),
    .B(_10858_),
    .X(_10859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11701_ (.A(\design_top.TIMER[14] ),
    .B(_10859_),
    .X(_10860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11702_ (.A(\design_top.TIMER[15] ),
    .B(_10860_),
    .X(_10861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11703_ (.A(\design_top.TIMER[17] ),
    .B(\design_top.TIMER[16] ),
    .C(_10846_),
    .D(_10861_),
    .X(_10862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11704_ (.A(\design_top.TIMER[21] ),
    .B(\design_top.TIMER[20] ),
    .C(_10862_),
    .X(_10863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11705_ (.A(\design_top.TIMER[23] ),
    .B(\design_top.TIMER[22] ),
    .C(_10863_),
    .X(_10864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11706_ (.A(\design_top.TIMER[25] ),
    .B(\design_top.TIMER[24] ),
    .C(_10864_),
    .X(_10865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11707_ (.A(\design_top.TIMER[26] ),
    .B(_10865_),
    .X(_10866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11708_ (.A(\design_top.TIMER[27] ),
    .B(_10866_),
    .X(_10867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11709_ (.A(\design_top.TIMER[29] ),
    .B(\design_top.TIMER[28] ),
    .C(_10845_),
    .D(_10867_),
    .X(_10868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11710_ (.A(_10844_),
    .B(_10868_),
    .X(_10869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11711_ (.A(_10869_),
    .Y(_10870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11712_ (.A(\design_top.IACK[7] ),
    .Y(_10871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11713_ (.A(_10831_),
    .X(_10872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11714_ (.A(_10872_),
    .X(_10873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _11715_ (.A1(\design_top.IREQ[7] ),
    .A2(_10870_),
    .B1(_10871_),
    .B2(_10869_),
    .C1(_10873_),
    .X(_07422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11716_ (.A(\design_top.DATAO[23] ),
    .Y(_10874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11717_ (.A(_10874_),
    .X(_10875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11718_ (.A(_10875_),
    .X(_10876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11719_ (.A(_02865_),
    .B(_10766_),
    .X(_10877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11720_ (.A(_10877_),
    .X(_10878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11721_ (.A(_10878_),
    .X(_10879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11722_ (.A(_10778_),
    .X(_02860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11723_ (.A(_01847_),
    .B(_02861_),
    .X(_10880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11724_ (.A(_02860_),
    .B(_10880_),
    .X(_10881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11725_ (.A(_10775_),
    .Y(_10882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11726_ (.A(_10882_),
    .X(_02651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11727_ (.A(_01837_),
    .B(_10772_),
    .X(_10883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11728_ (.A(_02651_),
    .B(_10883_),
    .X(_10884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11729_ (.A(_10884_),
    .X(_10885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11730_ (.A(_10881_),
    .B(_10885_),
    .X(_10886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11731_ (.A(_10879_),
    .B(_10886_),
    .X(_10887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11732_ (.A(_10887_),
    .X(_10888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _11733_ (.A(_10794_),
    .B(_10796_),
    .C_N(wbs_sel_i[3]),
    .X(_10889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11734_ (.A(_10889_),
    .X(_10890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11735_ (.A(_10890_),
    .X(_10891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11736_ (.A(_10891_),
    .X(_10892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11737_ (.A(wbs_adr_i[2]),
    .Y(_10893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11738_ (.A(_10893_),
    .X(_10894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11739_ (.A(wbs_adr_i[1]),
    .Y(_10895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11740_ (.A(_10895_),
    .X(_10896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11741_ (.A(_10787_),
    .B(_10894_),
    .C(_10896_),
    .D(_10790_),
    .X(_10897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11742_ (.A(_10897_),
    .X(_10898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11743_ (.A(_10898_),
    .X(_10899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11744_ (.A1(_10892_),
    .A2(_10899_),
    .B1(_10887_),
    .X(_10900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11745_ (.A(_10900_),
    .X(_10901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11746_ (.A1_N(_10876_),
    .A2_N(_10888_),
    .B1(\design_top.MEM[27][23] ),
    .B2(_10901_),
    .X(_07421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11747_ (.A(\design_top.DATAO[22] ),
    .Y(_10902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11748_ (.A(_10902_),
    .X(_10903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11749_ (.A(_10903_),
    .X(_10904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11750_ (.A1_N(_10904_),
    .A2_N(_10888_),
    .B1(\design_top.MEM[27][22] ),
    .B2(_10901_),
    .X(_07420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11751_ (.A(\design_top.DATAO[21] ),
    .Y(_10905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11752_ (.A(_10905_),
    .X(_10906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11753_ (.A(_10906_),
    .X(_10907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11754_ (.A1_N(_10907_),
    .A2_N(_10888_),
    .B1(\design_top.MEM[27][21] ),
    .B2(_10901_),
    .X(_07419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11755_ (.A(\design_top.DATAO[20] ),
    .Y(_10908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11756_ (.A(_10908_),
    .X(_10909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11757_ (.A(_10909_),
    .X(_10910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11758_ (.A1_N(_10910_),
    .A2_N(_10888_),
    .B1(\design_top.MEM[27][20] ),
    .B2(_10901_),
    .X(_07418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11759_ (.A(\design_top.DATAO[19] ),
    .Y(_10911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11760_ (.A(_10911_),
    .X(_10912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11761_ (.A(_10912_),
    .X(_10913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11762_ (.A1_N(_10913_),
    .A2_N(_10888_),
    .B1(\design_top.MEM[27][19] ),
    .B2(_10901_),
    .X(_07417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11763_ (.A(\design_top.DATAO[18] ),
    .Y(_10914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11764_ (.A(_10914_),
    .X(_10915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11765_ (.A(_10915_),
    .X(_10916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11766_ (.A1_N(_10916_),
    .A2_N(_10887_),
    .B1(\design_top.MEM[27][18] ),
    .B2(_10900_),
    .X(_07416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11767_ (.A(\design_top.DATAO[17] ),
    .Y(_10917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11768_ (.A(_10917_),
    .X(_10918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11769_ (.A(_10918_),
    .X(_10919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11770_ (.A1_N(_10919_),
    .A2_N(_10887_),
    .B1(\design_top.MEM[27][17] ),
    .B2(_10900_),
    .X(_07415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11771_ (.A(\design_top.DATAO[16] ),
    .Y(_10920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11772_ (.A(_10920_),
    .X(_10921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11773_ (.A(_10921_),
    .X(_10922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11774_ (.A1_N(_10922_),
    .A2_N(_10887_),
    .B1(\design_top.MEM[27][16] ),
    .B2(_10900_),
    .X(_07414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11775_ (.A(_10820_),
    .X(_10923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11776_ (.A(_10923_),
    .X(_10924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11777_ (.A(_02868_),
    .B(_10766_),
    .X(_10925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11778_ (.A(_10925_),
    .X(_10926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11779_ (.A(_10926_),
    .X(_10927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11780_ (.A(_10886_),
    .B(_10927_),
    .X(_10928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11781_ (.A(_10928_),
    .X(_10929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11782_ (.A1(_10892_),
    .A2(_10899_),
    .B1(_10928_),
    .X(_10930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11783_ (.A(_10930_),
    .X(_10931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11784_ (.A1_N(_10924_),
    .A2_N(_10929_),
    .B1(\design_top.MEM[27][31] ),
    .B2(_10931_),
    .X(_07413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11785_ (.A(\design_top.DATAO[30] ),
    .Y(_10932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11786_ (.A(_10932_),
    .X(_10933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11787_ (.A(_10933_),
    .X(_10934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11788_ (.A1_N(_10934_),
    .A2_N(_10929_),
    .B1(\design_top.MEM[27][30] ),
    .B2(_10931_),
    .X(_07412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11789_ (.A(\design_top.DATAO[29] ),
    .Y(_10935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11790_ (.A(_10935_),
    .X(_10936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11791_ (.A(_10936_),
    .X(_10937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11792_ (.A1_N(_10937_),
    .A2_N(_10929_),
    .B1(\design_top.MEM[27][29] ),
    .B2(_10931_),
    .X(_07411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11793_ (.A(\design_top.DATAO[28] ),
    .Y(_10938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11794_ (.A(_10938_),
    .X(_10939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11795_ (.A(_10939_),
    .X(_10940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11796_ (.A1_N(_10940_),
    .A2_N(_10929_),
    .B1(\design_top.MEM[27][28] ),
    .B2(_10931_),
    .X(_07410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11797_ (.A(\design_top.DATAO[27] ),
    .Y(_10941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11798_ (.A(_10941_),
    .X(_10942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11799_ (.A(_10942_),
    .X(_10943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11800_ (.A1_N(_10943_),
    .A2_N(_10929_),
    .B1(\design_top.MEM[27][27] ),
    .B2(_10931_),
    .X(_07409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11801_ (.A(\design_top.DATAO[26] ),
    .Y(_10944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11802_ (.A(_10944_),
    .X(_10945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11803_ (.A(_10945_),
    .X(_10946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11804_ (.A1_N(_10946_),
    .A2_N(_10928_),
    .B1(\design_top.MEM[27][26] ),
    .B2(_10930_),
    .X(_07408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11805_ (.A(\design_top.DATAO[25] ),
    .Y(_10947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11806_ (.A(_10947_),
    .X(_10948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11807_ (.A(_10948_),
    .X(_10949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11808_ (.A1_N(_10949_),
    .A2_N(_10928_),
    .B1(\design_top.MEM[27][25] ),
    .B2(_10930_),
    .X(_07407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11809_ (.A(\design_top.DATAO[24] ),
    .Y(_10950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11810_ (.A(_10950_),
    .X(_10951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11811_ (.A(_10951_),
    .X(_10952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11812_ (.A1_N(_10952_),
    .A2_N(_10928_),
    .B1(\design_top.MEM[27][24] ),
    .B2(_10930_),
    .X(_07406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11813_ (.A(\design_top.DATAO[15] ),
    .Y(_10953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11814_ (.A(_10953_),
    .X(_10954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11815_ (.A(_10954_),
    .X(_10955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11816_ (.A(_10881_),
    .X(_10956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11817_ (.A(_01837_),
    .Y(_02859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11818_ (.A(_02859_),
    .B(_10775_),
    .C(\design_top.DADDR[3] ),
    .X(_10957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11819_ (.A(_10957_),
    .X(_10958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11820_ (.A(_10956_),
    .B(_10958_),
    .X(_10959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11821_ (.A(_10769_),
    .B(_10959_),
    .X(_10960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11822_ (.A(_10960_),
    .X(_10961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11823_ (.A(_10799_),
    .X(_10962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11824_ (.A(wbs_adr_i[0]),
    .Y(_10963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11825_ (.A(_10963_),
    .X(_10964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11826_ (.A(_10787_),
    .B(_10894_),
    .C(_10896_),
    .D(_10964_),
    .X(_10965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11827_ (.A(_10965_),
    .X(_10966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11828_ (.A(_10966_),
    .X(_10967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11829_ (.A1(_10962_),
    .A2(_10967_),
    .B1(_10960_),
    .X(_10968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11830_ (.A(_10968_),
    .X(_10969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11831_ (.A1_N(_10955_),
    .A2_N(_10961_),
    .B1(\design_top.MEM[28][15] ),
    .B2(_10969_),
    .X(_07405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11832_ (.A1_N(_10589_),
    .A2_N(_10961_),
    .B1(\design_top.MEM[28][14] ),
    .B2(_10969_),
    .X(_07404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11833_ (.A1_N(_10804_),
    .A2_N(_10961_),
    .B1(\design_top.MEM[28][13] ),
    .B2(_10969_),
    .X(_07403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11834_ (.A1_N(_10807_),
    .A2_N(_10961_),
    .B1(\design_top.MEM[28][12] ),
    .B2(_10969_),
    .X(_07402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11835_ (.A1_N(_10810_),
    .A2_N(_10961_),
    .B1(\design_top.MEM[28][11] ),
    .B2(_10969_),
    .X(_07401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11836_ (.A1_N(_10813_),
    .A2_N(_10960_),
    .B1(\design_top.MEM[28][10] ),
    .B2(_10968_),
    .X(_07400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11837_ (.A1_N(_10816_),
    .A2_N(_10960_),
    .B1(\design_top.MEM[28][9] ),
    .B2(_10968_),
    .X(_07399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11838_ (.A1_N(_10819_),
    .A2_N(_10960_),
    .B1(\design_top.MEM[28][8] ),
    .B2(_10968_),
    .X(_07398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11839_ (.A(_10879_),
    .B(_10959_),
    .X(_10970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11840_ (.A(_10970_),
    .X(_10971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11841_ (.A1(_10962_),
    .A2(_10967_),
    .B1(_10970_),
    .X(_10972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11842_ (.A(_10972_),
    .X(_10973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11843_ (.A1_N(_10876_),
    .A2_N(_10971_),
    .B1(\design_top.MEM[28][23] ),
    .B2(_10973_),
    .X(_07397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11844_ (.A1_N(_10904_),
    .A2_N(_10971_),
    .B1(\design_top.MEM[28][22] ),
    .B2(_10973_),
    .X(_07396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11845_ (.A1_N(_10907_),
    .A2_N(_10971_),
    .B1(\design_top.MEM[28][21] ),
    .B2(_10973_),
    .X(_07395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11846_ (.A1_N(_10910_),
    .A2_N(_10971_),
    .B1(\design_top.MEM[28][20] ),
    .B2(_10973_),
    .X(_07394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11847_ (.A1_N(_10913_),
    .A2_N(_10971_),
    .B1(\design_top.MEM[28][19] ),
    .B2(_10973_),
    .X(_07393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11848_ (.A1_N(_10916_),
    .A2_N(_10970_),
    .B1(\design_top.MEM[28][18] ),
    .B2(_10972_),
    .X(_07392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11849_ (.A1_N(_10919_),
    .A2_N(_10970_),
    .B1(\design_top.MEM[28][17] ),
    .B2(_10972_),
    .X(_07391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11850_ (.A1_N(_10922_),
    .A2_N(_10970_),
    .B1(\design_top.MEM[28][16] ),
    .B2(_10972_),
    .X(_07390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11851_ (.A(_10927_),
    .B(_10959_),
    .X(_10974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11852_ (.A(_10974_),
    .X(_10975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11853_ (.A1(_10962_),
    .A2(_10967_),
    .B1(_10974_),
    .X(_10976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11854_ (.A(_10976_),
    .X(_10977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11855_ (.A1_N(_10924_),
    .A2_N(_10975_),
    .B1(\design_top.MEM[28][31] ),
    .B2(_10977_),
    .X(_07389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11856_ (.A1_N(_10934_),
    .A2_N(_10975_),
    .B1(\design_top.MEM[28][30] ),
    .B2(_10977_),
    .X(_07388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11857_ (.A1_N(_10937_),
    .A2_N(_10975_),
    .B1(\design_top.MEM[28][29] ),
    .B2(_10977_),
    .X(_07387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11858_ (.A1_N(_10940_),
    .A2_N(_10975_),
    .B1(\design_top.MEM[28][28] ),
    .B2(_10977_),
    .X(_07386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11859_ (.A1_N(_10943_),
    .A2_N(_10975_),
    .B1(\design_top.MEM[28][27] ),
    .B2(_10977_),
    .X(_07385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11860_ (.A1_N(_10946_),
    .A2_N(_10974_),
    .B1(\design_top.MEM[28][26] ),
    .B2(_10976_),
    .X(_07384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11861_ (.A1_N(_10949_),
    .A2_N(_10974_),
    .B1(\design_top.MEM[28][25] ),
    .B2(_10976_),
    .X(_07383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11862_ (.A1_N(_10952_),
    .A2_N(_10974_),
    .B1(\design_top.MEM[28][24] ),
    .B2(_10976_),
    .X(_07382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11863_ (.A(_02859_),
    .B(_10882_),
    .X(_10978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11864_ (.A(\design_top.DADDR[3] ),
    .B(_10978_),
    .X(_10979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11865_ (.A(_10979_),
    .X(_10980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11866_ (.A(_10956_),
    .B(_10980_),
    .X(_10981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11867_ (.A(_10769_),
    .B(_10981_),
    .X(_10982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11868_ (.A(_10982_),
    .X(_10983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11869_ (.A(_10966_),
    .X(_10984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _11870_ (.A(_10794_),
    .B(_10796_),
    .C_N(wbs_sel_i[1]),
    .X(_10985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11871_ (.A(_10985_),
    .X(_10986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11872_ (.A(_10986_),
    .X(_10987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11873_ (.A1(_10984_),
    .A2(_10987_),
    .B1(_10982_),
    .X(_10988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11874_ (.A(_10988_),
    .X(_10989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11875_ (.A1_N(_10955_),
    .A2_N(_10983_),
    .B1(\design_top.MEM[29][15] ),
    .B2(_10989_),
    .X(_07381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11876_ (.A1_N(_10589_),
    .A2_N(_10983_),
    .B1(\design_top.MEM[29][14] ),
    .B2(_10989_),
    .X(_07380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11877_ (.A1_N(_10804_),
    .A2_N(_10983_),
    .B1(\design_top.MEM[29][13] ),
    .B2(_10989_),
    .X(_07379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11878_ (.A1_N(_10807_),
    .A2_N(_10983_),
    .B1(\design_top.MEM[29][12] ),
    .B2(_10989_),
    .X(_07378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11879_ (.A1_N(_10810_),
    .A2_N(_10983_),
    .B1(\design_top.MEM[29][11] ),
    .B2(_10989_),
    .X(_07377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11880_ (.A1_N(_10813_),
    .A2_N(_10982_),
    .B1(\design_top.MEM[29][10] ),
    .B2(_10988_),
    .X(_07376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11881_ (.A1_N(_10816_),
    .A2_N(_10982_),
    .B1(\design_top.MEM[29][9] ),
    .B2(_10988_),
    .X(_07375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11882_ (.A1_N(_10819_),
    .A2_N(_10982_),
    .B1(\design_top.MEM[29][8] ),
    .B2(_10988_),
    .X(_07374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11883_ (.A(_10879_),
    .B(_10981_),
    .X(_10990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11884_ (.A(_10990_),
    .X(_10991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11885_ (.A(_10986_),
    .X(_10992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11886_ (.A1(_10984_),
    .A2(_10992_),
    .B1(_10990_),
    .X(_10993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11887_ (.A(_10993_),
    .X(_10994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11888_ (.A1_N(_10876_),
    .A2_N(_10991_),
    .B1(\design_top.MEM[29][23] ),
    .B2(_10994_),
    .X(_07373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11889_ (.A1_N(_10904_),
    .A2_N(_10991_),
    .B1(\design_top.MEM[29][22] ),
    .B2(_10994_),
    .X(_07372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11890_ (.A1_N(_10907_),
    .A2_N(_10991_),
    .B1(\design_top.MEM[29][21] ),
    .B2(_10994_),
    .X(_07371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11891_ (.A1_N(_10910_),
    .A2_N(_10991_),
    .B1(\design_top.MEM[29][20] ),
    .B2(_10994_),
    .X(_07370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11892_ (.A1_N(_10913_),
    .A2_N(_10991_),
    .B1(\design_top.MEM[29][19] ),
    .B2(_10994_),
    .X(_07369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11893_ (.A1_N(_10916_),
    .A2_N(_10990_),
    .B1(\design_top.MEM[29][18] ),
    .B2(_10993_),
    .X(_07368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11894_ (.A1_N(_10919_),
    .A2_N(_10990_),
    .B1(\design_top.MEM[29][17] ),
    .B2(_10993_),
    .X(_07367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11895_ (.A1_N(_10922_),
    .A2_N(_10990_),
    .B1(\design_top.MEM[29][16] ),
    .B2(_10993_),
    .X(_07366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11896_ (.A(_10927_),
    .B(_10981_),
    .X(_10995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11897_ (.A(_10995_),
    .X(_10996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11898_ (.A1(_10984_),
    .A2(_10992_),
    .B1(_10995_),
    .X(_10997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11899_ (.A(_10997_),
    .X(_10998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11900_ (.A1_N(_10924_),
    .A2_N(_10996_),
    .B1(\design_top.MEM[29][31] ),
    .B2(_10998_),
    .X(_07365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11901_ (.A1_N(_10934_),
    .A2_N(_10996_),
    .B1(\design_top.MEM[29][30] ),
    .B2(_10998_),
    .X(_07364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11902_ (.A1_N(_10937_),
    .A2_N(_10996_),
    .B1(\design_top.MEM[29][29] ),
    .B2(_10998_),
    .X(_07363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11903_ (.A1_N(_10940_),
    .A2_N(_10996_),
    .B1(\design_top.MEM[29][28] ),
    .B2(_10998_),
    .X(_07362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11904_ (.A1_N(_10943_),
    .A2_N(_10996_),
    .B1(\design_top.MEM[29][27] ),
    .B2(_10998_),
    .X(_07361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11905_ (.A1_N(_10946_),
    .A2_N(_10995_),
    .B1(\design_top.MEM[29][26] ),
    .B2(_10997_),
    .X(_07360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11906_ (.A1_N(_10949_),
    .A2_N(_10995_),
    .B1(\design_top.MEM[29][25] ),
    .B2(_10997_),
    .X(_07359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11907_ (.A1_N(_10952_),
    .A2_N(_10995_),
    .B1(\design_top.MEM[29][24] ),
    .B2(_10997_),
    .X(_07358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11908_ (.A(\design_top.DADDR[2] ),
    .B(_10883_),
    .X(_10999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11909_ (.A(_10999_),
    .X(_11000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11910_ (.A(_10783_),
    .B(_11000_),
    .X(_11001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11911_ (.A(_10769_),
    .B(_11001_),
    .X(_11002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11912_ (.A(_11002_),
    .X(_11003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _11913_ (.A(_10794_),
    .B(_10796_),
    .C_N(wbs_sel_i[2]),
    .X(_11004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11914_ (.A(_11004_),
    .X(_11005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11915_ (.A(_11005_),
    .X(_11006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11916_ (.A1(_10793_),
    .A2(_11006_),
    .B1(_11002_),
    .X(_11007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11917_ (.A(_11007_),
    .X(_11008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11918_ (.A1_N(_10955_),
    .A2_N(_11003_),
    .B1(\design_top.MEM[2][15] ),
    .B2(_11008_),
    .X(_07357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11919_ (.A1_N(_10589_),
    .A2_N(_11003_),
    .B1(\design_top.MEM[2][14] ),
    .B2(_11008_),
    .X(_07356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11920_ (.A1_N(_10804_),
    .A2_N(_11003_),
    .B1(\design_top.MEM[2][13] ),
    .B2(_11008_),
    .X(_07355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11921_ (.A1_N(_10807_),
    .A2_N(_11003_),
    .B1(\design_top.MEM[2][12] ),
    .B2(_11008_),
    .X(_07354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11922_ (.A1_N(_10810_),
    .A2_N(_11003_),
    .B1(\design_top.MEM[2][11] ),
    .B2(_11008_),
    .X(_07353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11923_ (.A1_N(_10813_),
    .A2_N(_11002_),
    .B1(\design_top.MEM[2][10] ),
    .B2(_11007_),
    .X(_07352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11924_ (.A1_N(_10816_),
    .A2_N(_11002_),
    .B1(\design_top.MEM[2][9] ),
    .B2(_11007_),
    .X(_07351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11925_ (.A1_N(_10819_),
    .A2_N(_11002_),
    .B1(\design_top.MEM[2][8] ),
    .B2(_11007_),
    .X(_07350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11926_ (.A(_10879_),
    .B(_11001_),
    .X(_11009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11927_ (.A(_11009_),
    .X(_11010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11928_ (.A(_11005_),
    .X(_11011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11929_ (.A1(_10793_),
    .A2(_11011_),
    .B1(_11009_),
    .X(_11012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11930_ (.A(_11012_),
    .X(_11013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11931_ (.A1_N(_10876_),
    .A2_N(_11010_),
    .B1(\design_top.MEM[2][23] ),
    .B2(_11013_),
    .X(_07349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11932_ (.A1_N(_10904_),
    .A2_N(_11010_),
    .B1(\design_top.MEM[2][22] ),
    .B2(_11013_),
    .X(_07348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11933_ (.A1_N(_10907_),
    .A2_N(_11010_),
    .B1(\design_top.MEM[2][21] ),
    .B2(_11013_),
    .X(_07347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11934_ (.A1_N(_10910_),
    .A2_N(_11010_),
    .B1(\design_top.MEM[2][20] ),
    .B2(_11013_),
    .X(_07346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11935_ (.A1_N(_10913_),
    .A2_N(_11010_),
    .B1(\design_top.MEM[2][19] ),
    .B2(_11013_),
    .X(_07345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11936_ (.A1_N(_10916_),
    .A2_N(_11009_),
    .B1(\design_top.MEM[2][18] ),
    .B2(_11012_),
    .X(_07344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11937_ (.A1_N(_10919_),
    .A2_N(_11009_),
    .B1(\design_top.MEM[2][17] ),
    .B2(_11012_),
    .X(_07343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11938_ (.A1_N(_10922_),
    .A2_N(_11009_),
    .B1(\design_top.MEM[2][16] ),
    .B2(_11012_),
    .X(_07342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11939_ (.A(_10927_),
    .B(_11001_),
    .X(_11014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11940_ (.A(_11014_),
    .X(_11015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11941_ (.A1(_10793_),
    .A2(_11011_),
    .B1(_11014_),
    .X(_11016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11942_ (.A(_11016_),
    .X(_11017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11943_ (.A1_N(_10924_),
    .A2_N(_11015_),
    .B1(\design_top.MEM[2][31] ),
    .B2(_11017_),
    .X(_07341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11944_ (.A1_N(_10934_),
    .A2_N(_11015_),
    .B1(\design_top.MEM[2][30] ),
    .B2(_11017_),
    .X(_07340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11945_ (.A1_N(_10937_),
    .A2_N(_11015_),
    .B1(\design_top.MEM[2][29] ),
    .B2(_11017_),
    .X(_07339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11946_ (.A1_N(_10940_),
    .A2_N(_11015_),
    .B1(\design_top.MEM[2][28] ),
    .B2(_11017_),
    .X(_07338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11947_ (.A1_N(_10943_),
    .A2_N(_11015_),
    .B1(\design_top.MEM[2][27] ),
    .B2(_11017_),
    .X(_07337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11948_ (.A1_N(_10946_),
    .A2_N(_11014_),
    .B1(\design_top.MEM[2][26] ),
    .B2(_11016_),
    .X(_07336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11949_ (.A1_N(_10949_),
    .A2_N(_11014_),
    .B1(\design_top.MEM[2][25] ),
    .B2(_11016_),
    .X(_07335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11950_ (.A1_N(_10952_),
    .A2_N(_11014_),
    .B1(\design_top.MEM[2][24] ),
    .B2(_11016_),
    .X(_07334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11951_ (.A(_10772_),
    .X(_02660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _11952_ (.A(_02660_),
    .B(_10775_),
    .C(_02859_),
    .X(_11018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11953_ (.A(_11018_),
    .X(_11019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11954_ (.A(_10956_),
    .B(_11019_),
    .X(_11020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11955_ (.A(_10769_),
    .B(_11020_),
    .X(_11021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11956_ (.A(_11021_),
    .X(_11022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11957_ (.A1(_10984_),
    .A2(_11011_),
    .B1(_11021_),
    .X(_11023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11958_ (.A(_11023_),
    .X(_11024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11959_ (.A1_N(_10955_),
    .A2_N(_11022_),
    .B1(\design_top.MEM[30][15] ),
    .B2(_11024_),
    .X(_07333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11960_ (.A1_N(_10589_),
    .A2_N(_11022_),
    .B1(\design_top.MEM[30][14] ),
    .B2(_11024_),
    .X(_07332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11961_ (.A1_N(_10804_),
    .A2_N(_11022_),
    .B1(\design_top.MEM[30][13] ),
    .B2(_11024_),
    .X(_07331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11962_ (.A1_N(_10807_),
    .A2_N(_11022_),
    .B1(\design_top.MEM[30][12] ),
    .B2(_11024_),
    .X(_07330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11963_ (.A1_N(_10810_),
    .A2_N(_11022_),
    .B1(\design_top.MEM[30][11] ),
    .B2(_11024_),
    .X(_07329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11964_ (.A1_N(_10813_),
    .A2_N(_11021_),
    .B1(\design_top.MEM[30][10] ),
    .B2(_11023_),
    .X(_07328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11965_ (.A1_N(_10816_),
    .A2_N(_11021_),
    .B1(\design_top.MEM[30][9] ),
    .B2(_11023_),
    .X(_07327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11966_ (.A1_N(_10819_),
    .A2_N(_11021_),
    .B1(\design_top.MEM[30][8] ),
    .B2(_11023_),
    .X(_07326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11967_ (.A(_10877_),
    .X(_11025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11968_ (.A(_11025_),
    .X(_11026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11969_ (.A(_11026_),
    .B(_11020_),
    .X(_11027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11970_ (.A(_11027_),
    .X(_11028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11971_ (.A1(_10984_),
    .A2(_11011_),
    .B1(_11027_),
    .X(_11029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11972_ (.A(_11029_),
    .X(_11030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11973_ (.A1_N(_10876_),
    .A2_N(_11028_),
    .B1(\design_top.MEM[30][23] ),
    .B2(_11030_),
    .X(_07325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11974_ (.A1_N(_10904_),
    .A2_N(_11028_),
    .B1(\design_top.MEM[30][22] ),
    .B2(_11030_),
    .X(_07324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11975_ (.A1_N(_10907_),
    .A2_N(_11028_),
    .B1(\design_top.MEM[30][21] ),
    .B2(_11030_),
    .X(_07323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11976_ (.A1_N(_10910_),
    .A2_N(_11028_),
    .B1(\design_top.MEM[30][20] ),
    .B2(_11030_),
    .X(_07322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11977_ (.A1_N(_10913_),
    .A2_N(_11028_),
    .B1(\design_top.MEM[30][19] ),
    .B2(_11030_),
    .X(_07321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11978_ (.A1_N(_10916_),
    .A2_N(_11027_),
    .B1(\design_top.MEM[30][18] ),
    .B2(_11029_),
    .X(_07320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11979_ (.A1_N(_10919_),
    .A2_N(_11027_),
    .B1(\design_top.MEM[30][17] ),
    .B2(_11029_),
    .X(_07319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11980_ (.A1_N(_10922_),
    .A2_N(_11027_),
    .B1(\design_top.MEM[30][16] ),
    .B2(_11029_),
    .X(_07318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11981_ (.A(_10925_),
    .X(_11031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11982_ (.A(_11031_),
    .X(_11032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11983_ (.A(_11032_),
    .B(_11020_),
    .X(_11033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11984_ (.A(_11033_),
    .X(_11034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11985_ (.A1(_10967_),
    .A2(_11011_),
    .B1(_11033_),
    .X(_11035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11986_ (.A(_11035_),
    .X(_11036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11987_ (.A1_N(_10924_),
    .A2_N(_11034_),
    .B1(\design_top.MEM[30][31] ),
    .B2(_11036_),
    .X(_07317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11988_ (.A1_N(_10934_),
    .A2_N(_11034_),
    .B1(\design_top.MEM[30][30] ),
    .B2(_11036_),
    .X(_07316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11989_ (.A1_N(_10937_),
    .A2_N(_11034_),
    .B1(\design_top.MEM[30][29] ),
    .B2(_11036_),
    .X(_07315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11990_ (.A1_N(_10940_),
    .A2_N(_11034_),
    .B1(\design_top.MEM[30][28] ),
    .B2(_11036_),
    .X(_07314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11991_ (.A1_N(_10943_),
    .A2_N(_11034_),
    .B1(\design_top.MEM[30][27] ),
    .B2(_11036_),
    .X(_07313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11992_ (.A1_N(_10946_),
    .A2_N(_11033_),
    .B1(\design_top.MEM[30][26] ),
    .B2(_11035_),
    .X(_07312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11993_ (.A1_N(_10949_),
    .A2_N(_11033_),
    .B1(\design_top.MEM[30][25] ),
    .B2(_11035_),
    .X(_07311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _11994_ (.A1_N(_10952_),
    .A2_N(_11033_),
    .B1(\design_top.MEM[30][24] ),
    .B2(_11035_),
    .X(_07310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11995_ (.A(_10767_),
    .X(_11037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11996_ (.A(_11037_),
    .X(_11038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11997_ (.A(_02660_),
    .B(_10978_),
    .X(_11039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11998_ (.A(_11039_),
    .X(_11040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11999_ (.A(_10956_),
    .B(_11040_),
    .X(_11041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12000_ (.A(_11038_),
    .B(_11041_),
    .X(_11042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12001_ (.A(_11042_),
    .X(_11043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12002_ (.A1(_10892_),
    .A2(_10967_),
    .B1(_11042_),
    .X(_11044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12003_ (.A(_11044_),
    .X(_11045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12004_ (.A1_N(_10955_),
    .A2_N(_11043_),
    .B1(\design_top.MEM[31][15] ),
    .B2(_11045_),
    .X(_07309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12005_ (.A(_10587_),
    .X(_11046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12006_ (.A(_11046_),
    .X(_11047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12007_ (.A1_N(_11047_),
    .A2_N(_11043_),
    .B1(\design_top.MEM[31][14] ),
    .B2(_11045_),
    .X(_07308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12008_ (.A(_10802_),
    .X(_11048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12009_ (.A(_11048_),
    .X(_11049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12010_ (.A1_N(_11049_),
    .A2_N(_11043_),
    .B1(\design_top.MEM[31][13] ),
    .B2(_11045_),
    .X(_07307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12011_ (.A(_10805_),
    .X(_11050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12012_ (.A(_11050_),
    .X(_11051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12013_ (.A1_N(_11051_),
    .A2_N(_11043_),
    .B1(\design_top.MEM[31][12] ),
    .B2(_11045_),
    .X(_07306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12014_ (.A(_10808_),
    .X(_11052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12015_ (.A(_11052_),
    .X(_11053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12016_ (.A1_N(_11053_),
    .A2_N(_11043_),
    .B1(\design_top.MEM[31][11] ),
    .B2(_11045_),
    .X(_07305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12017_ (.A(_10811_),
    .X(_11054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12018_ (.A(_11054_),
    .X(_11055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12019_ (.A1_N(_11055_),
    .A2_N(_11042_),
    .B1(\design_top.MEM[31][10] ),
    .B2(_11044_),
    .X(_07304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12020_ (.A(_10814_),
    .X(_11056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12021_ (.A(_11056_),
    .X(_11057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12022_ (.A1_N(_11057_),
    .A2_N(_11042_),
    .B1(\design_top.MEM[31][9] ),
    .B2(_11044_),
    .X(_07303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12023_ (.A(_10817_),
    .X(_11058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12024_ (.A(_11058_),
    .X(_11059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12025_ (.A1_N(_11059_),
    .A2_N(_11042_),
    .B1(\design_top.MEM[31][8] ),
    .B2(_11044_),
    .X(_07302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12026_ (.A(_10874_),
    .X(_11060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12027_ (.A(_11060_),
    .X(_11061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12028_ (.A(_11026_),
    .B(_11041_),
    .X(_11062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12029_ (.A(_11062_),
    .X(_11063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12030_ (.A1(_10892_),
    .A2(_10966_),
    .B1(_11062_),
    .X(_11064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12031_ (.A(_11064_),
    .X(_11065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12032_ (.A1_N(_11061_),
    .A2_N(_11063_),
    .B1(\design_top.MEM[31][23] ),
    .B2(_11065_),
    .X(_07301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12033_ (.A(_10902_),
    .X(_11066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12034_ (.A(_11066_),
    .X(_11067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12035_ (.A1_N(_11067_),
    .A2_N(_11063_),
    .B1(\design_top.MEM[31][22] ),
    .B2(_11065_),
    .X(_07300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12036_ (.A(_10905_),
    .X(_11068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12037_ (.A(_11068_),
    .X(_11069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12038_ (.A1_N(_11069_),
    .A2_N(_11063_),
    .B1(\design_top.MEM[31][21] ),
    .B2(_11065_),
    .X(_07299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12039_ (.A(_10908_),
    .X(_11070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12040_ (.A(_11070_),
    .X(_11071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12041_ (.A1_N(_11071_),
    .A2_N(_11063_),
    .B1(\design_top.MEM[31][20] ),
    .B2(_11065_),
    .X(_07298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12042_ (.A(_10911_),
    .X(_11072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12043_ (.A(_11072_),
    .X(_11073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12044_ (.A1_N(_11073_),
    .A2_N(_11063_),
    .B1(\design_top.MEM[31][19] ),
    .B2(_11065_),
    .X(_07297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12045_ (.A(_10914_),
    .X(_11074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12046_ (.A(_11074_),
    .X(_11075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12047_ (.A1_N(_11075_),
    .A2_N(_11062_),
    .B1(\design_top.MEM[31][18] ),
    .B2(_11064_),
    .X(_07296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12048_ (.A(_10917_),
    .X(_11076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12049_ (.A(_11076_),
    .X(_11077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12050_ (.A1_N(_11077_),
    .A2_N(_11062_),
    .B1(\design_top.MEM[31][17] ),
    .B2(_11064_),
    .X(_07295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12051_ (.A(_10920_),
    .X(_11078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12052_ (.A(_11078_),
    .X(_11079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12053_ (.A1_N(_11079_),
    .A2_N(_11062_),
    .B1(\design_top.MEM[31][16] ),
    .B2(_11064_),
    .X(_07294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12054_ (.A(_10820_),
    .X(_11080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12055_ (.A(_11080_),
    .X(_11081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12056_ (.A(_11032_),
    .B(_11041_),
    .X(_11082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12057_ (.A(_11082_),
    .X(_11083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12058_ (.A1(_10892_),
    .A2(_10966_),
    .B1(_11082_),
    .X(_11084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12059_ (.A(_11084_),
    .X(_11085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12060_ (.A1_N(_11081_),
    .A2_N(_11083_),
    .B1(\design_top.MEM[31][31] ),
    .B2(_11085_),
    .X(_07293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12061_ (.A(_10932_),
    .X(_11086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12062_ (.A(_11086_),
    .X(_11087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12063_ (.A1_N(_11087_),
    .A2_N(_11083_),
    .B1(\design_top.MEM[31][30] ),
    .B2(_11085_),
    .X(_07292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12064_ (.A(_10935_),
    .X(_11088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12065_ (.A(_11088_),
    .X(_11089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12066_ (.A1_N(_11089_),
    .A2_N(_11083_),
    .B1(\design_top.MEM[31][29] ),
    .B2(_11085_),
    .X(_07291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12067_ (.A(_10938_),
    .X(_11090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12068_ (.A(_11090_),
    .X(_11091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12069_ (.A1_N(_11091_),
    .A2_N(_11083_),
    .B1(\design_top.MEM[31][28] ),
    .B2(_11085_),
    .X(_07290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12070_ (.A(_10941_),
    .X(_11092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12071_ (.A(_11092_),
    .X(_11093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12072_ (.A1_N(_11093_),
    .A2_N(_11083_),
    .B1(\design_top.MEM[31][27] ),
    .B2(_11085_),
    .X(_07289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12073_ (.A(_10944_),
    .X(_11094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12074_ (.A(_11094_),
    .X(_11095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12075_ (.A1_N(_11095_),
    .A2_N(_11082_),
    .B1(\design_top.MEM[31][26] ),
    .B2(_11084_),
    .X(_07288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12076_ (.A(_10947_),
    .X(_11096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12077_ (.A(_11096_),
    .X(_11097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12078_ (.A1_N(_11097_),
    .A2_N(_11082_),
    .B1(\design_top.MEM[31][25] ),
    .B2(_11084_),
    .X(_07287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12079_ (.A(_10950_),
    .X(_11098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12080_ (.A(_11098_),
    .X(_11099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12081_ (.A1_N(_11099_),
    .A2_N(_11082_),
    .B1(\design_top.MEM[31][24] ),
    .B2(_11084_),
    .X(_07286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12082_ (.A(_10953_),
    .X(_11100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12083_ (.A(_11100_),
    .X(_11101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12084_ (.A(_10776_),
    .X(_11102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12085_ (.A(_02862_),
    .B(_03216_),
    .X(_11103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12086_ (.A(_03199_),
    .B(_11103_),
    .X(_11104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12087_ (.A(_11104_),
    .X(_11105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12088_ (.A(_11102_),
    .B(_11105_),
    .X(_11106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12089_ (.A(_11038_),
    .B(_11106_),
    .X(_11107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12090_ (.A(_11107_),
    .X(_11108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12091_ (.A(wbs_adr_i[3]),
    .Y(_11109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12092_ (.A(_11109_),
    .X(_11110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _12093_ (.A(_11110_),
    .B(_10788_),
    .C(_10789_),
    .D(_10790_),
    .X(_11111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12094_ (.A(_11111_),
    .X(_11112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12095_ (.A(_11112_),
    .X(_11113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12096_ (.A1(_10962_),
    .A2(_11113_),
    .B1(_11107_),
    .X(_11114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12097_ (.A(_11114_),
    .X(_11115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12098_ (.A1_N(_11101_),
    .A2_N(_11108_),
    .B1(\design_top.MEM[32][15] ),
    .B2(_11115_),
    .X(_07285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12099_ (.A1_N(_11047_),
    .A2_N(_11108_),
    .B1(\design_top.MEM[32][14] ),
    .B2(_11115_),
    .X(_07284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12100_ (.A1_N(_11049_),
    .A2_N(_11108_),
    .B1(\design_top.MEM[32][13] ),
    .B2(_11115_),
    .X(_07283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12101_ (.A1_N(_11051_),
    .A2_N(_11108_),
    .B1(\design_top.MEM[32][12] ),
    .B2(_11115_),
    .X(_07282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12102_ (.A1_N(_11053_),
    .A2_N(_11108_),
    .B1(\design_top.MEM[32][11] ),
    .B2(_11115_),
    .X(_07281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12103_ (.A1_N(_11055_),
    .A2_N(_11107_),
    .B1(\design_top.MEM[32][10] ),
    .B2(_11114_),
    .X(_07280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12104_ (.A1_N(_11057_),
    .A2_N(_11107_),
    .B1(\design_top.MEM[32][9] ),
    .B2(_11114_),
    .X(_07279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12105_ (.A1_N(_11059_),
    .A2_N(_11107_),
    .B1(\design_top.MEM[32][8] ),
    .B2(_11114_),
    .X(_07278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12106_ (.A(_11026_),
    .B(_11106_),
    .X(_11116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12107_ (.A(_11116_),
    .X(_11117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12108_ (.A1(_10962_),
    .A2(_11113_),
    .B1(_11116_),
    .X(_11118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12109_ (.A(_11118_),
    .X(_11119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12110_ (.A1_N(_11061_),
    .A2_N(_11117_),
    .B1(\design_top.MEM[32][23] ),
    .B2(_11119_),
    .X(_07277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12111_ (.A1_N(_11067_),
    .A2_N(_11117_),
    .B1(\design_top.MEM[32][22] ),
    .B2(_11119_),
    .X(_07276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12112_ (.A1_N(_11069_),
    .A2_N(_11117_),
    .B1(\design_top.MEM[32][21] ),
    .B2(_11119_),
    .X(_07275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12113_ (.A1_N(_11071_),
    .A2_N(_11117_),
    .B1(\design_top.MEM[32][20] ),
    .B2(_11119_),
    .X(_07274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12114_ (.A1_N(_11073_),
    .A2_N(_11117_),
    .B1(\design_top.MEM[32][19] ),
    .B2(_11119_),
    .X(_07273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12115_ (.A1_N(_11075_),
    .A2_N(_11116_),
    .B1(\design_top.MEM[32][18] ),
    .B2(_11118_),
    .X(_07272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12116_ (.A1_N(_11077_),
    .A2_N(_11116_),
    .B1(\design_top.MEM[32][17] ),
    .B2(_11118_),
    .X(_07271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12117_ (.A1_N(_11079_),
    .A2_N(_11116_),
    .B1(\design_top.MEM[32][16] ),
    .B2(_11118_),
    .X(_07270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12118_ (.A(_10784_),
    .B(_10879_),
    .X(_11120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12119_ (.A(_11120_),
    .X(_11121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12120_ (.A1(_10793_),
    .A2(_10799_),
    .B1(_11120_),
    .X(_11122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12121_ (.A(_11122_),
    .X(_11123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12122_ (.A1_N(_11061_),
    .A2_N(_11121_),
    .B1(\design_top.MEM[0][23] ),
    .B2(_11123_),
    .X(_07269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12123_ (.A1_N(_11067_),
    .A2_N(_11121_),
    .B1(\design_top.MEM[0][22] ),
    .B2(_11123_),
    .X(_07268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12124_ (.A1_N(_11069_),
    .A2_N(_11121_),
    .B1(\design_top.MEM[0][21] ),
    .B2(_11123_),
    .X(_07267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12125_ (.A1_N(_11071_),
    .A2_N(_11121_),
    .B1(\design_top.MEM[0][20] ),
    .B2(_11123_),
    .X(_07266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12126_ (.A1_N(_11073_),
    .A2_N(_11121_),
    .B1(\design_top.MEM[0][19] ),
    .B2(_11123_),
    .X(_07265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12127_ (.A1_N(_11075_),
    .A2_N(_11120_),
    .B1(\design_top.MEM[0][18] ),
    .B2(_11122_),
    .X(_07264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12128_ (.A1_N(_11077_),
    .A2_N(_11120_),
    .B1(\design_top.MEM[0][17] ),
    .B2(_11122_),
    .X(_07263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12129_ (.A1_N(_11079_),
    .A2_N(_11120_),
    .B1(\design_top.MEM[0][16] ),
    .B2(_11122_),
    .X(_07262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12130_ (.A(_10784_),
    .B(_10927_),
    .X(_11124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12131_ (.A(_11124_),
    .X(_11125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12132_ (.A(_10792_),
    .X(_11126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12133_ (.A1(_11126_),
    .A2(_10799_),
    .B1(_11124_),
    .X(_11127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12134_ (.A(_11127_),
    .X(_11128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12135_ (.A1_N(_11081_),
    .A2_N(_11125_),
    .B1(\design_top.MEM[0][31] ),
    .B2(_11128_),
    .X(_07261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12136_ (.A1_N(_11087_),
    .A2_N(_11125_),
    .B1(\design_top.MEM[0][30] ),
    .B2(_11128_),
    .X(_07260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12137_ (.A1_N(_11089_),
    .A2_N(_11125_),
    .B1(\design_top.MEM[0][29] ),
    .B2(_11128_),
    .X(_07259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12138_ (.A1_N(_11091_),
    .A2_N(_11125_),
    .B1(\design_top.MEM[0][28] ),
    .B2(_11128_),
    .X(_07258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12139_ (.A1_N(_11093_),
    .A2_N(_11125_),
    .B1(\design_top.MEM[0][27] ),
    .B2(_11128_),
    .X(_07257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12140_ (.A1_N(_11095_),
    .A2_N(_11124_),
    .B1(\design_top.MEM[0][26] ),
    .B2(_11127_),
    .X(_07256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12141_ (.A1_N(_11097_),
    .A2_N(_11124_),
    .B1(\design_top.MEM[0][25] ),
    .B2(_11127_),
    .X(_07255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12142_ (.A1_N(_11099_),
    .A2_N(_11124_),
    .B1(\design_top.MEM[0][24] ),
    .B2(_11127_),
    .X(_07254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12143_ (.A(_02860_),
    .B(_10781_),
    .X(_11129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12144_ (.A(_11129_),
    .X(_11130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12145_ (.A(_11000_),
    .B(_11130_),
    .X(_11131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12146_ (.A(_11038_),
    .B(_11131_),
    .X(_11132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12147_ (.A(_11132_),
    .X(_11133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12148_ (.A(_11004_),
    .X(_11134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12149_ (.A(_11134_),
    .X(_11135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12150_ (.A(_11135_),
    .X(_11136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _12151_ (.A(_10787_),
    .B(_10788_),
    .C(_10896_),
    .D(_10790_),
    .X(_11137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12152_ (.A(_11137_),
    .X(_11138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12153_ (.A(_11138_),
    .X(_11139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12154_ (.A1(_11136_),
    .A2(_11139_),
    .B1(_11132_),
    .X(_11140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12155_ (.A(_11140_),
    .X(_11141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12156_ (.A1_N(_11101_),
    .A2_N(_11133_),
    .B1(\design_top.MEM[10][15] ),
    .B2(_11141_),
    .X(_07253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12157_ (.A1_N(_11047_),
    .A2_N(_11133_),
    .B1(\design_top.MEM[10][14] ),
    .B2(_11141_),
    .X(_07252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12158_ (.A1_N(_11049_),
    .A2_N(_11133_),
    .B1(\design_top.MEM[10][13] ),
    .B2(_11141_),
    .X(_07251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12159_ (.A1_N(_11051_),
    .A2_N(_11133_),
    .B1(\design_top.MEM[10][12] ),
    .B2(_11141_),
    .X(_07250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12160_ (.A1_N(_11053_),
    .A2_N(_11133_),
    .B1(\design_top.MEM[10][11] ),
    .B2(_11141_),
    .X(_07249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12161_ (.A1_N(_11055_),
    .A2_N(_11132_),
    .B1(\design_top.MEM[10][10] ),
    .B2(_11140_),
    .X(_07248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12162_ (.A1_N(_11057_),
    .A2_N(_11132_),
    .B1(\design_top.MEM[10][9] ),
    .B2(_11140_),
    .X(_07247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12163_ (.A1_N(_11059_),
    .A2_N(_11132_),
    .B1(\design_top.MEM[10][8] ),
    .B2(_11140_),
    .X(_07246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12164_ (.A(_11026_),
    .B(_11131_),
    .X(_11142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12165_ (.A(_11142_),
    .X(_11143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12166_ (.A1(_11136_),
    .A2(_11139_),
    .B1(_11142_),
    .X(_11144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12167_ (.A(_11144_),
    .X(_11145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12168_ (.A1_N(_11061_),
    .A2_N(_11143_),
    .B1(\design_top.MEM[10][23] ),
    .B2(_11145_),
    .X(_07245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12169_ (.A1_N(_11067_),
    .A2_N(_11143_),
    .B1(\design_top.MEM[10][22] ),
    .B2(_11145_),
    .X(_07244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12170_ (.A1_N(_11069_),
    .A2_N(_11143_),
    .B1(\design_top.MEM[10][21] ),
    .B2(_11145_),
    .X(_07243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12171_ (.A1_N(_11071_),
    .A2_N(_11143_),
    .B1(\design_top.MEM[10][20] ),
    .B2(_11145_),
    .X(_07242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12172_ (.A1_N(_11073_),
    .A2_N(_11143_),
    .B1(\design_top.MEM[10][19] ),
    .B2(_11145_),
    .X(_07241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12173_ (.A1_N(_11075_),
    .A2_N(_11142_),
    .B1(\design_top.MEM[10][18] ),
    .B2(_11144_),
    .X(_07240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12174_ (.A1_N(_11077_),
    .A2_N(_11142_),
    .B1(\design_top.MEM[10][17] ),
    .B2(_11144_),
    .X(_07239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12175_ (.A1_N(_11079_),
    .A2_N(_11142_),
    .B1(\design_top.MEM[10][16] ),
    .B2(_11144_),
    .X(_07238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12176_ (.A(_11032_),
    .B(_11131_),
    .X(_11146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12177_ (.A(_11146_),
    .X(_11147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12178_ (.A1(_11136_),
    .A2(_11139_),
    .B1(_11146_),
    .X(_11148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12179_ (.A(_11148_),
    .X(_11149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12180_ (.A1_N(_11081_),
    .A2_N(_11147_),
    .B1(\design_top.MEM[10][31] ),
    .B2(_11149_),
    .X(_07237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12181_ (.A1_N(_11087_),
    .A2_N(_11147_),
    .B1(\design_top.MEM[10][30] ),
    .B2(_11149_),
    .X(_07236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12182_ (.A1_N(_11089_),
    .A2_N(_11147_),
    .B1(\design_top.MEM[10][29] ),
    .B2(_11149_),
    .X(_07235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12183_ (.A1_N(_11091_),
    .A2_N(_11147_),
    .B1(\design_top.MEM[10][28] ),
    .B2(_11149_),
    .X(_07234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12184_ (.A1_N(_11093_),
    .A2_N(_11147_),
    .B1(\design_top.MEM[10][27] ),
    .B2(_11149_),
    .X(_07233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12185_ (.A1_N(_11095_),
    .A2_N(_11146_),
    .B1(\design_top.MEM[10][26] ),
    .B2(_11148_),
    .X(_07232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12186_ (.A1_N(_11097_),
    .A2_N(_11146_),
    .B1(\design_top.MEM[10][25] ),
    .B2(_11148_),
    .X(_07231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12187_ (.A1_N(_11099_),
    .A2_N(_11146_),
    .B1(\design_top.MEM[10][24] ),
    .B2(_11148_),
    .X(_07230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12188_ (.A(_10885_),
    .B(_11130_),
    .X(_11150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12189_ (.A(_11038_),
    .B(_11150_),
    .X(_11151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12190_ (.A(_11151_),
    .X(_11152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12191_ (.A(_10891_),
    .X(_11153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12192_ (.A1(_11153_),
    .A2(_11139_),
    .B1(_11151_),
    .X(_11154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12193_ (.A(_11154_),
    .X(_11155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12194_ (.A1_N(_11101_),
    .A2_N(_11152_),
    .B1(\design_top.MEM[11][15] ),
    .B2(_11155_),
    .X(_07229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12195_ (.A1_N(_11047_),
    .A2_N(_11152_),
    .B1(\design_top.MEM[11][14] ),
    .B2(_11155_),
    .X(_07228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12196_ (.A1_N(_11049_),
    .A2_N(_11152_),
    .B1(\design_top.MEM[11][13] ),
    .B2(_11155_),
    .X(_07227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12197_ (.A1_N(_11051_),
    .A2_N(_11152_),
    .B1(\design_top.MEM[11][12] ),
    .B2(_11155_),
    .X(_07226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12198_ (.A1_N(_11053_),
    .A2_N(_11152_),
    .B1(\design_top.MEM[11][11] ),
    .B2(_11155_),
    .X(_07225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12199_ (.A1_N(_11055_),
    .A2_N(_11151_),
    .B1(\design_top.MEM[11][10] ),
    .B2(_11154_),
    .X(_07224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12200_ (.A1_N(_11057_),
    .A2_N(_11151_),
    .B1(\design_top.MEM[11][9] ),
    .B2(_11154_),
    .X(_07223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12201_ (.A1_N(_11059_),
    .A2_N(_11151_),
    .B1(\design_top.MEM[11][8] ),
    .B2(_11154_),
    .X(_07222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12202_ (.A(_11026_),
    .B(_11150_),
    .X(_11156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12203_ (.A(_11156_),
    .X(_11157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12204_ (.A1(_11153_),
    .A2(_11139_),
    .B1(_11156_),
    .X(_11158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12205_ (.A(_11158_),
    .X(_11159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12206_ (.A1_N(_11061_),
    .A2_N(_11157_),
    .B1(\design_top.MEM[11][23] ),
    .B2(_11159_),
    .X(_07221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12207_ (.A1_N(_11067_),
    .A2_N(_11157_),
    .B1(\design_top.MEM[11][22] ),
    .B2(_11159_),
    .X(_07220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12208_ (.A1_N(_11069_),
    .A2_N(_11157_),
    .B1(\design_top.MEM[11][21] ),
    .B2(_11159_),
    .X(_07219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12209_ (.A1_N(_11071_),
    .A2_N(_11157_),
    .B1(\design_top.MEM[11][20] ),
    .B2(_11159_),
    .X(_07218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12210_ (.A1_N(_11073_),
    .A2_N(_11157_),
    .B1(\design_top.MEM[11][19] ),
    .B2(_11159_),
    .X(_07217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12211_ (.A1_N(_11075_),
    .A2_N(_11156_),
    .B1(\design_top.MEM[11][18] ),
    .B2(_11158_),
    .X(_07216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12212_ (.A1_N(_11077_),
    .A2_N(_11156_),
    .B1(\design_top.MEM[11][17] ),
    .B2(_11158_),
    .X(_07215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12213_ (.A1_N(_11079_),
    .A2_N(_11156_),
    .B1(\design_top.MEM[11][16] ),
    .B2(_11158_),
    .X(_07214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12214_ (.A(_11032_),
    .B(_11150_),
    .X(_11160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12215_ (.A(_11160_),
    .X(_11161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12216_ (.A(_11138_),
    .X(_11162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12217_ (.A1(_11153_),
    .A2(_11162_),
    .B1(_11160_),
    .X(_11163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12218_ (.A(_11163_),
    .X(_11164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12219_ (.A1_N(_11081_),
    .A2_N(_11161_),
    .B1(\design_top.MEM[11][31] ),
    .B2(_11164_),
    .X(_07213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12220_ (.A1_N(_11087_),
    .A2_N(_11161_),
    .B1(\design_top.MEM[11][30] ),
    .B2(_11164_),
    .X(_07212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12221_ (.A1_N(_11089_),
    .A2_N(_11161_),
    .B1(\design_top.MEM[11][29] ),
    .B2(_11164_),
    .X(_07211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12222_ (.A1_N(_11091_),
    .A2_N(_11161_),
    .B1(\design_top.MEM[11][28] ),
    .B2(_11164_),
    .X(_07210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12223_ (.A1_N(_11093_),
    .A2_N(_11161_),
    .B1(\design_top.MEM[11][27] ),
    .B2(_11164_),
    .X(_07209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12224_ (.A1_N(_11095_),
    .A2_N(_11160_),
    .B1(\design_top.MEM[11][26] ),
    .B2(_11163_),
    .X(_07208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12225_ (.A1_N(_11097_),
    .A2_N(_11160_),
    .B1(\design_top.MEM[11][25] ),
    .B2(_11163_),
    .X(_07207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12226_ (.A1_N(_11099_),
    .A2_N(_11160_),
    .B1(\design_top.MEM[11][24] ),
    .B2(_11163_),
    .X(_07206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12227_ (.A(_10958_),
    .B(_11130_),
    .X(_11165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12228_ (.A(_11038_),
    .B(_11165_),
    .X(_11166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12229_ (.A(_11166_),
    .X(_11167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12230_ (.A(_10799_),
    .X(_11168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _12231_ (.A(_10787_),
    .B(_10788_),
    .C(_10896_),
    .D(_10964_),
    .X(_11169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12232_ (.A(_11169_),
    .X(_11170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12233_ (.A(_11170_),
    .X(_11171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12234_ (.A1(_11168_),
    .A2(_11171_),
    .B1(_11166_),
    .X(_11172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12235_ (.A(_11172_),
    .X(_11173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12236_ (.A1_N(_11101_),
    .A2_N(_11167_),
    .B1(\design_top.MEM[12][15] ),
    .B2(_11173_),
    .X(_07205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12237_ (.A1_N(_11047_),
    .A2_N(_11167_),
    .B1(\design_top.MEM[12][14] ),
    .B2(_11173_),
    .X(_07204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12238_ (.A1_N(_11049_),
    .A2_N(_11167_),
    .B1(\design_top.MEM[12][13] ),
    .B2(_11173_),
    .X(_07203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12239_ (.A1_N(_11051_),
    .A2_N(_11167_),
    .B1(\design_top.MEM[12][12] ),
    .B2(_11173_),
    .X(_07202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12240_ (.A1_N(_11053_),
    .A2_N(_11167_),
    .B1(\design_top.MEM[12][11] ),
    .B2(_11173_),
    .X(_07201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12241_ (.A1_N(_11055_),
    .A2_N(_11166_),
    .B1(\design_top.MEM[12][10] ),
    .B2(_11172_),
    .X(_07200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12242_ (.A1_N(_11057_),
    .A2_N(_11166_),
    .B1(\design_top.MEM[12][9] ),
    .B2(_11172_),
    .X(_07199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12243_ (.A1_N(_11059_),
    .A2_N(_11166_),
    .B1(\design_top.MEM[12][8] ),
    .B2(_11172_),
    .X(_07198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12244_ (.A(_11060_),
    .X(_11174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12245_ (.A(_11025_),
    .X(_11175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12246_ (.A(_11175_),
    .B(_11165_),
    .X(_11176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12247_ (.A(_11176_),
    .X(_11177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12248_ (.A1(_11168_),
    .A2(_11171_),
    .B1(_11176_),
    .X(_11178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12249_ (.A(_11178_),
    .X(_11179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12250_ (.A1_N(_11174_),
    .A2_N(_11177_),
    .B1(\design_top.MEM[12][23] ),
    .B2(_11179_),
    .X(_07197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12251_ (.A(_11066_),
    .X(_11180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12252_ (.A1_N(_11180_),
    .A2_N(_11177_),
    .B1(\design_top.MEM[12][22] ),
    .B2(_11179_),
    .X(_07196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12253_ (.A(_11068_),
    .X(_11181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12254_ (.A1_N(_11181_),
    .A2_N(_11177_),
    .B1(\design_top.MEM[12][21] ),
    .B2(_11179_),
    .X(_07195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12255_ (.A(_11070_),
    .X(_11182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12256_ (.A1_N(_11182_),
    .A2_N(_11177_),
    .B1(\design_top.MEM[12][20] ),
    .B2(_11179_),
    .X(_07194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12257_ (.A(_11072_),
    .X(_11183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12258_ (.A1_N(_11183_),
    .A2_N(_11177_),
    .B1(\design_top.MEM[12][19] ),
    .B2(_11179_),
    .X(_07193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12259_ (.A(_11074_),
    .X(_11184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12260_ (.A1_N(_11184_),
    .A2_N(_11176_),
    .B1(\design_top.MEM[12][18] ),
    .B2(_11178_),
    .X(_07192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12261_ (.A(_11076_),
    .X(_11185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12262_ (.A1_N(_11185_),
    .A2_N(_11176_),
    .B1(\design_top.MEM[12][17] ),
    .B2(_11178_),
    .X(_07191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12263_ (.A(_11078_),
    .X(_11186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12264_ (.A1_N(_11186_),
    .A2_N(_11176_),
    .B1(\design_top.MEM[12][16] ),
    .B2(_11178_),
    .X(_07190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12265_ (.A(_11032_),
    .B(_11165_),
    .X(_11187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12266_ (.A(_11187_),
    .X(_11188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12267_ (.A1(_11168_),
    .A2(_11171_),
    .B1(_11187_),
    .X(_11189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12268_ (.A(_11189_),
    .X(_11190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12269_ (.A1_N(_11081_),
    .A2_N(_11188_),
    .B1(\design_top.MEM[12][31] ),
    .B2(_11190_),
    .X(_07189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12270_ (.A1_N(_11087_),
    .A2_N(_11188_),
    .B1(\design_top.MEM[12][30] ),
    .B2(_11190_),
    .X(_07188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12271_ (.A1_N(_11089_),
    .A2_N(_11188_),
    .B1(\design_top.MEM[12][29] ),
    .B2(_11190_),
    .X(_07187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12272_ (.A1_N(_11091_),
    .A2_N(_11188_),
    .B1(\design_top.MEM[12][28] ),
    .B2(_11190_),
    .X(_07186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12273_ (.A1_N(_11093_),
    .A2_N(_11188_),
    .B1(\design_top.MEM[12][27] ),
    .B2(_11190_),
    .X(_07185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12274_ (.A1_N(_11095_),
    .A2_N(_11187_),
    .B1(\design_top.MEM[12][26] ),
    .B2(_11189_),
    .X(_07184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12275_ (.A1_N(_11097_),
    .A2_N(_11187_),
    .B1(\design_top.MEM[12][25] ),
    .B2(_11189_),
    .X(_07183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12276_ (.A1_N(_11099_),
    .A2_N(_11187_),
    .B1(\design_top.MEM[12][24] ),
    .B2(_11189_),
    .X(_07182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12277_ (.A(_11037_),
    .X(_11191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12278_ (.A(_10980_),
    .B(_11130_),
    .X(_11192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12279_ (.A(_11191_),
    .B(_11192_),
    .X(_11193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12280_ (.A(_11193_),
    .X(_11194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12281_ (.A(_10985_),
    .X(_11195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12282_ (.A(_11195_),
    .X(_11196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12283_ (.A(_11196_),
    .X(_11197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12284_ (.A1(_11197_),
    .A2(_11171_),
    .B1(_11193_),
    .X(_11198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12285_ (.A(_11198_),
    .X(_11199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12286_ (.A1_N(_11101_),
    .A2_N(_11194_),
    .B1(\design_top.MEM[13][15] ),
    .B2(_11199_),
    .X(_07181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12287_ (.A(_11046_),
    .X(_11200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12288_ (.A1_N(_11200_),
    .A2_N(_11194_),
    .B1(\design_top.MEM[13][14] ),
    .B2(_11199_),
    .X(_07180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12289_ (.A(_11048_),
    .X(_11201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12290_ (.A1_N(_11201_),
    .A2_N(_11194_),
    .B1(\design_top.MEM[13][13] ),
    .B2(_11199_),
    .X(_07179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12291_ (.A(_11050_),
    .X(_11202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12292_ (.A1_N(_11202_),
    .A2_N(_11194_),
    .B1(\design_top.MEM[13][12] ),
    .B2(_11199_),
    .X(_07178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12293_ (.A(_11052_),
    .X(_11203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12294_ (.A1_N(_11203_),
    .A2_N(_11194_),
    .B1(\design_top.MEM[13][11] ),
    .B2(_11199_),
    .X(_07177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12295_ (.A(_11054_),
    .X(_11204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12296_ (.A1_N(_11204_),
    .A2_N(_11193_),
    .B1(\design_top.MEM[13][10] ),
    .B2(_11198_),
    .X(_07176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12297_ (.A(_11056_),
    .X(_11205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12298_ (.A1_N(_11205_),
    .A2_N(_11193_),
    .B1(\design_top.MEM[13][9] ),
    .B2(_11198_),
    .X(_07175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12299_ (.A(_11058_),
    .X(_11206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12300_ (.A1_N(_11206_),
    .A2_N(_11193_),
    .B1(\design_top.MEM[13][8] ),
    .B2(_11198_),
    .X(_07174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12301_ (.A(_11175_),
    .B(_11192_),
    .X(_11207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12302_ (.A(_11207_),
    .X(_11208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12303_ (.A1(_11197_),
    .A2(_11171_),
    .B1(_11207_),
    .X(_11209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12304_ (.A(_11209_),
    .X(_11210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12305_ (.A1_N(_11174_),
    .A2_N(_11208_),
    .B1(\design_top.MEM[13][23] ),
    .B2(_11210_),
    .X(_07173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12306_ (.A1_N(_11180_),
    .A2_N(_11208_),
    .B1(\design_top.MEM[13][22] ),
    .B2(_11210_),
    .X(_07172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12307_ (.A1_N(_11181_),
    .A2_N(_11208_),
    .B1(\design_top.MEM[13][21] ),
    .B2(_11210_),
    .X(_07171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12308_ (.A1_N(_11182_),
    .A2_N(_11208_),
    .B1(\design_top.MEM[13][20] ),
    .B2(_11210_),
    .X(_07170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12309_ (.A1_N(_11183_),
    .A2_N(_11208_),
    .B1(\design_top.MEM[13][19] ),
    .B2(_11210_),
    .X(_07169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12310_ (.A1_N(_11184_),
    .A2_N(_11207_),
    .B1(\design_top.MEM[13][18] ),
    .B2(_11209_),
    .X(_07168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12311_ (.A1_N(_11185_),
    .A2_N(_11207_),
    .B1(\design_top.MEM[13][17] ),
    .B2(_11209_),
    .X(_07167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12312_ (.A1_N(_11186_),
    .A2_N(_11207_),
    .B1(\design_top.MEM[13][16] ),
    .B2(_11209_),
    .X(_07166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12313_ (.A(_11080_),
    .X(_11211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12314_ (.A(_11031_),
    .X(_11212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12315_ (.A(_11212_),
    .B(_11192_),
    .X(_11213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12316_ (.A(_11213_),
    .X(_11214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12317_ (.A(_11170_),
    .X(_11215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12318_ (.A1(_11197_),
    .A2(_11215_),
    .B1(_11213_),
    .X(_11216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12319_ (.A(_11216_),
    .X(_11217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12320_ (.A1_N(_11211_),
    .A2_N(_11214_),
    .B1(\design_top.MEM[13][31] ),
    .B2(_11217_),
    .X(_07165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12321_ (.A(_11086_),
    .X(_11218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12322_ (.A1_N(_11218_),
    .A2_N(_11214_),
    .B1(\design_top.MEM[13][30] ),
    .B2(_11217_),
    .X(_07164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12323_ (.A(_11088_),
    .X(_11219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12324_ (.A1_N(_11219_),
    .A2_N(_11214_),
    .B1(\design_top.MEM[13][29] ),
    .B2(_11217_),
    .X(_07163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12325_ (.A(_11090_),
    .X(_11220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12326_ (.A1_N(_11220_),
    .A2_N(_11214_),
    .B1(\design_top.MEM[13][28] ),
    .B2(_11217_),
    .X(_07162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12327_ (.A(_11092_),
    .X(_11221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12328_ (.A1_N(_11221_),
    .A2_N(_11214_),
    .B1(\design_top.MEM[13][27] ),
    .B2(_11217_),
    .X(_07161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12329_ (.A(_11094_),
    .X(_11222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12330_ (.A1_N(_11222_),
    .A2_N(_11213_),
    .B1(\design_top.MEM[13][26] ),
    .B2(_11216_),
    .X(_07160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12331_ (.A(_11096_),
    .X(_11223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12332_ (.A1_N(_11223_),
    .A2_N(_11213_),
    .B1(\design_top.MEM[13][25] ),
    .B2(_11216_),
    .X(_07159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12333_ (.A(_11098_),
    .X(_11224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12334_ (.A1_N(_11224_),
    .A2_N(_11213_),
    .B1(\design_top.MEM[13][24] ),
    .B2(_11216_),
    .X(_07158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12335_ (.A(_11100_),
    .X(_11225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12336_ (.A(_11019_),
    .B(_11130_),
    .X(_11226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12337_ (.A(_11191_),
    .B(_11226_),
    .X(_11227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12338_ (.A(_11227_),
    .X(_11228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12339_ (.A1(_11136_),
    .A2(_11215_),
    .B1(_11227_),
    .X(_11229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12340_ (.A(_11229_),
    .X(_11230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12341_ (.A1_N(_11225_),
    .A2_N(_11228_),
    .B1(\design_top.MEM[14][15] ),
    .B2(_11230_),
    .X(_07157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12342_ (.A1_N(_11200_),
    .A2_N(_11228_),
    .B1(\design_top.MEM[14][14] ),
    .B2(_11230_),
    .X(_07156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12343_ (.A1_N(_11201_),
    .A2_N(_11228_),
    .B1(\design_top.MEM[14][13] ),
    .B2(_11230_),
    .X(_07155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12344_ (.A1_N(_11202_),
    .A2_N(_11228_),
    .B1(\design_top.MEM[14][12] ),
    .B2(_11230_),
    .X(_07154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12345_ (.A1_N(_11203_),
    .A2_N(_11228_),
    .B1(\design_top.MEM[14][11] ),
    .B2(_11230_),
    .X(_07153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12346_ (.A1_N(_11204_),
    .A2_N(_11227_),
    .B1(\design_top.MEM[14][10] ),
    .B2(_11229_),
    .X(_07152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12347_ (.A1_N(_11205_),
    .A2_N(_11227_),
    .B1(\design_top.MEM[14][9] ),
    .B2(_11229_),
    .X(_07151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12348_ (.A1_N(_11206_),
    .A2_N(_11227_),
    .B1(\design_top.MEM[14][8] ),
    .B2(_11229_),
    .X(_07150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12349_ (.A(_11175_),
    .B(_11226_),
    .X(_11231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12350_ (.A(_11231_),
    .X(_11232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12351_ (.A1(_11136_),
    .A2(_11215_),
    .B1(_11231_),
    .X(_11233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12352_ (.A(_11233_),
    .X(_11234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12353_ (.A1_N(_11174_),
    .A2_N(_11232_),
    .B1(\design_top.MEM[14][23] ),
    .B2(_11234_),
    .X(_07149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12354_ (.A1_N(_11180_),
    .A2_N(_11232_),
    .B1(\design_top.MEM[14][22] ),
    .B2(_11234_),
    .X(_07148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12355_ (.A1_N(_11181_),
    .A2_N(_11232_),
    .B1(\design_top.MEM[14][21] ),
    .B2(_11234_),
    .X(_07147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12356_ (.A1_N(_11182_),
    .A2_N(_11232_),
    .B1(\design_top.MEM[14][20] ),
    .B2(_11234_),
    .X(_07146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12357_ (.A1_N(_11183_),
    .A2_N(_11232_),
    .B1(\design_top.MEM[14][19] ),
    .B2(_11234_),
    .X(_07145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12358_ (.A1_N(_11184_),
    .A2_N(_11231_),
    .B1(\design_top.MEM[14][18] ),
    .B2(_11233_),
    .X(_07144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12359_ (.A1_N(_11185_),
    .A2_N(_11231_),
    .B1(\design_top.MEM[14][17] ),
    .B2(_11233_),
    .X(_07143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12360_ (.A1_N(_11186_),
    .A2_N(_11231_),
    .B1(\design_top.MEM[14][16] ),
    .B2(_11233_),
    .X(_07142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12361_ (.A(_11212_),
    .B(_11226_),
    .X(_11235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12362_ (.A(_11235_),
    .X(_11236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12363_ (.A(_11135_),
    .X(_11237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12364_ (.A1(_11237_),
    .A2(_11215_),
    .B1(_11235_),
    .X(_11238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12365_ (.A(_11238_),
    .X(_11239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12366_ (.A1_N(_11211_),
    .A2_N(_11236_),
    .B1(\design_top.MEM[14][31] ),
    .B2(_11239_),
    .X(_07141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12367_ (.A1_N(_11218_),
    .A2_N(_11236_),
    .B1(\design_top.MEM[14][30] ),
    .B2(_11239_),
    .X(_07140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12368_ (.A1_N(_11219_),
    .A2_N(_11236_),
    .B1(\design_top.MEM[14][29] ),
    .B2(_11239_),
    .X(_07139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12369_ (.A1_N(_11220_),
    .A2_N(_11236_),
    .B1(\design_top.MEM[14][28] ),
    .B2(_11239_),
    .X(_07138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12370_ (.A1_N(_11221_),
    .A2_N(_11236_),
    .B1(\design_top.MEM[14][27] ),
    .B2(_11239_),
    .X(_07137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12371_ (.A1_N(_11222_),
    .A2_N(_11235_),
    .B1(\design_top.MEM[14][26] ),
    .B2(_11238_),
    .X(_07136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12372_ (.A1_N(_11223_),
    .A2_N(_11235_),
    .B1(\design_top.MEM[14][25] ),
    .B2(_11238_),
    .X(_07135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12373_ (.A1_N(_11224_),
    .A2_N(_11235_),
    .B1(\design_top.MEM[14][24] ),
    .B2(_11238_),
    .X(_07134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12374_ (.A(_11040_),
    .B(_11129_),
    .X(_11240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12375_ (.A(_11191_),
    .B(_11240_),
    .X(_11241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12376_ (.A(_11241_),
    .X(_11242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12377_ (.A1(_11153_),
    .A2(_11215_),
    .B1(_11241_),
    .X(_11243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12378_ (.A(_11243_),
    .X(_11244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12379_ (.A1_N(_11225_),
    .A2_N(_11242_),
    .B1(\design_top.MEM[15][15] ),
    .B2(_11244_),
    .X(_07133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12380_ (.A1_N(_11200_),
    .A2_N(_11242_),
    .B1(\design_top.MEM[15][14] ),
    .B2(_11244_),
    .X(_07132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12381_ (.A1_N(_11201_),
    .A2_N(_11242_),
    .B1(\design_top.MEM[15][13] ),
    .B2(_11244_),
    .X(_07131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12382_ (.A1_N(_11202_),
    .A2_N(_11242_),
    .B1(\design_top.MEM[15][12] ),
    .B2(_11244_),
    .X(_07130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12383_ (.A1_N(_11203_),
    .A2_N(_11242_),
    .B1(\design_top.MEM[15][11] ),
    .B2(_11244_),
    .X(_07129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12384_ (.A1_N(_11204_),
    .A2_N(_11241_),
    .B1(\design_top.MEM[15][10] ),
    .B2(_11243_),
    .X(_07128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12385_ (.A1_N(_11205_),
    .A2_N(_11241_),
    .B1(\design_top.MEM[15][9] ),
    .B2(_11243_),
    .X(_07127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12386_ (.A1_N(_11206_),
    .A2_N(_11241_),
    .B1(\design_top.MEM[15][8] ),
    .B2(_11243_),
    .X(_07126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12387_ (.A(_11175_),
    .B(_11240_),
    .X(_11245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12388_ (.A(_11245_),
    .X(_11246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12389_ (.A1(_11153_),
    .A2(_11170_),
    .B1(_11245_),
    .X(_11247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12390_ (.A(_11247_),
    .X(_11248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12391_ (.A1_N(_11174_),
    .A2_N(_11246_),
    .B1(\design_top.MEM[15][23] ),
    .B2(_11248_),
    .X(_07125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12392_ (.A1_N(_11180_),
    .A2_N(_11246_),
    .B1(\design_top.MEM[15][22] ),
    .B2(_11248_),
    .X(_07124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12393_ (.A1_N(_11181_),
    .A2_N(_11246_),
    .B1(\design_top.MEM[15][21] ),
    .B2(_11248_),
    .X(_07123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12394_ (.A1_N(_11182_),
    .A2_N(_11246_),
    .B1(\design_top.MEM[15][20] ),
    .B2(_11248_),
    .X(_07122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12395_ (.A1_N(_11183_),
    .A2_N(_11246_),
    .B1(\design_top.MEM[15][19] ),
    .B2(_11248_),
    .X(_07121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12396_ (.A1_N(_11184_),
    .A2_N(_11245_),
    .B1(\design_top.MEM[15][18] ),
    .B2(_11247_),
    .X(_07120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12397_ (.A1_N(_11185_),
    .A2_N(_11245_),
    .B1(\design_top.MEM[15][17] ),
    .B2(_11247_),
    .X(_07119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12398_ (.A1_N(_11186_),
    .A2_N(_11245_),
    .B1(\design_top.MEM[15][16] ),
    .B2(_11247_),
    .X(_07118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12399_ (.A(_11212_),
    .B(_11240_),
    .X(_11249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12400_ (.A(_11249_),
    .X(_11250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12401_ (.A(_10890_),
    .X(_11251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12402_ (.A(_11251_),
    .X(_11252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12403_ (.A1(_11252_),
    .A2(_11170_),
    .B1(_11249_),
    .X(_11253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12404_ (.A(_11253_),
    .X(_11254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12405_ (.A1_N(_11211_),
    .A2_N(_11250_),
    .B1(\design_top.MEM[15][31] ),
    .B2(_11254_),
    .X(_07117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12406_ (.A1_N(_11218_),
    .A2_N(_11250_),
    .B1(\design_top.MEM[15][30] ),
    .B2(_11254_),
    .X(_07116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12407_ (.A1_N(_11219_),
    .A2_N(_11250_),
    .B1(\design_top.MEM[15][29] ),
    .B2(_11254_),
    .X(_07115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12408_ (.A1_N(_11220_),
    .A2_N(_11250_),
    .B1(\design_top.MEM[15][28] ),
    .B2(_11254_),
    .X(_07114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12409_ (.A1_N(_11221_),
    .A2_N(_11250_),
    .B1(\design_top.MEM[15][27] ),
    .B2(_11254_),
    .X(_07113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12410_ (.A1_N(_11222_),
    .A2_N(_11249_),
    .B1(\design_top.MEM[15][26] ),
    .B2(_11253_),
    .X(_07112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12411_ (.A1_N(_11223_),
    .A2_N(_11249_),
    .B1(\design_top.MEM[15][25] ),
    .B2(_11253_),
    .X(_07111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12412_ (.A1_N(_11224_),
    .A2_N(_11249_),
    .B1(\design_top.MEM[15][24] ),
    .B2(_11253_),
    .X(_07110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12413_ (.A(_03199_),
    .B(_10880_),
    .X(_11255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12414_ (.A(_11255_),
    .X(_11256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12415_ (.A(_11102_),
    .B(_11256_),
    .X(_11257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12416_ (.A(_11191_),
    .B(_11257_),
    .X(_11258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12417_ (.A(_11258_),
    .X(_11259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _12418_ (.A(wbs_adr_i[3]),
    .B(_10894_),
    .C(_10789_),
    .D(_10790_),
    .X(_11260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12419_ (.A(_11260_),
    .X(_11261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12420_ (.A(_11261_),
    .X(_11262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12421_ (.A1(_11168_),
    .A2(_11262_),
    .B1(_11258_),
    .X(_11263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12422_ (.A(_11263_),
    .X(_11264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12423_ (.A1_N(_11225_),
    .A2_N(_11259_),
    .B1(\design_top.MEM[16][15] ),
    .B2(_11264_),
    .X(_07109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12424_ (.A1_N(_11200_),
    .A2_N(_11259_),
    .B1(\design_top.MEM[16][14] ),
    .B2(_11264_),
    .X(_07108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12425_ (.A1_N(_11201_),
    .A2_N(_11259_),
    .B1(\design_top.MEM[16][13] ),
    .B2(_11264_),
    .X(_07107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12426_ (.A1_N(_11202_),
    .A2_N(_11259_),
    .B1(\design_top.MEM[16][12] ),
    .B2(_11264_),
    .X(_07106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12427_ (.A1_N(_11203_),
    .A2_N(_11259_),
    .B1(\design_top.MEM[16][11] ),
    .B2(_11264_),
    .X(_07105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12428_ (.A1_N(_11204_),
    .A2_N(_11258_),
    .B1(\design_top.MEM[16][10] ),
    .B2(_11263_),
    .X(_07104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12429_ (.A1_N(_11205_),
    .A2_N(_11258_),
    .B1(\design_top.MEM[16][9] ),
    .B2(_11263_),
    .X(_07103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12430_ (.A1_N(_11206_),
    .A2_N(_11258_),
    .B1(\design_top.MEM[16][8] ),
    .B2(_11263_),
    .X(_07102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12431_ (.A(_11175_),
    .B(_11257_),
    .X(_11265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12432_ (.A(_11265_),
    .X(_11266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12433_ (.A1(_11168_),
    .A2(_11262_),
    .B1(_11265_),
    .X(_11267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12434_ (.A(_11267_),
    .X(_11268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12435_ (.A1_N(_11174_),
    .A2_N(_11266_),
    .B1(\design_top.MEM[16][23] ),
    .B2(_11268_),
    .X(_07101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12436_ (.A1_N(_11180_),
    .A2_N(_11266_),
    .B1(\design_top.MEM[16][22] ),
    .B2(_11268_),
    .X(_07100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12437_ (.A1_N(_11181_),
    .A2_N(_11266_),
    .B1(\design_top.MEM[16][21] ),
    .B2(_11268_),
    .X(_07099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12438_ (.A1_N(_11182_),
    .A2_N(_11266_),
    .B1(\design_top.MEM[16][20] ),
    .B2(_11268_),
    .X(_07098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12439_ (.A1_N(_11183_),
    .A2_N(_11266_),
    .B1(\design_top.MEM[16][19] ),
    .B2(_11268_),
    .X(_07097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12440_ (.A1_N(_11184_),
    .A2_N(_11265_),
    .B1(\design_top.MEM[16][18] ),
    .B2(_11267_),
    .X(_07096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12441_ (.A1_N(_11185_),
    .A2_N(_11265_),
    .B1(\design_top.MEM[16][17] ),
    .B2(_11267_),
    .X(_07095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12442_ (.A1_N(_11186_),
    .A2_N(_11265_),
    .B1(\design_top.MEM[16][16] ),
    .B2(_11267_),
    .X(_07094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12443_ (.A(_11212_),
    .B(_11257_),
    .X(_11269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12444_ (.A(_11269_),
    .X(_11270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12445_ (.A(_10798_),
    .X(_11271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12446_ (.A(_11271_),
    .X(_11272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12447_ (.A1(_11272_),
    .A2(_11262_),
    .B1(_11269_),
    .X(_11273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12448_ (.A(_11273_),
    .X(_11274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12449_ (.A1_N(_11211_),
    .A2_N(_11270_),
    .B1(\design_top.MEM[16][31] ),
    .B2(_11274_),
    .X(_07093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12450_ (.A1_N(_11218_),
    .A2_N(_11270_),
    .B1(\design_top.MEM[16][30] ),
    .B2(_11274_),
    .X(_07092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12451_ (.A1_N(_11219_),
    .A2_N(_11270_),
    .B1(\design_top.MEM[16][29] ),
    .B2(_11274_),
    .X(_07091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12452_ (.A1_N(_11220_),
    .A2_N(_11270_),
    .B1(\design_top.MEM[16][28] ),
    .B2(_11274_),
    .X(_07090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12453_ (.A1_N(_11221_),
    .A2_N(_11270_),
    .B1(\design_top.MEM[16][27] ),
    .B2(_11274_),
    .X(_07089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12454_ (.A1_N(_11222_),
    .A2_N(_11269_),
    .B1(\design_top.MEM[16][26] ),
    .B2(_11273_),
    .X(_07088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12455_ (.A1_N(_11223_),
    .A2_N(_11269_),
    .B1(\design_top.MEM[16][25] ),
    .B2(_11273_),
    .X(_07087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12456_ (.A1_N(_11224_),
    .A2_N(_11269_),
    .B1(\design_top.MEM[16][24] ),
    .B2(_11273_),
    .X(_07086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12457_ (.A(_10774_),
    .B(_02651_),
    .X(_11275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12458_ (.A(_11275_),
    .X(_11276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12459_ (.A(_11255_),
    .B(_11276_),
    .X(_11277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12460_ (.A(_11191_),
    .B(_11277_),
    .X(_11278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12461_ (.A(_11278_),
    .X(_11279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12462_ (.A1(_11197_),
    .A2(_11262_),
    .B1(_11278_),
    .X(_11280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12463_ (.A(_11280_),
    .X(_11281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12464_ (.A1_N(_11225_),
    .A2_N(_11279_),
    .B1(\design_top.MEM[17][15] ),
    .B2(_11281_),
    .X(_07085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12465_ (.A1_N(_11200_),
    .A2_N(_11279_),
    .B1(\design_top.MEM[17][14] ),
    .B2(_11281_),
    .X(_07084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12466_ (.A1_N(_11201_),
    .A2_N(_11279_),
    .B1(\design_top.MEM[17][13] ),
    .B2(_11281_),
    .X(_07083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12467_ (.A1_N(_11202_),
    .A2_N(_11279_),
    .B1(\design_top.MEM[17][12] ),
    .B2(_11281_),
    .X(_07082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12468_ (.A1_N(_11203_),
    .A2_N(_11279_),
    .B1(\design_top.MEM[17][11] ),
    .B2(_11281_),
    .X(_07081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12469_ (.A1_N(_11204_),
    .A2_N(_11278_),
    .B1(\design_top.MEM[17][10] ),
    .B2(_11280_),
    .X(_07080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12470_ (.A1_N(_11205_),
    .A2_N(_11278_),
    .B1(\design_top.MEM[17][9] ),
    .B2(_11280_),
    .X(_07079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12471_ (.A1_N(_11206_),
    .A2_N(_11278_),
    .B1(\design_top.MEM[17][8] ),
    .B2(_11280_),
    .X(_07078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12472_ (.A(_11212_),
    .B(_11106_),
    .X(_11282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12473_ (.A(_11282_),
    .X(_11283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12474_ (.A1(_11272_),
    .A2(_11113_),
    .B1(_11282_),
    .X(_11284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12475_ (.A(_11284_),
    .X(_11285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12476_ (.A1_N(_11211_),
    .A2_N(_11283_),
    .B1(\design_top.MEM[32][31] ),
    .B2(_11285_),
    .X(_07077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12477_ (.A1_N(_11218_),
    .A2_N(_11283_),
    .B1(\design_top.MEM[32][30] ),
    .B2(_11285_),
    .X(_07076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12478_ (.A1_N(_11219_),
    .A2_N(_11283_),
    .B1(\design_top.MEM[32][29] ),
    .B2(_11285_),
    .X(_07075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12479_ (.A1_N(_11220_),
    .A2_N(_11283_),
    .B1(\design_top.MEM[32][28] ),
    .B2(_11285_),
    .X(_07074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12480_ (.A1_N(_11221_),
    .A2_N(_11283_),
    .B1(\design_top.MEM[32][27] ),
    .B2(_11285_),
    .X(_07073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12481_ (.A1_N(_11222_),
    .A2_N(_11282_),
    .B1(\design_top.MEM[32][26] ),
    .B2(_11284_),
    .X(_07072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12482_ (.A1_N(_11223_),
    .A2_N(_11282_),
    .B1(\design_top.MEM[32][25] ),
    .B2(_11284_),
    .X(_07071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12483_ (.A1_N(_11224_),
    .A2_N(_11282_),
    .B1(\design_top.MEM[32][24] ),
    .B2(_11284_),
    .X(_07070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12484_ (.A(_11037_),
    .X(_11286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12485_ (.A(_11104_),
    .B(_11276_),
    .X(_11287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12486_ (.A(_11286_),
    .B(_11287_),
    .X(_11288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12487_ (.A(_11288_),
    .X(_11289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12488_ (.A1(_11197_),
    .A2(_11113_),
    .B1(_11288_),
    .X(_11290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12489_ (.A(_11290_),
    .X(_11291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12490_ (.A1_N(_11225_),
    .A2_N(_11289_),
    .B1(\design_top.MEM[33][15] ),
    .B2(_11291_),
    .X(_07069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12491_ (.A(_11046_),
    .X(_11292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12492_ (.A1_N(_11292_),
    .A2_N(_11289_),
    .B1(\design_top.MEM[33][14] ),
    .B2(_11291_),
    .X(_07068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12493_ (.A(_11048_),
    .X(_11293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12494_ (.A1_N(_11293_),
    .A2_N(_11289_),
    .B1(\design_top.MEM[33][13] ),
    .B2(_11291_),
    .X(_07067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12495_ (.A(_11050_),
    .X(_11294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12496_ (.A1_N(_11294_),
    .A2_N(_11289_),
    .B1(\design_top.MEM[33][12] ),
    .B2(_11291_),
    .X(_07066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12497_ (.A(_11052_),
    .X(_11295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12498_ (.A1_N(_11295_),
    .A2_N(_11289_),
    .B1(\design_top.MEM[33][11] ),
    .B2(_11291_),
    .X(_07065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12499_ (.A(_11054_),
    .X(_11296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12500_ (.A1_N(_11296_),
    .A2_N(_11288_),
    .B1(\design_top.MEM[33][10] ),
    .B2(_11290_),
    .X(_07064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12501_ (.A(_11056_),
    .X(_11297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12502_ (.A1_N(_11297_),
    .A2_N(_11288_),
    .B1(\design_top.MEM[33][9] ),
    .B2(_11290_),
    .X(_07063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12503_ (.A(_11058_),
    .X(_11298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12504_ (.A1_N(_11298_),
    .A2_N(_11288_),
    .B1(\design_top.MEM[33][8] ),
    .B2(_11290_),
    .X(_07062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12505_ (.A(_11060_),
    .X(_11299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12506_ (.A(_11025_),
    .X(_11300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12507_ (.A(_11300_),
    .B(_11287_),
    .X(_11301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12508_ (.A(_11301_),
    .X(_11302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12509_ (.A(_11196_),
    .X(_11303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12510_ (.A1(_11303_),
    .A2(_11113_),
    .B1(_11301_),
    .X(_11304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12511_ (.A(_11304_),
    .X(_11305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12512_ (.A1_N(_11299_),
    .A2_N(_11302_),
    .B1(\design_top.MEM[33][23] ),
    .B2(_11305_),
    .X(_07061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12513_ (.A(_11066_),
    .X(_11306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12514_ (.A1_N(_11306_),
    .A2_N(_11302_),
    .B1(\design_top.MEM[33][22] ),
    .B2(_11305_),
    .X(_07060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12515_ (.A(_11068_),
    .X(_11307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12516_ (.A1_N(_11307_),
    .A2_N(_11302_),
    .B1(\design_top.MEM[33][21] ),
    .B2(_11305_),
    .X(_07059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12517_ (.A(_11070_),
    .X(_11308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12518_ (.A1_N(_11308_),
    .A2_N(_11302_),
    .B1(\design_top.MEM[33][20] ),
    .B2(_11305_),
    .X(_07058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12519_ (.A(_11072_),
    .X(_11309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12520_ (.A1_N(_11309_),
    .A2_N(_11302_),
    .B1(\design_top.MEM[33][19] ),
    .B2(_11305_),
    .X(_07057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12521_ (.A(_11074_),
    .X(_11310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12522_ (.A1_N(_11310_),
    .A2_N(_11301_),
    .B1(\design_top.MEM[33][18] ),
    .B2(_11304_),
    .X(_07056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12523_ (.A(_11076_),
    .X(_11311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12524_ (.A1_N(_11311_),
    .A2_N(_11301_),
    .B1(\design_top.MEM[33][17] ),
    .B2(_11304_),
    .X(_07055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12525_ (.A(_11078_),
    .X(_11312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12526_ (.A1_N(_11312_),
    .A2_N(_11301_),
    .B1(\design_top.MEM[33][16] ),
    .B2(_11304_),
    .X(_07054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12527_ (.A(_11080_),
    .X(_11313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12528_ (.A(_11031_),
    .X(_11314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12529_ (.A(_11314_),
    .B(_11287_),
    .X(_11315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12530_ (.A(_11315_),
    .X(_11316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12531_ (.A(_11112_),
    .X(_11317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12532_ (.A1(_11303_),
    .A2(_11317_),
    .B1(_11315_),
    .X(_11318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12533_ (.A(_11318_),
    .X(_11319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12534_ (.A1_N(_11313_),
    .A2_N(_11316_),
    .B1(\design_top.MEM[33][31] ),
    .B2(_11319_),
    .X(_07053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12535_ (.A(_11086_),
    .X(_11320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12536_ (.A1_N(_11320_),
    .A2_N(_11316_),
    .B1(\design_top.MEM[33][30] ),
    .B2(_11319_),
    .X(_07052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12537_ (.A(_11088_),
    .X(_11321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12538_ (.A1_N(_11321_),
    .A2_N(_11316_),
    .B1(\design_top.MEM[33][29] ),
    .B2(_11319_),
    .X(_07051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12539_ (.A(_11090_),
    .X(_11322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12540_ (.A1_N(_11322_),
    .A2_N(_11316_),
    .B1(\design_top.MEM[33][28] ),
    .B2(_11319_),
    .X(_07050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12541_ (.A(_11092_),
    .X(_11323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12542_ (.A1_N(_11323_),
    .A2_N(_11316_),
    .B1(\design_top.MEM[33][27] ),
    .B2(_11319_),
    .X(_07049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12543_ (.A(_11094_),
    .X(_11324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12544_ (.A1_N(_11324_),
    .A2_N(_11315_),
    .B1(\design_top.MEM[33][26] ),
    .B2(_11318_),
    .X(_07048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12545_ (.A(_11096_),
    .X(_11325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12546_ (.A1_N(_11325_),
    .A2_N(_11315_),
    .B1(\design_top.MEM[33][25] ),
    .B2(_11318_),
    .X(_07047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12547_ (.A(_11098_),
    .X(_11326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12548_ (.A1_N(_11326_),
    .A2_N(_11315_),
    .B1(\design_top.MEM[33][24] ),
    .B2(_11318_),
    .X(_07046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12549_ (.A(_11000_),
    .B(_11105_),
    .X(_11327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12550_ (.A(_11314_),
    .B(_11327_),
    .X(_11328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12551_ (.A(_11328_),
    .X(_11329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12552_ (.A1(_11237_),
    .A2(_11317_),
    .B1(_11328_),
    .X(_11330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12553_ (.A(_11330_),
    .X(_11331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12554_ (.A1_N(_11313_),
    .A2_N(_11329_),
    .B1(\design_top.MEM[34][31] ),
    .B2(_11331_),
    .X(_07045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12555_ (.A1_N(_11320_),
    .A2_N(_11329_),
    .B1(\design_top.MEM[34][30] ),
    .B2(_11331_),
    .X(_07044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12556_ (.A1_N(_11321_),
    .A2_N(_11329_),
    .B1(\design_top.MEM[34][29] ),
    .B2(_11331_),
    .X(_07043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12557_ (.A1_N(_11322_),
    .A2_N(_11329_),
    .B1(\design_top.MEM[34][28] ),
    .B2(_11331_),
    .X(_07042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12558_ (.A1_N(_11323_),
    .A2_N(_11329_),
    .B1(\design_top.MEM[34][27] ),
    .B2(_11331_),
    .X(_07041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12559_ (.A1_N(_11324_),
    .A2_N(_11328_),
    .B1(\design_top.MEM[34][26] ),
    .B2(_11330_),
    .X(_07040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12560_ (.A1_N(_11325_),
    .A2_N(_11328_),
    .B1(\design_top.MEM[34][25] ),
    .B2(_11330_),
    .X(_07039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12561_ (.A1_N(_11326_),
    .A2_N(_11328_),
    .B1(\design_top.MEM[34][24] ),
    .B2(_11330_),
    .X(_07038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12562_ (.A(_11300_),
    .B(_11277_),
    .X(_11332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12563_ (.A(_11332_),
    .X(_11333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12564_ (.A1(_11303_),
    .A2(_11262_),
    .B1(_11332_),
    .X(_11334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12565_ (.A(_11334_),
    .X(_11335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12566_ (.A1_N(_11299_),
    .A2_N(_11333_),
    .B1(\design_top.MEM[17][23] ),
    .B2(_11335_),
    .X(_07037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12567_ (.A1_N(_11306_),
    .A2_N(_11333_),
    .B1(\design_top.MEM[17][22] ),
    .B2(_11335_),
    .X(_07036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12568_ (.A1_N(_11307_),
    .A2_N(_11333_),
    .B1(\design_top.MEM[17][21] ),
    .B2(_11335_),
    .X(_07035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12569_ (.A1_N(_11308_),
    .A2_N(_11333_),
    .B1(\design_top.MEM[17][20] ),
    .B2(_11335_),
    .X(_07034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12570_ (.A1_N(_11309_),
    .A2_N(_11333_),
    .B1(\design_top.MEM[17][19] ),
    .B2(_11335_),
    .X(_07033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12571_ (.A1_N(_11310_),
    .A2_N(_11332_),
    .B1(\design_top.MEM[17][18] ),
    .B2(_11334_),
    .X(_07032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12572_ (.A1_N(_11311_),
    .A2_N(_11332_),
    .B1(\design_top.MEM[17][17] ),
    .B2(_11334_),
    .X(_07031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12573_ (.A1_N(_11312_),
    .A2_N(_11332_),
    .B1(\design_top.MEM[17][16] ),
    .B2(_11334_),
    .X(_07030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12574_ (.A(_11314_),
    .B(_11277_),
    .X(_11336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12575_ (.A(_11336_),
    .X(_11337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12576_ (.A(_11261_),
    .X(_11338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12577_ (.A1(_11303_),
    .A2(_11338_),
    .B1(_11336_),
    .X(_11339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12578_ (.A(_11339_),
    .X(_11340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12579_ (.A1_N(_11313_),
    .A2_N(_11337_),
    .B1(\design_top.MEM[17][31] ),
    .B2(_11340_),
    .X(_07029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12580_ (.A1_N(_11320_),
    .A2_N(_11337_),
    .B1(\design_top.MEM[17][30] ),
    .B2(_11340_),
    .X(_07028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12581_ (.A1_N(_11321_),
    .A2_N(_11337_),
    .B1(\design_top.MEM[17][29] ),
    .B2(_11340_),
    .X(_07027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12582_ (.A1_N(_11322_),
    .A2_N(_11337_),
    .B1(\design_top.MEM[17][28] ),
    .B2(_11340_),
    .X(_07026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12583_ (.A1_N(_11323_),
    .A2_N(_11337_),
    .B1(\design_top.MEM[17][27] ),
    .B2(_11340_),
    .X(_07025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12584_ (.A1_N(_11324_),
    .A2_N(_11336_),
    .B1(\design_top.MEM[17][26] ),
    .B2(_11339_),
    .X(_07024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12585_ (.A1_N(_11325_),
    .A2_N(_11336_),
    .B1(\design_top.MEM[17][25] ),
    .B2(_11339_),
    .X(_07023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12586_ (.A1_N(_11326_),
    .A2_N(_11336_),
    .B1(\design_top.MEM[17][24] ),
    .B2(_11339_),
    .X(_07022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12587_ (.A(_11100_),
    .X(_11341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12588_ (.A(_11000_),
    .B(_11256_),
    .X(_11342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12589_ (.A(_11286_),
    .B(_11342_),
    .X(_11343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12590_ (.A(_11343_),
    .X(_11344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12591_ (.A1(_11237_),
    .A2(_11338_),
    .B1(_11343_),
    .X(_11345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12592_ (.A(_11345_),
    .X(_11346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12593_ (.A1_N(_11341_),
    .A2_N(_11344_),
    .B1(\design_top.MEM[18][15] ),
    .B2(_11346_),
    .X(_07021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12594_ (.A1_N(_11292_),
    .A2_N(_11344_),
    .B1(\design_top.MEM[18][14] ),
    .B2(_11346_),
    .X(_07020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12595_ (.A1_N(_11293_),
    .A2_N(_11344_),
    .B1(\design_top.MEM[18][13] ),
    .B2(_11346_),
    .X(_07019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12596_ (.A1_N(_11294_),
    .A2_N(_11344_),
    .B1(\design_top.MEM[18][12] ),
    .B2(_11346_),
    .X(_07018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12597_ (.A1_N(_11295_),
    .A2_N(_11344_),
    .B1(\design_top.MEM[18][11] ),
    .B2(_11346_),
    .X(_07017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12598_ (.A1_N(_11296_),
    .A2_N(_11343_),
    .B1(\design_top.MEM[18][10] ),
    .B2(_11345_),
    .X(_07016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12599_ (.A1_N(_11297_),
    .A2_N(_11343_),
    .B1(\design_top.MEM[18][9] ),
    .B2(_11345_),
    .X(_07015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12600_ (.A1_N(_11298_),
    .A2_N(_11343_),
    .B1(\design_top.MEM[18][8] ),
    .B2(_11345_),
    .X(_07014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12601_ (.A(_11300_),
    .B(_11342_),
    .X(_11347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12602_ (.A(_11347_),
    .X(_11348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12603_ (.A1(_11237_),
    .A2(_11338_),
    .B1(_11347_),
    .X(_11349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12604_ (.A(_11349_),
    .X(_11350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12605_ (.A1_N(_11299_),
    .A2_N(_11348_),
    .B1(\design_top.MEM[18][23] ),
    .B2(_11350_),
    .X(_07013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12606_ (.A1_N(_11306_),
    .A2_N(_11348_),
    .B1(\design_top.MEM[18][22] ),
    .B2(_11350_),
    .X(_07012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12607_ (.A1_N(_11307_),
    .A2_N(_11348_),
    .B1(\design_top.MEM[18][21] ),
    .B2(_11350_),
    .X(_07011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12608_ (.A1_N(_11308_),
    .A2_N(_11348_),
    .B1(\design_top.MEM[18][20] ),
    .B2(_11350_),
    .X(_07010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12609_ (.A1_N(_11309_),
    .A2_N(_11348_),
    .B1(\design_top.MEM[18][19] ),
    .B2(_11350_),
    .X(_07009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12610_ (.A1_N(_11310_),
    .A2_N(_11347_),
    .B1(\design_top.MEM[18][18] ),
    .B2(_11349_),
    .X(_07008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12611_ (.A1_N(_11311_),
    .A2_N(_11347_),
    .B1(\design_top.MEM[18][17] ),
    .B2(_11349_),
    .X(_07007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12612_ (.A1_N(_11312_),
    .A2_N(_11347_),
    .B1(\design_top.MEM[18][16] ),
    .B2(_11349_),
    .X(_07006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12613_ (.A(_11314_),
    .B(_11342_),
    .X(_11351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12614_ (.A(_11351_),
    .X(_11352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12615_ (.A1(_11237_),
    .A2(_11338_),
    .B1(_11351_),
    .X(_11353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12616_ (.A(_11353_),
    .X(_11354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12617_ (.A1_N(_11313_),
    .A2_N(_11352_),
    .B1(\design_top.MEM[18][31] ),
    .B2(_11354_),
    .X(_07005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12618_ (.A1_N(_11320_),
    .A2_N(_11352_),
    .B1(\design_top.MEM[18][30] ),
    .B2(_11354_),
    .X(_07004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12619_ (.A1_N(_11321_),
    .A2_N(_11352_),
    .B1(\design_top.MEM[18][29] ),
    .B2(_11354_),
    .X(_07003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12620_ (.A1_N(_11322_),
    .A2_N(_11352_),
    .B1(\design_top.MEM[18][28] ),
    .B2(_11354_),
    .X(_07002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12621_ (.A1_N(_11323_),
    .A2_N(_11352_),
    .B1(\design_top.MEM[18][27] ),
    .B2(_11354_),
    .X(_07001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12622_ (.A1_N(_11324_),
    .A2_N(_11351_),
    .B1(\design_top.MEM[18][26] ),
    .B2(_11353_),
    .X(_07000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12623_ (.A1_N(_11325_),
    .A2_N(_11351_),
    .B1(\design_top.MEM[18][25] ),
    .B2(_11353_),
    .X(_06999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12624_ (.A1_N(_11326_),
    .A2_N(_11351_),
    .B1(\design_top.MEM[18][24] ),
    .B2(_11353_),
    .X(_06998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12625_ (.A(_10885_),
    .B(_11256_),
    .X(_11355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12626_ (.A(_11286_),
    .B(_11355_),
    .X(_11356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12627_ (.A(_11356_),
    .X(_11357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12628_ (.A1(_11252_),
    .A2(_11338_),
    .B1(_11356_),
    .X(_11358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12629_ (.A(_11358_),
    .X(_11359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12630_ (.A1_N(_11341_),
    .A2_N(_11357_),
    .B1(\design_top.MEM[19][15] ),
    .B2(_11359_),
    .X(_06997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12631_ (.A1_N(_11292_),
    .A2_N(_11357_),
    .B1(\design_top.MEM[19][14] ),
    .B2(_11359_),
    .X(_06996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12632_ (.A1_N(_11293_),
    .A2_N(_11357_),
    .B1(\design_top.MEM[19][13] ),
    .B2(_11359_),
    .X(_06995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12633_ (.A1_N(_11294_),
    .A2_N(_11357_),
    .B1(\design_top.MEM[19][12] ),
    .B2(_11359_),
    .X(_06994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12634_ (.A1_N(_11295_),
    .A2_N(_11357_),
    .B1(\design_top.MEM[19][11] ),
    .B2(_11359_),
    .X(_06993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12635_ (.A1_N(_11296_),
    .A2_N(_11356_),
    .B1(\design_top.MEM[19][10] ),
    .B2(_11358_),
    .X(_06992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12636_ (.A1_N(_11297_),
    .A2_N(_11356_),
    .B1(\design_top.MEM[19][9] ),
    .B2(_11358_),
    .X(_06991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12637_ (.A1_N(_11298_),
    .A2_N(_11356_),
    .B1(\design_top.MEM[19][8] ),
    .B2(_11358_),
    .X(_06990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12638_ (.A(_11300_),
    .B(_11355_),
    .X(_11360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12639_ (.A(_11360_),
    .X(_11361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12640_ (.A1(_11252_),
    .A2(_11261_),
    .B1(_11360_),
    .X(_11362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12641_ (.A(_11362_),
    .X(_11363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12642_ (.A1_N(_11299_),
    .A2_N(_11361_),
    .B1(\design_top.MEM[19][23] ),
    .B2(_11363_),
    .X(_06989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12643_ (.A1_N(_11306_),
    .A2_N(_11361_),
    .B1(\design_top.MEM[19][22] ),
    .B2(_11363_),
    .X(_06988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12644_ (.A1_N(_11307_),
    .A2_N(_11361_),
    .B1(\design_top.MEM[19][21] ),
    .B2(_11363_),
    .X(_06987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12645_ (.A1_N(_11308_),
    .A2_N(_11361_),
    .B1(\design_top.MEM[19][20] ),
    .B2(_11363_),
    .X(_06986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12646_ (.A1_N(_11309_),
    .A2_N(_11361_),
    .B1(\design_top.MEM[19][19] ),
    .B2(_11363_),
    .X(_06985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12647_ (.A1_N(_11310_),
    .A2_N(_11360_),
    .B1(\design_top.MEM[19][18] ),
    .B2(_11362_),
    .X(_06984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12648_ (.A1_N(_11311_),
    .A2_N(_11360_),
    .B1(\design_top.MEM[19][17] ),
    .B2(_11362_),
    .X(_06983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12649_ (.A1_N(_11312_),
    .A2_N(_11360_),
    .B1(\design_top.MEM[19][16] ),
    .B2(_11362_),
    .X(_06982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12650_ (.A(_11314_),
    .B(_11355_),
    .X(_11364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12651_ (.A(_11364_),
    .X(_11365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12652_ (.A1(_11252_),
    .A2(_11261_),
    .B1(_11364_),
    .X(_11366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12653_ (.A(_11366_),
    .X(_11367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12654_ (.A1_N(_11313_),
    .A2_N(_11365_),
    .B1(\design_top.MEM[19][31] ),
    .B2(_11367_),
    .X(_06981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12655_ (.A1_N(_11320_),
    .A2_N(_11365_),
    .B1(\design_top.MEM[19][30] ),
    .B2(_11367_),
    .X(_06980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12656_ (.A1_N(_11321_),
    .A2_N(_11365_),
    .B1(\design_top.MEM[19][29] ),
    .B2(_11367_),
    .X(_06979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12657_ (.A1_N(_11322_),
    .A2_N(_11365_),
    .B1(\design_top.MEM[19][28] ),
    .B2(_11367_),
    .X(_06978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12658_ (.A1_N(_11323_),
    .A2_N(_11365_),
    .B1(\design_top.MEM[19][27] ),
    .B2(_11367_),
    .X(_06977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12659_ (.A1_N(_11324_),
    .A2_N(_11364_),
    .B1(\design_top.MEM[19][26] ),
    .B2(_11366_),
    .X(_06976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12660_ (.A1_N(_11325_),
    .A2_N(_11364_),
    .B1(\design_top.MEM[19][25] ),
    .B2(_11366_),
    .X(_06975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12661_ (.A1_N(_11326_),
    .A2_N(_11364_),
    .B1(\design_top.MEM[19][24] ),
    .B2(_11366_),
    .X(_06974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12662_ (.A(_11286_),
    .B(_11327_),
    .X(_07432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12663_ (.A(_07432_),
    .X(_07433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12664_ (.A(_11134_),
    .X(_07434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12665_ (.A(_07434_),
    .X(_07435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12666_ (.A1(_07435_),
    .A2(_11317_),
    .B1(_07432_),
    .X(_07436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12667_ (.A(_07436_),
    .X(_07437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12668_ (.A1_N(_11341_),
    .A2_N(_07433_),
    .B1(\design_top.MEM[34][15] ),
    .B2(_07437_),
    .X(_06973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12669_ (.A1_N(_11292_),
    .A2_N(_07433_),
    .B1(\design_top.MEM[34][14] ),
    .B2(_07437_),
    .X(_06972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12670_ (.A1_N(_11293_),
    .A2_N(_07433_),
    .B1(\design_top.MEM[34][13] ),
    .B2(_07437_),
    .X(_06971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12671_ (.A1_N(_11294_),
    .A2_N(_07433_),
    .B1(\design_top.MEM[34][12] ),
    .B2(_07437_),
    .X(_06970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12672_ (.A1_N(_11295_),
    .A2_N(_07433_),
    .B1(\design_top.MEM[34][11] ),
    .B2(_07437_),
    .X(_06969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12673_ (.A1_N(_11296_),
    .A2_N(_07432_),
    .B1(\design_top.MEM[34][10] ),
    .B2(_07436_),
    .X(_06968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12674_ (.A1_N(_11297_),
    .A2_N(_07432_),
    .B1(\design_top.MEM[34][9] ),
    .B2(_07436_),
    .X(_06967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12675_ (.A1_N(_11298_),
    .A2_N(_07432_),
    .B1(\design_top.MEM[34][8] ),
    .B2(_07436_),
    .X(_06966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12676_ (.A(_11300_),
    .B(_11327_),
    .X(_07438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12677_ (.A(_07438_),
    .X(_07439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12678_ (.A1(_07435_),
    .A2(_11317_),
    .B1(_07438_),
    .X(_07440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12679_ (.A(_07440_),
    .X(_07441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12680_ (.A1_N(_11299_),
    .A2_N(_07439_),
    .B1(\design_top.MEM[34][23] ),
    .B2(_07441_),
    .X(_06965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12681_ (.A1_N(_11306_),
    .A2_N(_07439_),
    .B1(\design_top.MEM[34][22] ),
    .B2(_07441_),
    .X(_06964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12682_ (.A1_N(_11307_),
    .A2_N(_07439_),
    .B1(\design_top.MEM[34][21] ),
    .B2(_07441_),
    .X(_06963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12683_ (.A1_N(_11308_),
    .A2_N(_07439_),
    .B1(\design_top.MEM[34][20] ),
    .B2(_07441_),
    .X(_06962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12684_ (.A1_N(_11309_),
    .A2_N(_07439_),
    .B1(\design_top.MEM[34][19] ),
    .B2(_07441_),
    .X(_06961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12685_ (.A1_N(_11310_),
    .A2_N(_07438_),
    .B1(\design_top.MEM[34][18] ),
    .B2(_07440_),
    .X(_06960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12686_ (.A1_N(_11311_),
    .A2_N(_07438_),
    .B1(\design_top.MEM[34][17] ),
    .B2(_07440_),
    .X(_06959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12687_ (.A1_N(_11312_),
    .A2_N(_07438_),
    .B1(\design_top.MEM[34][16] ),
    .B2(_07440_),
    .X(_06958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12688_ (.A(_10885_),
    .B(_11105_),
    .X(_07442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12689_ (.A(_11286_),
    .B(_07442_),
    .X(_07443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12690_ (.A(_07443_),
    .X(_07444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12691_ (.A1(_11252_),
    .A2(_11317_),
    .B1(_07443_),
    .X(_07445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12692_ (.A(_07445_),
    .X(_07446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12693_ (.A1_N(_11341_),
    .A2_N(_07444_),
    .B1(\design_top.MEM[35][15] ),
    .B2(_07446_),
    .X(_06957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12694_ (.A1_N(_11292_),
    .A2_N(_07444_),
    .B1(\design_top.MEM[35][14] ),
    .B2(_07446_),
    .X(_06956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12695_ (.A1_N(_11293_),
    .A2_N(_07444_),
    .B1(\design_top.MEM[35][13] ),
    .B2(_07446_),
    .X(_06955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12696_ (.A1_N(_11294_),
    .A2_N(_07444_),
    .B1(\design_top.MEM[35][12] ),
    .B2(_07446_),
    .X(_06954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12697_ (.A1_N(_11295_),
    .A2_N(_07444_),
    .B1(\design_top.MEM[35][11] ),
    .B2(_07446_),
    .X(_06953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12698_ (.A1_N(_11296_),
    .A2_N(_07443_),
    .B1(\design_top.MEM[35][10] ),
    .B2(_07445_),
    .X(_06952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12699_ (.A1_N(_11297_),
    .A2_N(_07443_),
    .B1(\design_top.MEM[35][9] ),
    .B2(_07445_),
    .X(_06951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12700_ (.A1_N(_11298_),
    .A2_N(_07443_),
    .B1(\design_top.MEM[35][8] ),
    .B2(_07445_),
    .X(_06950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12701_ (.A(_11060_),
    .X(_07447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12702_ (.A(_11025_),
    .X(_07448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12703_ (.A(_02860_),
    .B(_11103_),
    .X(_07449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12704_ (.A(_07449_),
    .X(_07450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12705_ (.A(_10980_),
    .B(_07450_),
    .X(_07451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12706_ (.A(_07448_),
    .B(_07451_),
    .X(_07452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12707_ (.A(_07452_),
    .X(_07453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _12708_ (.A(_11110_),
    .B(_10788_),
    .C(_10896_),
    .D(_10964_),
    .X(_07454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12709_ (.A(_07454_),
    .X(_07455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12710_ (.A(_07455_),
    .X(_07456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12711_ (.A1(_11303_),
    .A2(_07456_),
    .B1(_07452_),
    .X(_07457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12712_ (.A(_07457_),
    .X(_07458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12713_ (.A1_N(_07447_),
    .A2_N(_07453_),
    .B1(\design_top.MEM[45][23] ),
    .B2(_07458_),
    .X(_06949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12714_ (.A(_11066_),
    .X(_07459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12715_ (.A1_N(_07459_),
    .A2_N(_07453_),
    .B1(\design_top.MEM[45][22] ),
    .B2(_07458_),
    .X(_06948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12716_ (.A(_11068_),
    .X(_07460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12717_ (.A1_N(_07460_),
    .A2_N(_07453_),
    .B1(\design_top.MEM[45][21] ),
    .B2(_07458_),
    .X(_06947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12718_ (.A(_11070_),
    .X(_07461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12719_ (.A1_N(_07461_),
    .A2_N(_07453_),
    .B1(\design_top.MEM[45][20] ),
    .B2(_07458_),
    .X(_06946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12720_ (.A(_11072_),
    .X(_07462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12721_ (.A1_N(_07462_),
    .A2_N(_07453_),
    .B1(\design_top.MEM[45][19] ),
    .B2(_07458_),
    .X(_06945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12722_ (.A(_11074_),
    .X(_07463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12723_ (.A1_N(_07463_),
    .A2_N(_07452_),
    .B1(\design_top.MEM[45][18] ),
    .B2(_07457_),
    .X(_06944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12724_ (.A(_11076_),
    .X(_07464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12725_ (.A1_N(_07464_),
    .A2_N(_07452_),
    .B1(\design_top.MEM[45][17] ),
    .B2(_07457_),
    .X(_06943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12726_ (.A(_11078_),
    .X(_07465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12727_ (.A1_N(_07465_),
    .A2_N(_07452_),
    .B1(\design_top.MEM[45][16] ),
    .B2(_07457_),
    .X(_06942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12728_ (.A(_07448_),
    .B(_07442_),
    .X(_07466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12729_ (.A(_07466_),
    .X(_07467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12730_ (.A(_11251_),
    .X(_07468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12731_ (.A1(_07468_),
    .A2(_11112_),
    .B1(_07466_),
    .X(_07469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12732_ (.A(_07469_),
    .X(_07470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12733_ (.A1_N(_07447_),
    .A2_N(_07467_),
    .B1(\design_top.MEM[35][23] ),
    .B2(_07470_),
    .X(_06941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12734_ (.A1_N(_07459_),
    .A2_N(_07467_),
    .B1(\design_top.MEM[35][22] ),
    .B2(_07470_),
    .X(_06940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12735_ (.A1_N(_07460_),
    .A2_N(_07467_),
    .B1(\design_top.MEM[35][21] ),
    .B2(_07470_),
    .X(_06939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12736_ (.A1_N(_07461_),
    .A2_N(_07467_),
    .B1(\design_top.MEM[35][20] ),
    .B2(_07470_),
    .X(_06938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12737_ (.A1_N(_07462_),
    .A2_N(_07467_),
    .B1(\design_top.MEM[35][19] ),
    .B2(_07470_),
    .X(_06937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12738_ (.A1_N(_07463_),
    .A2_N(_07466_),
    .B1(\design_top.MEM[35][18] ),
    .B2(_07469_),
    .X(_06936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12739_ (.A1_N(_07464_),
    .A2_N(_07466_),
    .B1(\design_top.MEM[35][17] ),
    .B2(_07469_),
    .X(_06935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12740_ (.A1_N(_07465_),
    .A2_N(_07466_),
    .B1(\design_top.MEM[35][16] ),
    .B2(_07469_),
    .X(_06934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12741_ (.A(_11037_),
    .X(_07471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12742_ (.A(_10958_),
    .B(_11256_),
    .X(_07472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12743_ (.A(_07471_),
    .B(_07472_),
    .X(_07473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12744_ (.A(_07473_),
    .X(_07474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _12745_ (.A(wbs_adr_i[3]),
    .B(_10894_),
    .C(_10789_),
    .D(_10964_),
    .X(_07475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12746_ (.A(_07475_),
    .X(_07476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12747_ (.A(_07476_),
    .X(_07477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12748_ (.A1(_11272_),
    .A2(_07477_),
    .B1(_07473_),
    .X(_07478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12749_ (.A(_07478_),
    .X(_07479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12750_ (.A1_N(_11341_),
    .A2_N(_07474_),
    .B1(\design_top.MEM[20][15] ),
    .B2(_07479_),
    .X(_06933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12751_ (.A(_11046_),
    .X(_07480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12752_ (.A1_N(_07480_),
    .A2_N(_07474_),
    .B1(\design_top.MEM[20][14] ),
    .B2(_07479_),
    .X(_06932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12753_ (.A(_11048_),
    .X(_07481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12754_ (.A1_N(_07481_),
    .A2_N(_07474_),
    .B1(\design_top.MEM[20][13] ),
    .B2(_07479_),
    .X(_06931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12755_ (.A(_11050_),
    .X(_07482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12756_ (.A1_N(_07482_),
    .A2_N(_07474_),
    .B1(\design_top.MEM[20][12] ),
    .B2(_07479_),
    .X(_06930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12757_ (.A(_11052_),
    .X(_07483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12758_ (.A1_N(_07483_),
    .A2_N(_07474_),
    .B1(\design_top.MEM[20][11] ),
    .B2(_07479_),
    .X(_06929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12759_ (.A(_11054_),
    .X(_07484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12760_ (.A1_N(_07484_),
    .A2_N(_07473_),
    .B1(\design_top.MEM[20][10] ),
    .B2(_07478_),
    .X(_06928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12761_ (.A(_11056_),
    .X(_07485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12762_ (.A1_N(_07485_),
    .A2_N(_07473_),
    .B1(\design_top.MEM[20][9] ),
    .B2(_07478_),
    .X(_06927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12763_ (.A(_11058_),
    .X(_07486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12764_ (.A1_N(_07486_),
    .A2_N(_07473_),
    .B1(\design_top.MEM[20][8] ),
    .B2(_07478_),
    .X(_06926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12765_ (.A(_11080_),
    .X(_07487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12766_ (.A(_11031_),
    .X(_07488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12767_ (.A(_07488_),
    .B(_07442_),
    .X(_07489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12768_ (.A(_07489_),
    .X(_07490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12769_ (.A1(_07468_),
    .A2(_11112_),
    .B1(_07489_),
    .X(_07491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12770_ (.A(_07491_),
    .X(_07492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12771_ (.A1_N(_07487_),
    .A2_N(_07490_),
    .B1(\design_top.MEM[35][31] ),
    .B2(_07492_),
    .X(_06925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12772_ (.A(_11086_),
    .X(_07493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12773_ (.A1_N(_07493_),
    .A2_N(_07490_),
    .B1(\design_top.MEM[35][30] ),
    .B2(_07492_),
    .X(_06924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12774_ (.A(_11088_),
    .X(_07494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12775_ (.A1_N(_07494_),
    .A2_N(_07490_),
    .B1(\design_top.MEM[35][29] ),
    .B2(_07492_),
    .X(_06923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12776_ (.A(_11090_),
    .X(_07495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12777_ (.A1_N(_07495_),
    .A2_N(_07490_),
    .B1(\design_top.MEM[35][28] ),
    .B2(_07492_),
    .X(_06922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12778_ (.A(_11092_),
    .X(_07496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12779_ (.A1_N(_07496_),
    .A2_N(_07490_),
    .B1(\design_top.MEM[35][27] ),
    .B2(_07492_),
    .X(_06921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12780_ (.A(_11094_),
    .X(_07497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12781_ (.A1_N(_07497_),
    .A2_N(_07489_),
    .B1(\design_top.MEM[35][26] ),
    .B2(_07491_),
    .X(_06920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12782_ (.A(_11096_),
    .X(_07498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12783_ (.A1_N(_07498_),
    .A2_N(_07489_),
    .B1(\design_top.MEM[35][25] ),
    .B2(_07491_),
    .X(_06919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12784_ (.A(_11098_),
    .X(_07499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12785_ (.A1_N(_07499_),
    .A2_N(_07489_),
    .B1(\design_top.MEM[35][24] ),
    .B2(_07491_),
    .X(_06918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12786_ (.A(_07448_),
    .B(_07472_),
    .X(_07500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12787_ (.A(_07500_),
    .X(_07501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12788_ (.A1(_11272_),
    .A2(_07477_),
    .B1(_07500_),
    .X(_07502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12789_ (.A(_07502_),
    .X(_07503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12790_ (.A1_N(_07447_),
    .A2_N(_07501_),
    .B1(\design_top.MEM[20][23] ),
    .B2(_07503_),
    .X(_06917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12791_ (.A1_N(_07459_),
    .A2_N(_07501_),
    .B1(\design_top.MEM[20][22] ),
    .B2(_07503_),
    .X(_06916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12792_ (.A1_N(_07460_),
    .A2_N(_07501_),
    .B1(\design_top.MEM[20][21] ),
    .B2(_07503_),
    .X(_06915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12793_ (.A1_N(_07461_),
    .A2_N(_07501_),
    .B1(\design_top.MEM[20][20] ),
    .B2(_07503_),
    .X(_06914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12794_ (.A1_N(_07462_),
    .A2_N(_07501_),
    .B1(\design_top.MEM[20][19] ),
    .B2(_07503_),
    .X(_06913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12795_ (.A1_N(_07463_),
    .A2_N(_07500_),
    .B1(\design_top.MEM[20][18] ),
    .B2(_07502_),
    .X(_06912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12796_ (.A1_N(_07464_),
    .A2_N(_07500_),
    .B1(\design_top.MEM[20][17] ),
    .B2(_07502_),
    .X(_06911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12797_ (.A1_N(_07465_),
    .A2_N(_07500_),
    .B1(\design_top.MEM[20][16] ),
    .B2(_07502_),
    .X(_06910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12798_ (.A(_11100_),
    .X(_07504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12799_ (.A(_10980_),
    .B(_11256_),
    .X(_07505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12800_ (.A(_07471_),
    .B(_07505_),
    .X(_07506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12801_ (.A(_07506_),
    .X(_07507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12802_ (.A(_11195_),
    .X(_07508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12803_ (.A(_07508_),
    .X(_07509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12804_ (.A1(_07509_),
    .A2(_07477_),
    .B1(_07506_),
    .X(_07510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12805_ (.A(_07510_),
    .X(_07511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12806_ (.A1_N(_07504_),
    .A2_N(_07507_),
    .B1(\design_top.MEM[21][15] ),
    .B2(_07511_),
    .X(_06909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12807_ (.A1_N(_07480_),
    .A2_N(_07507_),
    .B1(\design_top.MEM[21][14] ),
    .B2(_07511_),
    .X(_06908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12808_ (.A1_N(_07481_),
    .A2_N(_07507_),
    .B1(\design_top.MEM[21][13] ),
    .B2(_07511_),
    .X(_06907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12809_ (.A1_N(_07482_),
    .A2_N(_07507_),
    .B1(\design_top.MEM[21][12] ),
    .B2(_07511_),
    .X(_06906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12810_ (.A1_N(_07483_),
    .A2_N(_07507_),
    .B1(\design_top.MEM[21][11] ),
    .B2(_07511_),
    .X(_06905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12811_ (.A1_N(_07484_),
    .A2_N(_07506_),
    .B1(\design_top.MEM[21][10] ),
    .B2(_07510_),
    .X(_06904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12812_ (.A1_N(_07485_),
    .A2_N(_07506_),
    .B1(\design_top.MEM[21][9] ),
    .B2(_07510_),
    .X(_06903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12813_ (.A1_N(_07486_),
    .A2_N(_07506_),
    .B1(\design_top.MEM[21][8] ),
    .B2(_07510_),
    .X(_06902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12814_ (.A(_07448_),
    .B(_07505_),
    .X(_07512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12815_ (.A(_07512_),
    .X(_07513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12816_ (.A1(_07509_),
    .A2(_07477_),
    .B1(_07512_),
    .X(_07514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12817_ (.A(_07514_),
    .X(_07515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12818_ (.A1_N(_07447_),
    .A2_N(_07513_),
    .B1(\design_top.MEM[21][23] ),
    .B2(_07515_),
    .X(_06901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12819_ (.A1_N(_07459_),
    .A2_N(_07513_),
    .B1(\design_top.MEM[21][22] ),
    .B2(_07515_),
    .X(_06900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12820_ (.A1_N(_07460_),
    .A2_N(_07513_),
    .B1(\design_top.MEM[21][21] ),
    .B2(_07515_),
    .X(_06899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12821_ (.A1_N(_07461_),
    .A2_N(_07513_),
    .B1(\design_top.MEM[21][20] ),
    .B2(_07515_),
    .X(_06898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12822_ (.A1_N(_07462_),
    .A2_N(_07513_),
    .B1(\design_top.MEM[21][19] ),
    .B2(_07515_),
    .X(_06897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12823_ (.A1_N(_07463_),
    .A2_N(_07512_),
    .B1(\design_top.MEM[21][18] ),
    .B2(_07514_),
    .X(_06896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12824_ (.A1_N(_07464_),
    .A2_N(_07512_),
    .B1(\design_top.MEM[21][17] ),
    .B2(_07514_),
    .X(_06895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12825_ (.A1_N(_07465_),
    .A2_N(_07512_),
    .B1(\design_top.MEM[21][16] ),
    .B2(_07514_),
    .X(_06894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12826_ (.A(_10958_),
    .B(_11105_),
    .X(_07516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12827_ (.A(_07471_),
    .B(_07516_),
    .X(_07517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12828_ (.A(_07517_),
    .X(_07518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _12829_ (.A(_11110_),
    .B(wbs_adr_i[2]),
    .C(_10789_),
    .D(_10964_),
    .X(_07519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12830_ (.A(_07519_),
    .X(_07520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12831_ (.A(_07520_),
    .X(_07521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12832_ (.A1(_11272_),
    .A2(_07521_),
    .B1(_07517_),
    .X(_07522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12833_ (.A(_07522_),
    .X(_07523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12834_ (.A1_N(_07504_),
    .A2_N(_07518_),
    .B1(\design_top.MEM[36][15] ),
    .B2(_07523_),
    .X(_06893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12835_ (.A1_N(_07480_),
    .A2_N(_07518_),
    .B1(\design_top.MEM[36][14] ),
    .B2(_07523_),
    .X(_06892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12836_ (.A1_N(_07481_),
    .A2_N(_07518_),
    .B1(\design_top.MEM[36][13] ),
    .B2(_07523_),
    .X(_06891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12837_ (.A1_N(_07482_),
    .A2_N(_07518_),
    .B1(\design_top.MEM[36][12] ),
    .B2(_07523_),
    .X(_06890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12838_ (.A1_N(_07483_),
    .A2_N(_07518_),
    .B1(\design_top.MEM[36][11] ),
    .B2(_07523_),
    .X(_06889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12839_ (.A1_N(_07484_),
    .A2_N(_07517_),
    .B1(\design_top.MEM[36][10] ),
    .B2(_07522_),
    .X(_06888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12840_ (.A1_N(_07485_),
    .A2_N(_07517_),
    .B1(\design_top.MEM[36][9] ),
    .B2(_07522_),
    .X(_06887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12841_ (.A1_N(_07486_),
    .A2_N(_07517_),
    .B1(\design_top.MEM[36][8] ),
    .B2(_07522_),
    .X(_06886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12842_ (.A(_07488_),
    .B(_07505_),
    .X(_07524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12843_ (.A(_07524_),
    .X(_07525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12844_ (.A1(_07509_),
    .A2(_07477_),
    .B1(_07524_),
    .X(_07526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12845_ (.A(_07526_),
    .X(_07527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12846_ (.A1_N(_07487_),
    .A2_N(_07525_),
    .B1(\design_top.MEM[21][31] ),
    .B2(_07527_),
    .X(_06885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12847_ (.A1_N(_07493_),
    .A2_N(_07525_),
    .B1(\design_top.MEM[21][30] ),
    .B2(_07527_),
    .X(_06884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12848_ (.A1_N(_07494_),
    .A2_N(_07525_),
    .B1(\design_top.MEM[21][29] ),
    .B2(_07527_),
    .X(_06883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12849_ (.A1_N(_07495_),
    .A2_N(_07525_),
    .B1(\design_top.MEM[21][28] ),
    .B2(_07527_),
    .X(_06882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12850_ (.A1_N(_07496_),
    .A2_N(_07525_),
    .B1(\design_top.MEM[21][27] ),
    .B2(_07527_),
    .X(_06881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12851_ (.A1_N(_07497_),
    .A2_N(_07524_),
    .B1(\design_top.MEM[21][26] ),
    .B2(_07526_),
    .X(_06880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12852_ (.A1_N(_07498_),
    .A2_N(_07524_),
    .B1(\design_top.MEM[21][25] ),
    .B2(_07526_),
    .X(_06879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12853_ (.A1_N(_07499_),
    .A2_N(_07524_),
    .B1(\design_top.MEM[21][24] ),
    .B2(_07526_),
    .X(_06878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12854_ (.A(_11019_),
    .B(_11255_),
    .X(_07528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12855_ (.A(_07471_),
    .B(_07528_),
    .X(_07529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12856_ (.A(_07529_),
    .X(_07530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12857_ (.A(_07476_),
    .X(_07531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12858_ (.A1(_07435_),
    .A2(_07531_),
    .B1(_07529_),
    .X(_07532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12859_ (.A(_07532_),
    .X(_07533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12860_ (.A1_N(_07504_),
    .A2_N(_07530_),
    .B1(\design_top.MEM[22][15] ),
    .B2(_07533_),
    .X(_06877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12861_ (.A1_N(_07480_),
    .A2_N(_07530_),
    .B1(\design_top.MEM[22][14] ),
    .B2(_07533_),
    .X(_06876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12862_ (.A1_N(_07481_),
    .A2_N(_07530_),
    .B1(\design_top.MEM[22][13] ),
    .B2(_07533_),
    .X(_06875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12863_ (.A1_N(_07482_),
    .A2_N(_07530_),
    .B1(\design_top.MEM[22][12] ),
    .B2(_07533_),
    .X(_06874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12864_ (.A1_N(_07483_),
    .A2_N(_07530_),
    .B1(\design_top.MEM[22][11] ),
    .B2(_07533_),
    .X(_06873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12865_ (.A1_N(_07484_),
    .A2_N(_07529_),
    .B1(\design_top.MEM[22][10] ),
    .B2(_07532_),
    .X(_06872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12866_ (.A1_N(_07485_),
    .A2_N(_07529_),
    .B1(\design_top.MEM[22][9] ),
    .B2(_07532_),
    .X(_06871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12867_ (.A1_N(_07486_),
    .A2_N(_07529_),
    .B1(\design_top.MEM[22][8] ),
    .B2(_07532_),
    .X(_06870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12868_ (.A(_07448_),
    .B(_07528_),
    .X(_07534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12869_ (.A(_07534_),
    .X(_07535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12870_ (.A1(_07435_),
    .A2(_07531_),
    .B1(_07534_),
    .X(_07536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12871_ (.A(_07536_),
    .X(_07537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12872_ (.A1_N(_07447_),
    .A2_N(_07535_),
    .B1(\design_top.MEM[22][23] ),
    .B2(_07537_),
    .X(_06869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12873_ (.A1_N(_07459_),
    .A2_N(_07535_),
    .B1(\design_top.MEM[22][22] ),
    .B2(_07537_),
    .X(_06868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12874_ (.A1_N(_07460_),
    .A2_N(_07535_),
    .B1(\design_top.MEM[22][21] ),
    .B2(_07537_),
    .X(_06867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12875_ (.A1_N(_07461_),
    .A2_N(_07535_),
    .B1(\design_top.MEM[22][20] ),
    .B2(_07537_),
    .X(_06866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12876_ (.A1_N(_07462_),
    .A2_N(_07535_),
    .B1(\design_top.MEM[22][19] ),
    .B2(_07537_),
    .X(_06865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12877_ (.A1_N(_07463_),
    .A2_N(_07534_),
    .B1(\design_top.MEM[22][18] ),
    .B2(_07536_),
    .X(_06864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12878_ (.A1_N(_07464_),
    .A2_N(_07534_),
    .B1(\design_top.MEM[22][17] ),
    .B2(_07536_),
    .X(_06863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12879_ (.A1_N(_07465_),
    .A2_N(_07534_),
    .B1(\design_top.MEM[22][16] ),
    .B2(_07536_),
    .X(_06862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12880_ (.A(_11060_),
    .X(_07538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12881_ (.A(_11025_),
    .X(_07539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12882_ (.A(_07539_),
    .B(_07516_),
    .X(_07540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12883_ (.A(_07540_),
    .X(_07541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12884_ (.A(_11271_),
    .X(_07542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12885_ (.A1(_07542_),
    .A2(_07521_),
    .B1(_07540_),
    .X(_07543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12886_ (.A(_07543_),
    .X(_07544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12887_ (.A1_N(_07538_),
    .A2_N(_07541_),
    .B1(\design_top.MEM[36][23] ),
    .B2(_07544_),
    .X(_06861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12888_ (.A(_11066_),
    .X(_07545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12889_ (.A1_N(_07545_),
    .A2_N(_07541_),
    .B1(\design_top.MEM[36][22] ),
    .B2(_07544_),
    .X(_06860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12890_ (.A(_11068_),
    .X(_07546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12891_ (.A1_N(_07546_),
    .A2_N(_07541_),
    .B1(\design_top.MEM[36][21] ),
    .B2(_07544_),
    .X(_06859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12892_ (.A(_11070_),
    .X(_07547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12893_ (.A1_N(_07547_),
    .A2_N(_07541_),
    .B1(\design_top.MEM[36][20] ),
    .B2(_07544_),
    .X(_06858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12894_ (.A(_11072_),
    .X(_07548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12895_ (.A1_N(_07548_),
    .A2_N(_07541_),
    .B1(\design_top.MEM[36][19] ),
    .B2(_07544_),
    .X(_06857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12896_ (.A(_11074_),
    .X(_07549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12897_ (.A1_N(_07549_),
    .A2_N(_07540_),
    .B1(\design_top.MEM[36][18] ),
    .B2(_07543_),
    .X(_06856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12898_ (.A(_11076_),
    .X(_07550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12899_ (.A1_N(_07550_),
    .A2_N(_07540_),
    .B1(\design_top.MEM[36][17] ),
    .B2(_07543_),
    .X(_06855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12900_ (.A(_11078_),
    .X(_07551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12901_ (.A1_N(_07551_),
    .A2_N(_07540_),
    .B1(\design_top.MEM[36][16] ),
    .B2(_07543_),
    .X(_06854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12902_ (.A(_07488_),
    .B(_07516_),
    .X(_07552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12903_ (.A(_07552_),
    .X(_07553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12904_ (.A1(_07542_),
    .A2(_07521_),
    .B1(_07552_),
    .X(_07554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12905_ (.A(_07554_),
    .X(_07555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12906_ (.A1_N(_07487_),
    .A2_N(_07553_),
    .B1(\design_top.MEM[36][31] ),
    .B2(_07555_),
    .X(_06853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12907_ (.A1_N(_07493_),
    .A2_N(_07553_),
    .B1(\design_top.MEM[36][30] ),
    .B2(_07555_),
    .X(_06852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12908_ (.A1_N(_07494_),
    .A2_N(_07553_),
    .B1(\design_top.MEM[36][29] ),
    .B2(_07555_),
    .X(_06851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12909_ (.A1_N(_07495_),
    .A2_N(_07553_),
    .B1(\design_top.MEM[36][28] ),
    .B2(_07555_),
    .X(_06850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12910_ (.A1_N(_07496_),
    .A2_N(_07553_),
    .B1(\design_top.MEM[36][27] ),
    .B2(_07555_),
    .X(_06849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12911_ (.A1_N(_07497_),
    .A2_N(_07552_),
    .B1(\design_top.MEM[36][26] ),
    .B2(_07554_),
    .X(_06848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12912_ (.A1_N(_07498_),
    .A2_N(_07552_),
    .B1(\design_top.MEM[36][25] ),
    .B2(_07554_),
    .X(_06847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12913_ (.A1_N(_07499_),
    .A2_N(_07552_),
    .B1(\design_top.MEM[36][24] ),
    .B2(_07554_),
    .X(_06846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12914_ (.A(_02862_),
    .B(_02861_),
    .X(_07556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12915_ (.A(_03199_),
    .B(_07556_),
    .X(_07557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12916_ (.A(_07557_),
    .X(_07558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12917_ (.A(_10999_),
    .B(_07558_),
    .X(_07559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12918_ (.A(_07488_),
    .B(_07559_),
    .X(_07560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12919_ (.A(_07560_),
    .X(_07561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _12920_ (.A(_11110_),
    .B(_10894_),
    .C(wbs_adr_i[1]),
    .D(wbs_adr_i[0]),
    .X(_07562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12921_ (.A(_07562_),
    .X(_07563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12922_ (.A(_07563_),
    .X(_07564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12923_ (.A1(_07435_),
    .A2(_07564_),
    .B1(_07560_),
    .X(_07565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12924_ (.A(_07565_),
    .X(_07566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12925_ (.A1_N(_07487_),
    .A2_N(_07561_),
    .B1(\design_top.MEM[50][31] ),
    .B2(_07566_),
    .X(_06845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12926_ (.A1_N(_07493_),
    .A2_N(_07561_),
    .B1(\design_top.MEM[50][30] ),
    .B2(_07566_),
    .X(_06844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12927_ (.A1_N(_07494_),
    .A2_N(_07561_),
    .B1(\design_top.MEM[50][29] ),
    .B2(_07566_),
    .X(_06843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12928_ (.A1_N(_07495_),
    .A2_N(_07561_),
    .B1(\design_top.MEM[50][28] ),
    .B2(_07566_),
    .X(_06842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12929_ (.A1_N(_07496_),
    .A2_N(_07561_),
    .B1(\design_top.MEM[50][27] ),
    .B2(_07566_),
    .X(_06841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12930_ (.A1_N(_07497_),
    .A2_N(_07560_),
    .B1(\design_top.MEM[50][26] ),
    .B2(_07565_),
    .X(_06840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12931_ (.A1_N(_07498_),
    .A2_N(_07560_),
    .B1(\design_top.MEM[50][25] ),
    .B2(_07565_),
    .X(_06839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12932_ (.A1_N(_07499_),
    .A2_N(_07560_),
    .B1(\design_top.MEM[50][24] ),
    .B2(_07565_),
    .X(_06838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12933_ (.A(_11019_),
    .B(_07558_),
    .X(_07567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12934_ (.A(_07471_),
    .B(_07567_),
    .X(_07568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12935_ (.A(_07568_),
    .X(_07569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12936_ (.A(_07434_),
    .X(_07570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _12937_ (.A(_11110_),
    .B(_10893_),
    .C(wbs_adr_i[1]),
    .D(_10963_),
    .X(_07571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12938_ (.A(_07571_),
    .X(_07572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12939_ (.A(_07572_),
    .X(_07573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12940_ (.A1(_07570_),
    .A2(_07573_),
    .B1(_07568_),
    .X(_07574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12941_ (.A(_07574_),
    .X(_07575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12942_ (.A1_N(_07504_),
    .A2_N(_07569_),
    .B1(\design_top.MEM[54][15] ),
    .B2(_07575_),
    .X(_06837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12943_ (.A1_N(_07480_),
    .A2_N(_07569_),
    .B1(\design_top.MEM[54][14] ),
    .B2(_07575_),
    .X(_06836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12944_ (.A1_N(_07481_),
    .A2_N(_07569_),
    .B1(\design_top.MEM[54][13] ),
    .B2(_07575_),
    .X(_06835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12945_ (.A1_N(_07482_),
    .A2_N(_07569_),
    .B1(\design_top.MEM[54][12] ),
    .B2(_07575_),
    .X(_06834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12946_ (.A1_N(_07483_),
    .A2_N(_07569_),
    .B1(\design_top.MEM[54][11] ),
    .B2(_07575_),
    .X(_06833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12947_ (.A1_N(_07484_),
    .A2_N(_07568_),
    .B1(\design_top.MEM[54][10] ),
    .B2(_07574_),
    .X(_06832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12948_ (.A1_N(_07485_),
    .A2_N(_07568_),
    .B1(\design_top.MEM[54][9] ),
    .B2(_07574_),
    .X(_06831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12949_ (.A1_N(_07486_),
    .A2_N(_07568_),
    .B1(\design_top.MEM[54][8] ),
    .B2(_07574_),
    .X(_06830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12950_ (.A(_11037_),
    .X(_07576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12951_ (.A(_10884_),
    .B(_07558_),
    .X(_07577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12952_ (.A(_07576_),
    .B(_07577_),
    .X(_07578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12953_ (.A(_07578_),
    .X(_07579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12954_ (.A1(_07468_),
    .A2(_07564_),
    .B1(_07578_),
    .X(_07580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12955_ (.A(_07580_),
    .X(_07581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12956_ (.A1_N(_07504_),
    .A2_N(_07579_),
    .B1(\design_top.MEM[51][15] ),
    .B2(_07581_),
    .X(_06829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12957_ (.A(_11046_),
    .X(_07582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12958_ (.A1_N(_07582_),
    .A2_N(_07579_),
    .B1(\design_top.MEM[51][14] ),
    .B2(_07581_),
    .X(_06828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12959_ (.A(_11048_),
    .X(_07583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12960_ (.A1_N(_07583_),
    .A2_N(_07579_),
    .B1(\design_top.MEM[51][13] ),
    .B2(_07581_),
    .X(_06827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12961_ (.A(_11050_),
    .X(_07584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12962_ (.A1_N(_07584_),
    .A2_N(_07579_),
    .B1(\design_top.MEM[51][12] ),
    .B2(_07581_),
    .X(_06826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12963_ (.A(_11052_),
    .X(_07585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12964_ (.A1_N(_07585_),
    .A2_N(_07579_),
    .B1(\design_top.MEM[51][11] ),
    .B2(_07581_),
    .X(_06825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12965_ (.A(_11054_),
    .X(_07586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12966_ (.A1_N(_07586_),
    .A2_N(_07578_),
    .B1(\design_top.MEM[51][10] ),
    .B2(_07580_),
    .X(_06824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12967_ (.A(_11056_),
    .X(_07587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12968_ (.A1_N(_07587_),
    .A2_N(_07578_),
    .B1(\design_top.MEM[51][9] ),
    .B2(_07580_),
    .X(_06823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12969_ (.A(_11058_),
    .X(_07588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12970_ (.A1_N(_07588_),
    .A2_N(_07578_),
    .B1(\design_top.MEM[51][8] ),
    .B2(_07580_),
    .X(_06822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12971_ (.A(_07539_),
    .B(_07577_),
    .X(_07589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12972_ (.A(_07589_),
    .X(_07590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12973_ (.A1(_07468_),
    .A2(_07564_),
    .B1(_07589_),
    .X(_07591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12974_ (.A(_07591_),
    .X(_07592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12975_ (.A1_N(_07538_),
    .A2_N(_07590_),
    .B1(\design_top.MEM[51][23] ),
    .B2(_07592_),
    .X(_06821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12976_ (.A1_N(_07545_),
    .A2_N(_07590_),
    .B1(\design_top.MEM[51][22] ),
    .B2(_07592_),
    .X(_06820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12977_ (.A1_N(_07546_),
    .A2_N(_07590_),
    .B1(\design_top.MEM[51][21] ),
    .B2(_07592_),
    .X(_06819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12978_ (.A1_N(_07547_),
    .A2_N(_07590_),
    .B1(\design_top.MEM[51][20] ),
    .B2(_07592_),
    .X(_06818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12979_ (.A1_N(_07548_),
    .A2_N(_07590_),
    .B1(\design_top.MEM[51][19] ),
    .B2(_07592_),
    .X(_06817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12980_ (.A1_N(_07549_),
    .A2_N(_07589_),
    .B1(\design_top.MEM[51][18] ),
    .B2(_07591_),
    .X(_06816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12981_ (.A1_N(_07550_),
    .A2_N(_07589_),
    .B1(\design_top.MEM[51][17] ),
    .B2(_07591_),
    .X(_06815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12982_ (.A1_N(_07551_),
    .A2_N(_07589_),
    .B1(\design_top.MEM[51][16] ),
    .B2(_07591_),
    .X(_06814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12983_ (.A(_07488_),
    .B(_07577_),
    .X(_07593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12984_ (.A(_07593_),
    .X(_07594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12985_ (.A1(_07468_),
    .A2(_07564_),
    .B1(_07593_),
    .X(_07595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12986_ (.A(_07595_),
    .X(_07596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12987_ (.A1_N(_07487_),
    .A2_N(_07594_),
    .B1(\design_top.MEM[51][31] ),
    .B2(_07596_),
    .X(_06813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12988_ (.A1_N(_07493_),
    .A2_N(_07594_),
    .B1(\design_top.MEM[51][30] ),
    .B2(_07596_),
    .X(_06812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12989_ (.A1_N(_07494_),
    .A2_N(_07594_),
    .B1(\design_top.MEM[51][29] ),
    .B2(_07596_),
    .X(_06811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12990_ (.A1_N(_07495_),
    .A2_N(_07594_),
    .B1(\design_top.MEM[51][28] ),
    .B2(_07596_),
    .X(_06810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12991_ (.A1_N(_07496_),
    .A2_N(_07594_),
    .B1(\design_top.MEM[51][27] ),
    .B2(_07596_),
    .X(_06809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12992_ (.A1_N(_07497_),
    .A2_N(_07593_),
    .B1(\design_top.MEM[51][26] ),
    .B2(_07595_),
    .X(_06808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12993_ (.A1_N(_07498_),
    .A2_N(_07593_),
    .B1(\design_top.MEM[51][25] ),
    .B2(_07595_),
    .X(_06807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12994_ (.A1_N(_07499_),
    .A2_N(_07593_),
    .B1(\design_top.MEM[51][24] ),
    .B2(_07595_),
    .X(_06806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12995_ (.A(_07539_),
    .B(_07567_),
    .X(_07597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12996_ (.A(_07597_),
    .X(_07598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _12997_ (.A1(_07570_),
    .A2(_07573_),
    .B1(_07597_),
    .X(_07599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12998_ (.A(_07599_),
    .X(_07600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _12999_ (.A1_N(_07538_),
    .A2_N(_07598_),
    .B1(\design_top.MEM[54][23] ),
    .B2(_07600_),
    .X(_06805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13000_ (.A1_N(_07545_),
    .A2_N(_07598_),
    .B1(\design_top.MEM[54][22] ),
    .B2(_07600_),
    .X(_06804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13001_ (.A1_N(_07546_),
    .A2_N(_07598_),
    .B1(\design_top.MEM[54][21] ),
    .B2(_07600_),
    .X(_06803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13002_ (.A1_N(_07547_),
    .A2_N(_07598_),
    .B1(\design_top.MEM[54][20] ),
    .B2(_07600_),
    .X(_06802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13003_ (.A1_N(_07548_),
    .A2_N(_07598_),
    .B1(\design_top.MEM[54][19] ),
    .B2(_07600_),
    .X(_06801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13004_ (.A1_N(_07549_),
    .A2_N(_07597_),
    .B1(\design_top.MEM[54][18] ),
    .B2(_07599_),
    .X(_06800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13005_ (.A1_N(_07550_),
    .A2_N(_07597_),
    .B1(\design_top.MEM[54][17] ),
    .B2(_07599_),
    .X(_06799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13006_ (.A1_N(_07551_),
    .A2_N(_07597_),
    .B1(\design_top.MEM[54][16] ),
    .B2(_07599_),
    .X(_06798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13007_ (.A(_11100_),
    .X(_07601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13008_ (.A(_10957_),
    .B(_07558_),
    .X(_07602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13009_ (.A(_07576_),
    .B(_07602_),
    .X(_07603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13010_ (.A(_07603_),
    .X(_07604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13011_ (.A1(_07542_),
    .A2(_07573_),
    .B1(_07603_),
    .X(_07605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13012_ (.A(_07605_),
    .X(_07606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13013_ (.A1_N(_07601_),
    .A2_N(_07604_),
    .B1(\design_top.MEM[52][15] ),
    .B2(_07606_),
    .X(_06797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13014_ (.A1_N(_07582_),
    .A2_N(_07604_),
    .B1(\design_top.MEM[52][14] ),
    .B2(_07606_),
    .X(_06796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13015_ (.A1_N(_07583_),
    .A2_N(_07604_),
    .B1(\design_top.MEM[52][13] ),
    .B2(_07606_),
    .X(_06795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13016_ (.A1_N(_07584_),
    .A2_N(_07604_),
    .B1(\design_top.MEM[52][12] ),
    .B2(_07606_),
    .X(_06794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13017_ (.A1_N(_07585_),
    .A2_N(_07604_),
    .B1(\design_top.MEM[52][11] ),
    .B2(_07606_),
    .X(_06793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13018_ (.A1_N(_07586_),
    .A2_N(_07603_),
    .B1(\design_top.MEM[52][10] ),
    .B2(_07605_),
    .X(_06792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13019_ (.A1_N(_07587_),
    .A2_N(_07603_),
    .B1(\design_top.MEM[52][9] ),
    .B2(_07605_),
    .X(_06791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13020_ (.A1_N(_07588_),
    .A2_N(_07603_),
    .B1(\design_top.MEM[52][8] ),
    .B2(_07605_),
    .X(_06790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13021_ (.A(_11080_),
    .X(_07607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13022_ (.A(_11031_),
    .X(_07608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13023_ (.A(_07608_),
    .B(_07567_),
    .X(_07609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13024_ (.A(_07609_),
    .X(_07610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13025_ (.A1(_07570_),
    .A2(_07573_),
    .B1(_07609_),
    .X(_07611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13026_ (.A(_07611_),
    .X(_07612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13027_ (.A1_N(_07607_),
    .A2_N(_07610_),
    .B1(\design_top.MEM[54][31] ),
    .B2(_07612_),
    .X(_06789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13028_ (.A(_11086_),
    .X(_07613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13029_ (.A1_N(_07613_),
    .A2_N(_07610_),
    .B1(\design_top.MEM[54][30] ),
    .B2(_07612_),
    .X(_06788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13030_ (.A(_11088_),
    .X(_07614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13031_ (.A1_N(_07614_),
    .A2_N(_07610_),
    .B1(\design_top.MEM[54][29] ),
    .B2(_07612_),
    .X(_06787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13032_ (.A(_11090_),
    .X(_07615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13033_ (.A1_N(_07615_),
    .A2_N(_07610_),
    .B1(\design_top.MEM[54][28] ),
    .B2(_07612_),
    .X(_06786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13034_ (.A(_11092_),
    .X(_07616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13035_ (.A1_N(_07616_),
    .A2_N(_07610_),
    .B1(\design_top.MEM[54][27] ),
    .B2(_07612_),
    .X(_06785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13036_ (.A(_11094_),
    .X(_07617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13037_ (.A1_N(_07617_),
    .A2_N(_07609_),
    .B1(\design_top.MEM[54][26] ),
    .B2(_07611_),
    .X(_06784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13038_ (.A(_11096_),
    .X(_07618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13039_ (.A1_N(_07618_),
    .A2_N(_07609_),
    .B1(\design_top.MEM[54][25] ),
    .B2(_07611_),
    .X(_06783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13040_ (.A(_11098_),
    .X(_07619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13041_ (.A1_N(_07619_),
    .A2_N(_07609_),
    .B1(\design_top.MEM[54][24] ),
    .B2(_07611_),
    .X(_06782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13042_ (.A(_07539_),
    .B(_07602_),
    .X(_07620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13043_ (.A(_07620_),
    .X(_07621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13044_ (.A1(_07542_),
    .A2(_07573_),
    .B1(_07620_),
    .X(_07622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13045_ (.A(_07622_),
    .X(_07623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13046_ (.A1_N(_07538_),
    .A2_N(_07621_),
    .B1(\design_top.MEM[52][23] ),
    .B2(_07623_),
    .X(_06781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13047_ (.A1_N(_07545_),
    .A2_N(_07621_),
    .B1(\design_top.MEM[52][22] ),
    .B2(_07623_),
    .X(_06780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13048_ (.A1_N(_07546_),
    .A2_N(_07621_),
    .B1(\design_top.MEM[52][21] ),
    .B2(_07623_),
    .X(_06779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13049_ (.A1_N(_07547_),
    .A2_N(_07621_),
    .B1(\design_top.MEM[52][20] ),
    .B2(_07623_),
    .X(_06778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13050_ (.A1_N(_07548_),
    .A2_N(_07621_),
    .B1(\design_top.MEM[52][19] ),
    .B2(_07623_),
    .X(_06777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13051_ (.A1_N(_07549_),
    .A2_N(_07620_),
    .B1(\design_top.MEM[52][18] ),
    .B2(_07622_),
    .X(_06776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13052_ (.A1_N(_07550_),
    .A2_N(_07620_),
    .B1(\design_top.MEM[52][17] ),
    .B2(_07622_),
    .X(_06775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13053_ (.A1_N(_07551_),
    .A2_N(_07620_),
    .B1(\design_top.MEM[52][16] ),
    .B2(_07622_),
    .X(_06774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13054_ (.A(_11040_),
    .B(_07558_),
    .X(_07624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13055_ (.A(_07539_),
    .B(_07624_),
    .X(_07625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13056_ (.A(_07625_),
    .X(_07626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13057_ (.A(_11251_),
    .X(_07627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13058_ (.A(_07572_),
    .X(_07628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13059_ (.A1(_07627_),
    .A2(_07628_),
    .B1(_07625_),
    .X(_07629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13060_ (.A(_07629_),
    .X(_07630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13061_ (.A1_N(_07538_),
    .A2_N(_07626_),
    .B1(\design_top.MEM[55][23] ),
    .B2(_07630_),
    .X(_06773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13062_ (.A1_N(_07545_),
    .A2_N(_07626_),
    .B1(\design_top.MEM[55][22] ),
    .B2(_07630_),
    .X(_06772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13063_ (.A1_N(_07546_),
    .A2_N(_07626_),
    .B1(\design_top.MEM[55][21] ),
    .B2(_07630_),
    .X(_06771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13064_ (.A1_N(_07547_),
    .A2_N(_07626_),
    .B1(\design_top.MEM[55][20] ),
    .B2(_07630_),
    .X(_06770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13065_ (.A1_N(_07548_),
    .A2_N(_07626_),
    .B1(\design_top.MEM[55][19] ),
    .B2(_07630_),
    .X(_06769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13066_ (.A1_N(_07549_),
    .A2_N(_07625_),
    .B1(\design_top.MEM[55][18] ),
    .B2(_07629_),
    .X(_06768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13067_ (.A1_N(_07550_),
    .A2_N(_07625_),
    .B1(\design_top.MEM[55][17] ),
    .B2(_07629_),
    .X(_06767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13068_ (.A1_N(_07551_),
    .A2_N(_07625_),
    .B1(\design_top.MEM[55][16] ),
    .B2(_07629_),
    .X(_06766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13069_ (.A(_07608_),
    .B(_07624_),
    .X(_07631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13070_ (.A(_07631_),
    .X(_07632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13071_ (.A1(_07627_),
    .A2(_07628_),
    .B1(_07631_),
    .X(_07633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13072_ (.A(_07633_),
    .X(_07634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13073_ (.A1_N(_07607_),
    .A2_N(_07632_),
    .B1(\design_top.MEM[55][31] ),
    .B2(_07634_),
    .X(_06765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13074_ (.A1_N(_07613_),
    .A2_N(_07632_),
    .B1(\design_top.MEM[55][30] ),
    .B2(_07634_),
    .X(_06764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13075_ (.A1_N(_07614_),
    .A2_N(_07632_),
    .B1(\design_top.MEM[55][29] ),
    .B2(_07634_),
    .X(_06763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13076_ (.A1_N(_07615_),
    .A2_N(_07632_),
    .B1(\design_top.MEM[55][28] ),
    .B2(_07634_),
    .X(_06762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13077_ (.A1_N(_07616_),
    .A2_N(_07632_),
    .B1(\design_top.MEM[55][27] ),
    .B2(_07634_),
    .X(_06761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13078_ (.A1_N(_07617_),
    .A2_N(_07631_),
    .B1(\design_top.MEM[55][26] ),
    .B2(_07633_),
    .X(_06760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13079_ (.A1_N(_07618_),
    .A2_N(_07631_),
    .B1(\design_top.MEM[55][25] ),
    .B2(_07633_),
    .X(_06759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13080_ (.A1_N(_07619_),
    .A2_N(_07631_),
    .B1(\design_top.MEM[55][24] ),
    .B2(_07633_),
    .X(_06758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13081_ (.A(_07608_),
    .B(_07602_),
    .X(_07635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13082_ (.A(_07635_),
    .X(_07636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13083_ (.A1(_07542_),
    .A2(_07628_),
    .B1(_07635_),
    .X(_07637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13084_ (.A(_07637_),
    .X(_07638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13085_ (.A1_N(_07607_),
    .A2_N(_07636_),
    .B1(\design_top.MEM[52][31] ),
    .B2(_07638_),
    .X(_06757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13086_ (.A1_N(_07613_),
    .A2_N(_07636_),
    .B1(\design_top.MEM[52][30] ),
    .B2(_07638_),
    .X(_06756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13087_ (.A1_N(_07614_),
    .A2_N(_07636_),
    .B1(\design_top.MEM[52][29] ),
    .B2(_07638_),
    .X(_06755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13088_ (.A1_N(_07615_),
    .A2_N(_07636_),
    .B1(\design_top.MEM[52][28] ),
    .B2(_07638_),
    .X(_06754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13089_ (.A1_N(_07616_),
    .A2_N(_07636_),
    .B1(\design_top.MEM[52][27] ),
    .B2(_07638_),
    .X(_06753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13090_ (.A1_N(_07617_),
    .A2_N(_07635_),
    .B1(\design_top.MEM[52][26] ),
    .B2(_07637_),
    .X(_06752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13091_ (.A1_N(_07618_),
    .A2_N(_07635_),
    .B1(\design_top.MEM[52][25] ),
    .B2(_07637_),
    .X(_06751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13092_ (.A1_N(_07619_),
    .A2_N(_07635_),
    .B1(\design_top.MEM[52][24] ),
    .B2(_07637_),
    .X(_06750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13093_ (.A(_10874_),
    .X(_07639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13094_ (.A(_07639_),
    .X(_07640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13095_ (.A(_10877_),
    .X(_07641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13096_ (.A(_07641_),
    .X(_07642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13097_ (.A(_10979_),
    .B(_07557_),
    .X(_07643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13098_ (.A(_07642_),
    .B(_07643_),
    .X(_07644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13099_ (.A(_07644_),
    .X(_07645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13100_ (.A1(_07509_),
    .A2(_07628_),
    .B1(_07644_),
    .X(_07646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13101_ (.A(_07646_),
    .X(_07647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13102_ (.A1_N(_07640_),
    .A2_N(_07645_),
    .B1(\design_top.MEM[53][23] ),
    .B2(_07647_),
    .X(_06749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13103_ (.A(_10902_),
    .X(_07648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13104_ (.A(_07648_),
    .X(_07649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13105_ (.A1_N(_07649_),
    .A2_N(_07645_),
    .B1(\design_top.MEM[53][22] ),
    .B2(_07647_),
    .X(_06748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13106_ (.A(_10905_),
    .X(_07650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13107_ (.A(_07650_),
    .X(_07651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13108_ (.A1_N(_07651_),
    .A2_N(_07645_),
    .B1(\design_top.MEM[53][21] ),
    .B2(_07647_),
    .X(_06747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13109_ (.A(_10908_),
    .X(_07652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13110_ (.A(_07652_),
    .X(_07653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13111_ (.A1_N(_07653_),
    .A2_N(_07645_),
    .B1(\design_top.MEM[53][20] ),
    .B2(_07647_),
    .X(_06746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13112_ (.A(_10911_),
    .X(_07654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13113_ (.A(_07654_),
    .X(_07655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13114_ (.A1_N(_07655_),
    .A2_N(_07645_),
    .B1(\design_top.MEM[53][19] ),
    .B2(_07647_),
    .X(_06745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13115_ (.A(_10914_),
    .X(_07656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13116_ (.A(_07656_),
    .X(_07657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13117_ (.A1_N(_07657_),
    .A2_N(_07644_),
    .B1(\design_top.MEM[53][18] ),
    .B2(_07646_),
    .X(_06744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13118_ (.A(_10917_),
    .X(_07658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13119_ (.A(_07658_),
    .X(_07659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13120_ (.A1_N(_07659_),
    .A2_N(_07644_),
    .B1(\design_top.MEM[53][17] ),
    .B2(_07646_),
    .X(_06743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13121_ (.A(_10920_),
    .X(_07660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13122_ (.A(_07660_),
    .X(_07661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13123_ (.A1_N(_07661_),
    .A2_N(_07644_),
    .B1(\design_top.MEM[53][16] ),
    .B2(_07646_),
    .X(_06742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13124_ (.A(_07608_),
    .B(_07643_),
    .X(_07662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13125_ (.A(_07662_),
    .X(_07663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13126_ (.A1(_07509_),
    .A2(_07628_),
    .B1(_07662_),
    .X(_07664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13127_ (.A(_07664_),
    .X(_07665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13128_ (.A1_N(_07607_),
    .A2_N(_07663_),
    .B1(\design_top.MEM[53][31] ),
    .B2(_07665_),
    .X(_06741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13129_ (.A1_N(_07613_),
    .A2_N(_07663_),
    .B1(\design_top.MEM[53][30] ),
    .B2(_07665_),
    .X(_06740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13130_ (.A1_N(_07614_),
    .A2_N(_07663_),
    .B1(\design_top.MEM[53][29] ),
    .B2(_07665_),
    .X(_06739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13131_ (.A1_N(_07615_),
    .A2_N(_07663_),
    .B1(\design_top.MEM[53][28] ),
    .B2(_07665_),
    .X(_06738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13132_ (.A1_N(_07616_),
    .A2_N(_07663_),
    .B1(\design_top.MEM[53][27] ),
    .B2(_07665_),
    .X(_06737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13133_ (.A1_N(_07617_),
    .A2_N(_07662_),
    .B1(\design_top.MEM[53][26] ),
    .B2(_07664_),
    .X(_06736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13134_ (.A1_N(_07618_),
    .A2_N(_07662_),
    .B1(\design_top.MEM[53][25] ),
    .B2(_07664_),
    .X(_06735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13135_ (.A1_N(_07619_),
    .A2_N(_07662_),
    .B1(\design_top.MEM[53][24] ),
    .B2(_07664_),
    .X(_06734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13136_ (.A(_07576_),
    .B(_07643_),
    .X(_07666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13137_ (.A(_07666_),
    .X(_07667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13138_ (.A(_07508_),
    .X(_07668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13139_ (.A1(_07668_),
    .A2(_07572_),
    .B1(_07666_),
    .X(_07669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13140_ (.A(_07669_),
    .X(_07670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13141_ (.A1_N(_07601_),
    .A2_N(_07667_),
    .B1(\design_top.MEM[53][15] ),
    .B2(_07670_),
    .X(_06733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13142_ (.A1_N(_07582_),
    .A2_N(_07667_),
    .B1(\design_top.MEM[53][14] ),
    .B2(_07670_),
    .X(_06732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13143_ (.A1_N(_07583_),
    .A2_N(_07667_),
    .B1(\design_top.MEM[53][13] ),
    .B2(_07670_),
    .X(_06731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13144_ (.A1_N(_07584_),
    .A2_N(_07667_),
    .B1(\design_top.MEM[53][12] ),
    .B2(_07670_),
    .X(_06730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13145_ (.A1_N(_07585_),
    .A2_N(_07667_),
    .B1(\design_top.MEM[53][11] ),
    .B2(_07670_),
    .X(_06729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13146_ (.A1_N(_07586_),
    .A2_N(_07666_),
    .B1(\design_top.MEM[53][10] ),
    .B2(_07669_),
    .X(_06728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13147_ (.A1_N(_07587_),
    .A2_N(_07666_),
    .B1(\design_top.MEM[53][9] ),
    .B2(_07669_),
    .X(_06727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13148_ (.A1_N(_07588_),
    .A2_N(_07666_),
    .B1(\design_top.MEM[53][8] ),
    .B2(_07669_),
    .X(_06726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13149_ (.A(_11018_),
    .B(_11105_),
    .X(_07671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13150_ (.A(_07608_),
    .B(_07671_),
    .X(_07672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13151_ (.A(_07672_),
    .X(_07673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13152_ (.A1(_07570_),
    .A2(_07521_),
    .B1(_07672_),
    .X(_07674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13153_ (.A(_07674_),
    .X(_07675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13154_ (.A1_N(_07607_),
    .A2_N(_07673_),
    .B1(\design_top.MEM[38][31] ),
    .B2(_07675_),
    .X(_06725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13155_ (.A1_N(_07613_),
    .A2_N(_07673_),
    .B1(\design_top.MEM[38][30] ),
    .B2(_07675_),
    .X(_06724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13156_ (.A1_N(_07614_),
    .A2_N(_07673_),
    .B1(\design_top.MEM[38][29] ),
    .B2(_07675_),
    .X(_06723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13157_ (.A1_N(_07615_),
    .A2_N(_07673_),
    .B1(\design_top.MEM[38][28] ),
    .B2(_07675_),
    .X(_06722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13158_ (.A1_N(_07616_),
    .A2_N(_07673_),
    .B1(\design_top.MEM[38][27] ),
    .B2(_07675_),
    .X(_06721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13159_ (.A1_N(_07617_),
    .A2_N(_07672_),
    .B1(\design_top.MEM[38][26] ),
    .B2(_07674_),
    .X(_06720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13160_ (.A1_N(_07618_),
    .A2_N(_07672_),
    .B1(\design_top.MEM[38][25] ),
    .B2(_07674_),
    .X(_06719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13161_ (.A1_N(_07619_),
    .A2_N(_07672_),
    .B1(\design_top.MEM[38][24] ),
    .B2(_07674_),
    .X(_06718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13162_ (.A(_10820_),
    .X(_07676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13163_ (.A(_07676_),
    .X(_07677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13164_ (.A(_10925_),
    .X(_07678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13165_ (.A(_07678_),
    .X(_07679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13166_ (.A(_07679_),
    .B(_07451_),
    .X(_07680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13167_ (.A(_07680_),
    .X(_07681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13168_ (.A1(_07668_),
    .A2(_07456_),
    .B1(_07680_),
    .X(_07682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13169_ (.A(_07682_),
    .X(_07683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13170_ (.A1_N(_07677_),
    .A2_N(_07681_),
    .B1(\design_top.MEM[45][31] ),
    .B2(_07683_),
    .X(_06717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13171_ (.A(_10932_),
    .X(_07684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13172_ (.A(_07684_),
    .X(_07685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13173_ (.A1_N(_07685_),
    .A2_N(_07681_),
    .B1(\design_top.MEM[45][30] ),
    .B2(_07683_),
    .X(_06716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13174_ (.A(_10935_),
    .X(_07686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13175_ (.A(_07686_),
    .X(_07687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13176_ (.A1_N(_07687_),
    .A2_N(_07681_),
    .B1(\design_top.MEM[45][29] ),
    .B2(_07683_),
    .X(_06715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13177_ (.A(_10938_),
    .X(_07688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13178_ (.A(_07688_),
    .X(_07689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13179_ (.A1_N(_07689_),
    .A2_N(_07681_),
    .B1(\design_top.MEM[45][28] ),
    .B2(_07683_),
    .X(_06714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13180_ (.A(_10941_),
    .X(_07690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13181_ (.A(_07690_),
    .X(_07691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13182_ (.A1_N(_07691_),
    .A2_N(_07681_),
    .B1(\design_top.MEM[45][27] ),
    .B2(_07683_),
    .X(_06713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13183_ (.A(_10944_),
    .X(_07692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13184_ (.A(_07692_),
    .X(_07693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13185_ (.A1_N(_07693_),
    .A2_N(_07680_),
    .B1(\design_top.MEM[45][26] ),
    .B2(_07682_),
    .X(_06712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13186_ (.A(_10947_),
    .X(_07694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13187_ (.A(_07694_),
    .X(_07695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13188_ (.A1_N(_07695_),
    .A2_N(_07680_),
    .B1(\design_top.MEM[45][25] ),
    .B2(_07682_),
    .X(_06711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13189_ (.A(_10950_),
    .X(_07696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13190_ (.A(_07696_),
    .X(_07697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13191_ (.A1_N(_07697_),
    .A2_N(_07680_),
    .B1(\design_top.MEM[45][24] ),
    .B2(_07682_),
    .X(_06710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13192_ (.A(_11040_),
    .B(_11104_),
    .X(_07698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13193_ (.A(_07576_),
    .B(_07698_),
    .X(_07699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13194_ (.A(_07699_),
    .X(_07700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13195_ (.A1(_07627_),
    .A2(_07521_),
    .B1(_07699_),
    .X(_07701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13196_ (.A(_07701_),
    .X(_07702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13197_ (.A1_N(_07601_),
    .A2_N(_07700_),
    .B1(\design_top.MEM[39][15] ),
    .B2(_07702_),
    .X(_06709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13198_ (.A1_N(_07582_),
    .A2_N(_07700_),
    .B1(\design_top.MEM[39][14] ),
    .B2(_07702_),
    .X(_06708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13199_ (.A1_N(_07583_),
    .A2_N(_07700_),
    .B1(\design_top.MEM[39][13] ),
    .B2(_07702_),
    .X(_06707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13200_ (.A1_N(_07584_),
    .A2_N(_07700_),
    .B1(\design_top.MEM[39][12] ),
    .B2(_07702_),
    .X(_06706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13201_ (.A1_N(_07585_),
    .A2_N(_07700_),
    .B1(\design_top.MEM[39][11] ),
    .B2(_07702_),
    .X(_06705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13202_ (.A1_N(_07586_),
    .A2_N(_07699_),
    .B1(\design_top.MEM[39][10] ),
    .B2(_07701_),
    .X(_06704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13203_ (.A1_N(_07587_),
    .A2_N(_07699_),
    .B1(\design_top.MEM[39][9] ),
    .B2(_07701_),
    .X(_06703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13204_ (.A1_N(_07588_),
    .A2_N(_07699_),
    .B1(\design_top.MEM[39][8] ),
    .B2(_07701_),
    .X(_06702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13205_ (.A(_11018_),
    .B(_07450_),
    .X(_07703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13206_ (.A(_07576_),
    .B(_07703_),
    .X(_07704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13207_ (.A(_07704_),
    .X(_07705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13208_ (.A1(_07570_),
    .A2(_07456_),
    .B1(_07704_),
    .X(_07706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13209_ (.A(_07706_),
    .X(_07707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13210_ (.A1_N(_07601_),
    .A2_N(_07705_),
    .B1(\design_top.MEM[46][15] ),
    .B2(_07707_),
    .X(_06701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13211_ (.A1_N(_07582_),
    .A2_N(_07705_),
    .B1(\design_top.MEM[46][14] ),
    .B2(_07707_),
    .X(_06700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13212_ (.A1_N(_07583_),
    .A2_N(_07705_),
    .B1(\design_top.MEM[46][13] ),
    .B2(_07707_),
    .X(_06699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13213_ (.A1_N(_07584_),
    .A2_N(_07705_),
    .B1(\design_top.MEM[46][12] ),
    .B2(_07707_),
    .X(_06698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13214_ (.A1_N(_07585_),
    .A2_N(_07705_),
    .B1(\design_top.MEM[46][11] ),
    .B2(_07707_),
    .X(_06697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13215_ (.A1_N(_07586_),
    .A2_N(_07704_),
    .B1(\design_top.MEM[46][10] ),
    .B2(_07706_),
    .X(_06696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13216_ (.A1_N(_07587_),
    .A2_N(_07704_),
    .B1(\design_top.MEM[46][9] ),
    .B2(_07706_),
    .X(_06695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13217_ (.A1_N(_07588_),
    .A2_N(_07704_),
    .B1(\design_top.MEM[46][8] ),
    .B2(_07706_),
    .X(_06694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13218_ (.A(_07642_),
    .B(_07698_),
    .X(_07708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13219_ (.A(_07708_),
    .X(_07709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13220_ (.A(_07520_),
    .X(_07710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13221_ (.A1(_07627_),
    .A2(_07710_),
    .B1(_07708_),
    .X(_07711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13222_ (.A(_07711_),
    .X(_07712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13223_ (.A1_N(_07640_),
    .A2_N(_07709_),
    .B1(\design_top.MEM[39][23] ),
    .B2(_07712_),
    .X(_06693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13224_ (.A1_N(_07649_),
    .A2_N(_07709_),
    .B1(\design_top.MEM[39][22] ),
    .B2(_07712_),
    .X(_06692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13225_ (.A1_N(_07651_),
    .A2_N(_07709_),
    .B1(\design_top.MEM[39][21] ),
    .B2(_07712_),
    .X(_06691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13226_ (.A1_N(_07653_),
    .A2_N(_07709_),
    .B1(\design_top.MEM[39][20] ),
    .B2(_07712_),
    .X(_06690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13227_ (.A1_N(_07655_),
    .A2_N(_07709_),
    .B1(\design_top.MEM[39][19] ),
    .B2(_07712_),
    .X(_06689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13228_ (.A1_N(_07657_),
    .A2_N(_07708_),
    .B1(\design_top.MEM[39][18] ),
    .B2(_07711_),
    .X(_06688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13229_ (.A1_N(_07659_),
    .A2_N(_07708_),
    .B1(\design_top.MEM[39][17] ),
    .B2(_07711_),
    .X(_06687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13230_ (.A1_N(_07661_),
    .A2_N(_07708_),
    .B1(\design_top.MEM[39][16] ),
    .B2(_07711_),
    .X(_06686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13231_ (.A(_07642_),
    .B(_07703_),
    .X(_07713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13232_ (.A(_07713_),
    .X(_07714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13233_ (.A(_07434_),
    .X(_07715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13234_ (.A1(_07715_),
    .A2(_07456_),
    .B1(_07713_),
    .X(_07716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13235_ (.A(_07716_),
    .X(_07717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13236_ (.A1_N(_07640_),
    .A2_N(_07714_),
    .B1(\design_top.MEM[46][23] ),
    .B2(_07717_),
    .X(_06685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13237_ (.A1_N(_07649_),
    .A2_N(_07714_),
    .B1(\design_top.MEM[46][22] ),
    .B2(_07717_),
    .X(_06684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13238_ (.A1_N(_07651_),
    .A2_N(_07714_),
    .B1(\design_top.MEM[46][21] ),
    .B2(_07717_),
    .X(_06683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13239_ (.A1_N(_07653_),
    .A2_N(_07714_),
    .B1(\design_top.MEM[46][20] ),
    .B2(_07717_),
    .X(_06682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13240_ (.A1_N(_07655_),
    .A2_N(_07714_),
    .B1(\design_top.MEM[46][19] ),
    .B2(_07717_),
    .X(_06681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13241_ (.A1_N(_07657_),
    .A2_N(_07713_),
    .B1(\design_top.MEM[46][18] ),
    .B2(_07716_),
    .X(_06680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13242_ (.A1_N(_07659_),
    .A2_N(_07713_),
    .B1(\design_top.MEM[46][17] ),
    .B2(_07716_),
    .X(_06679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13243_ (.A1_N(_07661_),
    .A2_N(_07713_),
    .B1(\design_top.MEM[46][16] ),
    .B2(_07716_),
    .X(_06678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13244_ (.A(_07679_),
    .B(_07703_),
    .X(_07718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13245_ (.A(_07718_),
    .X(_07719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13246_ (.A1(_07715_),
    .A2(_07456_),
    .B1(_07718_),
    .X(_07720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13247_ (.A(_07720_),
    .X(_07721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13248_ (.A1_N(_07677_),
    .A2_N(_07719_),
    .B1(\design_top.MEM[46][31] ),
    .B2(_07721_),
    .X(_06677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13249_ (.A1_N(_07685_),
    .A2_N(_07719_),
    .B1(\design_top.MEM[46][30] ),
    .B2(_07721_),
    .X(_06676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13250_ (.A1_N(_07687_),
    .A2_N(_07719_),
    .B1(\design_top.MEM[46][29] ),
    .B2(_07721_),
    .X(_06675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13251_ (.A1_N(_07689_),
    .A2_N(_07719_),
    .B1(\design_top.MEM[46][28] ),
    .B2(_07721_),
    .X(_06674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13252_ (.A1_N(_07691_),
    .A2_N(_07719_),
    .B1(\design_top.MEM[46][27] ),
    .B2(_07721_),
    .X(_06673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13253_ (.A1_N(_07693_),
    .A2_N(_07718_),
    .B1(\design_top.MEM[46][26] ),
    .B2(_07720_),
    .X(_06672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13254_ (.A1_N(_07695_),
    .A2_N(_07718_),
    .B1(\design_top.MEM[46][25] ),
    .B2(_07720_),
    .X(_06671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13255_ (.A1_N(_07697_),
    .A2_N(_07718_),
    .B1(\design_top.MEM[46][24] ),
    .B2(_07720_),
    .X(_06670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13256_ (.A(_07679_),
    .B(_07698_),
    .X(_07722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13257_ (.A(_07722_),
    .X(_07723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13258_ (.A1(_07627_),
    .A2(_07710_),
    .B1(_07722_),
    .X(_07724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13259_ (.A(_07724_),
    .X(_07725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13260_ (.A1_N(_07677_),
    .A2_N(_07723_),
    .B1(\design_top.MEM[39][31] ),
    .B2(_07725_),
    .X(_06669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13261_ (.A1_N(_07685_),
    .A2_N(_07723_),
    .B1(\design_top.MEM[39][30] ),
    .B2(_07725_),
    .X(_06668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13262_ (.A1_N(_07687_),
    .A2_N(_07723_),
    .B1(\design_top.MEM[39][29] ),
    .B2(_07725_),
    .X(_06667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13263_ (.A1_N(_07689_),
    .A2_N(_07723_),
    .B1(\design_top.MEM[39][28] ),
    .B2(_07725_),
    .X(_06666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13264_ (.A1_N(_07691_),
    .A2_N(_07723_),
    .B1(\design_top.MEM[39][27] ),
    .B2(_07725_),
    .X(_06665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13265_ (.A1_N(_07693_),
    .A2_N(_07722_),
    .B1(\design_top.MEM[39][26] ),
    .B2(_07724_),
    .X(_06664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13266_ (.A1_N(_07695_),
    .A2_N(_07722_),
    .B1(\design_top.MEM[39][25] ),
    .B2(_07724_),
    .X(_06663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13267_ (.A1_N(_07697_),
    .A2_N(_07722_),
    .B1(\design_top.MEM[39][24] ),
    .B2(_07724_),
    .X(_06662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13268_ (.A(_10767_),
    .X(_07726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13269_ (.A(_07726_),
    .X(_07727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13270_ (.A(_11039_),
    .B(_07450_),
    .X(_07728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13271_ (.A(_07727_),
    .B(_07728_),
    .X(_07729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13272_ (.A(_07729_),
    .X(_07730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13273_ (.A(_11251_),
    .X(_07731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13274_ (.A(_07455_),
    .X(_07732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13275_ (.A1(_07731_),
    .A2(_07732_),
    .B1(_07729_),
    .X(_07733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13276_ (.A(_07733_),
    .X(_07734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13277_ (.A1_N(_07601_),
    .A2_N(_07730_),
    .B1(\design_top.MEM[47][15] ),
    .B2(_07734_),
    .X(_06661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13278_ (.A(_10587_),
    .X(_07735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13279_ (.A(_07735_),
    .X(_07736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13280_ (.A1_N(_07736_),
    .A2_N(_07730_),
    .B1(\design_top.MEM[47][14] ),
    .B2(_07734_),
    .X(_06660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13281_ (.A(_10802_),
    .X(_07737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13282_ (.A(_07737_),
    .X(_07738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13283_ (.A1_N(_07738_),
    .A2_N(_07730_),
    .B1(\design_top.MEM[47][13] ),
    .B2(_07734_),
    .X(_06659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13284_ (.A(_10805_),
    .X(_07739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13285_ (.A(_07739_),
    .X(_07740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13286_ (.A1_N(_07740_),
    .A2_N(_07730_),
    .B1(\design_top.MEM[47][12] ),
    .B2(_07734_),
    .X(_06658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13287_ (.A(_10808_),
    .X(_07741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13288_ (.A(_07741_),
    .X(_07742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13289_ (.A1_N(_07742_),
    .A2_N(_07730_),
    .B1(\design_top.MEM[47][11] ),
    .B2(_07734_),
    .X(_06657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13290_ (.A(_10811_),
    .X(_07743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13291_ (.A(_07743_),
    .X(_07744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13292_ (.A1_N(_07744_),
    .A2_N(_07729_),
    .B1(\design_top.MEM[47][10] ),
    .B2(_07733_),
    .X(_06656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13293_ (.A(_10814_),
    .X(_07745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13294_ (.A(_07745_),
    .X(_07746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13295_ (.A1_N(_07746_),
    .A2_N(_07729_),
    .B1(\design_top.MEM[47][9] ),
    .B2(_07733_),
    .X(_06655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13296_ (.A(_10817_),
    .X(_07747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13297_ (.A(_07747_),
    .X(_07748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13298_ (.A1_N(_07748_),
    .A2_N(_07729_),
    .B1(\design_top.MEM[47][8] ),
    .B2(_07733_),
    .X(_06654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13299_ (.A(_10953_),
    .X(_07749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13300_ (.A(_07749_),
    .X(_07750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13301_ (.A(_10783_),
    .B(_10885_),
    .X(_07751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13302_ (.A(_07727_),
    .B(_07751_),
    .X(_07752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13303_ (.A(_07752_),
    .X(_07753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13304_ (.A1(_11126_),
    .A2(_10891_),
    .B1(_07752_),
    .X(_07754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13305_ (.A(_07754_),
    .X(_07755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13306_ (.A1_N(_07750_),
    .A2_N(_07753_),
    .B1(\design_top.MEM[3][15] ),
    .B2(_07755_),
    .X(_06653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13307_ (.A1_N(_07736_),
    .A2_N(_07753_),
    .B1(\design_top.MEM[3][14] ),
    .B2(_07755_),
    .X(_06652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13308_ (.A1_N(_07738_),
    .A2_N(_07753_),
    .B1(\design_top.MEM[3][13] ),
    .B2(_07755_),
    .X(_06651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13309_ (.A1_N(_07740_),
    .A2_N(_07753_),
    .B1(\design_top.MEM[3][12] ),
    .B2(_07755_),
    .X(_06650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13310_ (.A1_N(_07742_),
    .A2_N(_07753_),
    .B1(\design_top.MEM[3][11] ),
    .B2(_07755_),
    .X(_06649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13311_ (.A1_N(_07744_),
    .A2_N(_07752_),
    .B1(\design_top.MEM[3][10] ),
    .B2(_07754_),
    .X(_06648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13312_ (.A1_N(_07746_),
    .A2_N(_07752_),
    .B1(\design_top.MEM[3][9] ),
    .B2(_07754_),
    .X(_06647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13313_ (.A1_N(_07748_),
    .A2_N(_07752_),
    .B1(\design_top.MEM[3][8] ),
    .B2(_07754_),
    .X(_06646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13314_ (.A(_07642_),
    .B(_07751_),
    .X(_07756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13315_ (.A(_07756_),
    .X(_07757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13316_ (.A1(_11126_),
    .A2(_10891_),
    .B1(_07756_),
    .X(_07758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13317_ (.A(_07758_),
    .X(_07759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13318_ (.A1_N(_07640_),
    .A2_N(_07757_),
    .B1(\design_top.MEM[3][23] ),
    .B2(_07759_),
    .X(_06645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13319_ (.A1_N(_07649_),
    .A2_N(_07757_),
    .B1(\design_top.MEM[3][22] ),
    .B2(_07759_),
    .X(_06644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13320_ (.A1_N(_07651_),
    .A2_N(_07757_),
    .B1(\design_top.MEM[3][21] ),
    .B2(_07759_),
    .X(_06643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13321_ (.A1_N(_07653_),
    .A2_N(_07757_),
    .B1(\design_top.MEM[3][20] ),
    .B2(_07759_),
    .X(_06642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13322_ (.A1_N(_07655_),
    .A2_N(_07757_),
    .B1(\design_top.MEM[3][19] ),
    .B2(_07759_),
    .X(_06641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13323_ (.A1_N(_07657_),
    .A2_N(_07756_),
    .B1(\design_top.MEM[3][18] ),
    .B2(_07758_),
    .X(_06640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13324_ (.A1_N(_07659_),
    .A2_N(_07756_),
    .B1(\design_top.MEM[3][17] ),
    .B2(_07758_),
    .X(_06639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13325_ (.A1_N(_07661_),
    .A2_N(_07756_),
    .B1(\design_top.MEM[3][16] ),
    .B2(_07758_),
    .X(_06638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13326_ (.A(_07679_),
    .B(_07751_),
    .X(_07760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13327_ (.A(_07760_),
    .X(_07761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13328_ (.A1(_11126_),
    .A2(_10891_),
    .B1(_07760_),
    .X(_07762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13329_ (.A(_07762_),
    .X(_07763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13330_ (.A1_N(_07677_),
    .A2_N(_07761_),
    .B1(\design_top.MEM[3][31] ),
    .B2(_07763_),
    .X(_06637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13331_ (.A1_N(_07685_),
    .A2_N(_07761_),
    .B1(\design_top.MEM[3][30] ),
    .B2(_07763_),
    .X(_06636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13332_ (.A1_N(_07687_),
    .A2_N(_07761_),
    .B1(\design_top.MEM[3][29] ),
    .B2(_07763_),
    .X(_06635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13333_ (.A1_N(_07689_),
    .A2_N(_07761_),
    .B1(\design_top.MEM[3][28] ),
    .B2(_07763_),
    .X(_06634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13334_ (.A1_N(_07691_),
    .A2_N(_07761_),
    .B1(\design_top.MEM[3][27] ),
    .B2(_07763_),
    .X(_06633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13335_ (.A1_N(_07693_),
    .A2_N(_07760_),
    .B1(\design_top.MEM[3][26] ),
    .B2(_07762_),
    .X(_06632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13336_ (.A1_N(_07695_),
    .A2_N(_07760_),
    .B1(\design_top.MEM[3][25] ),
    .B2(_07762_),
    .X(_06631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13337_ (.A1_N(_07697_),
    .A2_N(_07760_),
    .B1(\design_top.MEM[3][24] ),
    .B2(_07762_),
    .X(_06630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13338_ (.A(_07642_),
    .B(_07728_),
    .X(_07764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13339_ (.A(_07764_),
    .X(_07765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13340_ (.A1(_07731_),
    .A2(_07732_),
    .B1(_07764_),
    .X(_07766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13341_ (.A(_07766_),
    .X(_07767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13342_ (.A1_N(_07640_),
    .A2_N(_07765_),
    .B1(\design_top.MEM[47][23] ),
    .B2(_07767_),
    .X(_06629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13343_ (.A1_N(_07649_),
    .A2_N(_07765_),
    .B1(\design_top.MEM[47][22] ),
    .B2(_07767_),
    .X(_06628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13344_ (.A1_N(_07651_),
    .A2_N(_07765_),
    .B1(\design_top.MEM[47][21] ),
    .B2(_07767_),
    .X(_06627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13345_ (.A1_N(_07653_),
    .A2_N(_07765_),
    .B1(\design_top.MEM[47][20] ),
    .B2(_07767_),
    .X(_06626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13346_ (.A1_N(_07655_),
    .A2_N(_07765_),
    .B1(\design_top.MEM[47][19] ),
    .B2(_07767_),
    .X(_06625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13347_ (.A1_N(_07657_),
    .A2_N(_07764_),
    .B1(\design_top.MEM[47][18] ),
    .B2(_07766_),
    .X(_06624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13348_ (.A1_N(_07659_),
    .A2_N(_07764_),
    .B1(\design_top.MEM[47][17] ),
    .B2(_07766_),
    .X(_06623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13349_ (.A1_N(_07661_),
    .A2_N(_07764_),
    .B1(\design_top.MEM[47][16] ),
    .B2(_07766_),
    .X(_06622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13350_ (.A(_07679_),
    .B(_07728_),
    .X(_07768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13351_ (.A(_07768_),
    .X(_07769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13352_ (.A1(_07731_),
    .A2(_07732_),
    .B1(_07768_),
    .X(_07770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13353_ (.A(_07770_),
    .X(_07771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13354_ (.A1_N(_07677_),
    .A2_N(_07769_),
    .B1(\design_top.MEM[47][31] ),
    .B2(_07771_),
    .X(_06621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13355_ (.A1_N(_07685_),
    .A2_N(_07769_),
    .B1(\design_top.MEM[47][30] ),
    .B2(_07771_),
    .X(_06620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13356_ (.A1_N(_07687_),
    .A2_N(_07769_),
    .B1(\design_top.MEM[47][29] ),
    .B2(_07771_),
    .X(_06619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13357_ (.A1_N(_07689_),
    .A2_N(_07769_),
    .B1(\design_top.MEM[47][28] ),
    .B2(_07771_),
    .X(_06618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13358_ (.A1_N(_07691_),
    .A2_N(_07769_),
    .B1(\design_top.MEM[47][27] ),
    .B2(_07771_),
    .X(_06617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13359_ (.A1_N(_07693_),
    .A2_N(_07768_),
    .B1(\design_top.MEM[47][26] ),
    .B2(_07770_),
    .X(_06616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13360_ (.A1_N(_07695_),
    .A2_N(_07768_),
    .B1(\design_top.MEM[47][25] ),
    .B2(_07770_),
    .X(_06615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13361_ (.A1_N(_07697_),
    .A2_N(_07768_),
    .B1(\design_top.MEM[47][24] ),
    .B2(_07770_),
    .X(_06614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13362_ (.A(_11102_),
    .B(_07450_),
    .X(_07772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13363_ (.A(_07727_),
    .B(_07772_),
    .X(_07773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13364_ (.A(_07773_),
    .X(_07774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13365_ (.A(_11271_),
    .X(_07775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _13366_ (.A(_11109_),
    .B(wbs_adr_i[2]),
    .C(_10895_),
    .D(wbs_adr_i[0]),
    .X(_07776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13367_ (.A(_07776_),
    .X(_07777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13368_ (.A(_07777_),
    .X(_07778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13369_ (.A1(_07775_),
    .A2(_07778_),
    .B1(_07773_),
    .X(_07779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13370_ (.A(_07779_),
    .X(_07780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13371_ (.A1_N(_07750_),
    .A2_N(_07774_),
    .B1(\design_top.MEM[40][15] ),
    .B2(_07780_),
    .X(_06613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13372_ (.A1_N(_07736_),
    .A2_N(_07774_),
    .B1(\design_top.MEM[40][14] ),
    .B2(_07780_),
    .X(_06612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13373_ (.A1_N(_07738_),
    .A2_N(_07774_),
    .B1(\design_top.MEM[40][13] ),
    .B2(_07780_),
    .X(_06611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13374_ (.A1_N(_07740_),
    .A2_N(_07774_),
    .B1(\design_top.MEM[40][12] ),
    .B2(_07780_),
    .X(_06610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13375_ (.A1_N(_07742_),
    .A2_N(_07774_),
    .B1(\design_top.MEM[40][11] ),
    .B2(_07780_),
    .X(_06609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13376_ (.A1_N(_07744_),
    .A2_N(_07773_),
    .B1(\design_top.MEM[40][10] ),
    .B2(_07779_),
    .X(_06608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13377_ (.A1_N(_07746_),
    .A2_N(_07773_),
    .B1(\design_top.MEM[40][9] ),
    .B2(_07779_),
    .X(_06607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13378_ (.A1_N(_07748_),
    .A2_N(_07773_),
    .B1(\design_top.MEM[40][8] ),
    .B2(_07779_),
    .X(_06606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13379_ (.A(_11102_),
    .B(_07557_),
    .X(_07781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13380_ (.A(_07727_),
    .B(_07781_),
    .X(_07782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13381_ (.A(_07782_),
    .X(_07783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13382_ (.A1(_07775_),
    .A2(_07564_),
    .B1(_07782_),
    .X(_07784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13383_ (.A(_07784_),
    .X(_07785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13384_ (.A1_N(_07750_),
    .A2_N(_07783_),
    .B1(\design_top.MEM[48][15] ),
    .B2(_07785_),
    .X(_06605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13385_ (.A1_N(_07736_),
    .A2_N(_07783_),
    .B1(\design_top.MEM[48][14] ),
    .B2(_07785_),
    .X(_06604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13386_ (.A1_N(_07738_),
    .A2_N(_07783_),
    .B1(\design_top.MEM[48][13] ),
    .B2(_07785_),
    .X(_06603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13387_ (.A1_N(_07740_),
    .A2_N(_07783_),
    .B1(\design_top.MEM[48][12] ),
    .B2(_07785_),
    .X(_06602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13388_ (.A1_N(_07742_),
    .A2_N(_07783_),
    .B1(\design_top.MEM[48][11] ),
    .B2(_07785_),
    .X(_06601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13389_ (.A1_N(_07744_),
    .A2_N(_07782_),
    .B1(\design_top.MEM[48][10] ),
    .B2(_07784_),
    .X(_06600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13390_ (.A1_N(_07746_),
    .A2_N(_07782_),
    .B1(\design_top.MEM[48][9] ),
    .B2(_07784_),
    .X(_06599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13391_ (.A1_N(_07748_),
    .A2_N(_07782_),
    .B1(\design_top.MEM[48][8] ),
    .B2(_07784_),
    .X(_06598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13392_ (.A(_07639_),
    .X(_07786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13393_ (.A(_07641_),
    .X(_07787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13394_ (.A(_07787_),
    .B(_07772_),
    .X(_07788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13395_ (.A(_07788_),
    .X(_07789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13396_ (.A1(_07775_),
    .A2(_07778_),
    .B1(_07788_),
    .X(_07790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13397_ (.A(_07790_),
    .X(_07791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13398_ (.A1_N(_07786_),
    .A2_N(_07789_),
    .B1(\design_top.MEM[40][23] ),
    .B2(_07791_),
    .X(_06597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13399_ (.A(_07648_),
    .X(_07792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13400_ (.A1_N(_07792_),
    .A2_N(_07789_),
    .B1(\design_top.MEM[40][22] ),
    .B2(_07791_),
    .X(_06596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13401_ (.A(_07650_),
    .X(_07793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13402_ (.A1_N(_07793_),
    .A2_N(_07789_),
    .B1(\design_top.MEM[40][21] ),
    .B2(_07791_),
    .X(_06595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13403_ (.A(_07652_),
    .X(_07794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13404_ (.A1_N(_07794_),
    .A2_N(_07789_),
    .B1(\design_top.MEM[40][20] ),
    .B2(_07791_),
    .X(_06594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13405_ (.A(_07654_),
    .X(_07795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13406_ (.A1_N(_07795_),
    .A2_N(_07789_),
    .B1(\design_top.MEM[40][19] ),
    .B2(_07791_),
    .X(_06593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13407_ (.A(_07656_),
    .X(_07796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13408_ (.A1_N(_07796_),
    .A2_N(_07788_),
    .B1(\design_top.MEM[40][18] ),
    .B2(_07790_),
    .X(_06592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13409_ (.A(_07658_),
    .X(_07797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13410_ (.A1_N(_07797_),
    .A2_N(_07788_),
    .B1(\design_top.MEM[40][17] ),
    .B2(_07790_),
    .X(_06591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13411_ (.A(_07660_),
    .X(_07798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13412_ (.A1_N(_07798_),
    .A2_N(_07788_),
    .B1(\design_top.MEM[40][16] ),
    .B2(_07790_),
    .X(_06590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13413_ (.A(_07676_),
    .X(_07799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13414_ (.A(_07678_),
    .X(_07800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13415_ (.A(_07800_),
    .B(_07772_),
    .X(_07801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13416_ (.A(_07801_),
    .X(_07802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13417_ (.A1(_07775_),
    .A2(_07778_),
    .B1(_07801_),
    .X(_07803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13418_ (.A(_07803_),
    .X(_07804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13419_ (.A1_N(_07799_),
    .A2_N(_07802_),
    .B1(\design_top.MEM[40][31] ),
    .B2(_07804_),
    .X(_06589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13420_ (.A(_07684_),
    .X(_07805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13421_ (.A1_N(_07805_),
    .A2_N(_07802_),
    .B1(\design_top.MEM[40][30] ),
    .B2(_07804_),
    .X(_06588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13422_ (.A(_07686_),
    .X(_07806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13423_ (.A1_N(_07806_),
    .A2_N(_07802_),
    .B1(\design_top.MEM[40][29] ),
    .B2(_07804_),
    .X(_06587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13424_ (.A(_07688_),
    .X(_07807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13425_ (.A1_N(_07807_),
    .A2_N(_07802_),
    .B1(\design_top.MEM[40][28] ),
    .B2(_07804_),
    .X(_06586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13426_ (.A(_07690_),
    .X(_07808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13427_ (.A1_N(_07808_),
    .A2_N(_07802_),
    .B1(\design_top.MEM[40][27] ),
    .B2(_07804_),
    .X(_06585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13428_ (.A(_07692_),
    .X(_07809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13429_ (.A1_N(_07809_),
    .A2_N(_07801_),
    .B1(\design_top.MEM[40][26] ),
    .B2(_07803_),
    .X(_06584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13430_ (.A(_07694_),
    .X(_07810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13431_ (.A1_N(_07810_),
    .A2_N(_07801_),
    .B1(\design_top.MEM[40][25] ),
    .B2(_07803_),
    .X(_06583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13432_ (.A(_07696_),
    .X(_07811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13433_ (.A1_N(_07811_),
    .A2_N(_07801_),
    .B1(\design_top.MEM[40][24] ),
    .B2(_07803_),
    .X(_06582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13434_ (.A(_07787_),
    .B(_07781_),
    .X(_07812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13435_ (.A(_07812_),
    .X(_07813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13436_ (.A(_07563_),
    .X(_07814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13437_ (.A1(_07775_),
    .A2(_07814_),
    .B1(_07812_),
    .X(_07815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13438_ (.A(_07815_),
    .X(_07816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13439_ (.A1_N(_07786_),
    .A2_N(_07813_),
    .B1(\design_top.MEM[48][23] ),
    .B2(_07816_),
    .X(_06581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13440_ (.A1_N(_07792_),
    .A2_N(_07813_),
    .B1(\design_top.MEM[48][22] ),
    .B2(_07816_),
    .X(_06580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13441_ (.A1_N(_07793_),
    .A2_N(_07813_),
    .B1(\design_top.MEM[48][21] ),
    .B2(_07816_),
    .X(_06579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13442_ (.A1_N(_07794_),
    .A2_N(_07813_),
    .B1(\design_top.MEM[48][20] ),
    .B2(_07816_),
    .X(_06578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13443_ (.A1_N(_07795_),
    .A2_N(_07813_),
    .B1(\design_top.MEM[48][19] ),
    .B2(_07816_),
    .X(_06577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13444_ (.A1_N(_07796_),
    .A2_N(_07812_),
    .B1(\design_top.MEM[48][18] ),
    .B2(_07815_),
    .X(_06576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13445_ (.A1_N(_07797_),
    .A2_N(_07812_),
    .B1(\design_top.MEM[48][17] ),
    .B2(_07815_),
    .X(_06575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13446_ (.A1_N(_07798_),
    .A2_N(_07812_),
    .B1(\design_top.MEM[48][16] ),
    .B2(_07815_),
    .X(_06574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13447_ (.A(_07800_),
    .B(_07781_),
    .X(_07817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13448_ (.A(_07817_),
    .X(_07818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13449_ (.A(_11271_),
    .X(_07819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13450_ (.A1(_07819_),
    .A2(_07814_),
    .B1(_07817_),
    .X(_07820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13451_ (.A(_07820_),
    .X(_07821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13452_ (.A1_N(_07799_),
    .A2_N(_07818_),
    .B1(\design_top.MEM[48][31] ),
    .B2(_07821_),
    .X(_06573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13453_ (.A1_N(_07805_),
    .A2_N(_07818_),
    .B1(\design_top.MEM[48][30] ),
    .B2(_07821_),
    .X(_06572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13454_ (.A1_N(_07806_),
    .A2_N(_07818_),
    .B1(\design_top.MEM[48][29] ),
    .B2(_07821_),
    .X(_06571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13455_ (.A1_N(_07807_),
    .A2_N(_07818_),
    .B1(\design_top.MEM[48][28] ),
    .B2(_07821_),
    .X(_06570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13456_ (.A1_N(_07808_),
    .A2_N(_07818_),
    .B1(\design_top.MEM[48][27] ),
    .B2(_07821_),
    .X(_06569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13457_ (.A1_N(_07809_),
    .A2_N(_07817_),
    .B1(\design_top.MEM[48][26] ),
    .B2(_07820_),
    .X(_06568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13458_ (.A1_N(_07810_),
    .A2_N(_07817_),
    .B1(\design_top.MEM[48][25] ),
    .B2(_07820_),
    .X(_06567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13459_ (.A1_N(_07811_),
    .A2_N(_07817_),
    .B1(\design_top.MEM[48][24] ),
    .B2(_07820_),
    .X(_06566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13460_ (.A(_11275_),
    .B(_07450_),
    .X(_07822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13461_ (.A(_07727_),
    .B(_07822_),
    .X(_07823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13462_ (.A(_07823_),
    .X(_07824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13463_ (.A1(_07668_),
    .A2(_07778_),
    .B1(_07823_),
    .X(_07825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13464_ (.A(_07825_),
    .X(_07826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13465_ (.A1_N(_07750_),
    .A2_N(_07824_),
    .B1(\design_top.MEM[41][15] ),
    .B2(_07826_),
    .X(_06565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13466_ (.A1_N(_07736_),
    .A2_N(_07824_),
    .B1(\design_top.MEM[41][14] ),
    .B2(_07826_),
    .X(_06564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13467_ (.A1_N(_07738_),
    .A2_N(_07824_),
    .B1(\design_top.MEM[41][13] ),
    .B2(_07826_),
    .X(_06563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13468_ (.A1_N(_07740_),
    .A2_N(_07824_),
    .B1(\design_top.MEM[41][12] ),
    .B2(_07826_),
    .X(_06562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13469_ (.A1_N(_07742_),
    .A2_N(_07824_),
    .B1(\design_top.MEM[41][11] ),
    .B2(_07826_),
    .X(_06561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13470_ (.A1_N(_07744_),
    .A2_N(_07823_),
    .B1(\design_top.MEM[41][10] ),
    .B2(_07825_),
    .X(_06560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13471_ (.A1_N(_07746_),
    .A2_N(_07823_),
    .B1(\design_top.MEM[41][9] ),
    .B2(_07825_),
    .X(_06559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13472_ (.A1_N(_07748_),
    .A2_N(_07823_),
    .B1(\design_top.MEM[41][8] ),
    .B2(_07825_),
    .X(_06558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13473_ (.A(_07726_),
    .X(_07827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13474_ (.A(_11275_),
    .B(_07557_),
    .X(_07828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13475_ (.A(_07827_),
    .B(_07828_),
    .X(_07829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13476_ (.A(_07829_),
    .X(_07830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13477_ (.A1(_07668_),
    .A2(_07814_),
    .B1(_07829_),
    .X(_07831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13478_ (.A(_07831_),
    .X(_07832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13479_ (.A1_N(_07750_),
    .A2_N(_07830_),
    .B1(\design_top.MEM[49][15] ),
    .B2(_07832_),
    .X(_06557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13480_ (.A(_07735_),
    .X(_07833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13481_ (.A1_N(_07833_),
    .A2_N(_07830_),
    .B1(\design_top.MEM[49][14] ),
    .B2(_07832_),
    .X(_06556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13482_ (.A(_07737_),
    .X(_07834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13483_ (.A1_N(_07834_),
    .A2_N(_07830_),
    .B1(\design_top.MEM[49][13] ),
    .B2(_07832_),
    .X(_06555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13484_ (.A(_07739_),
    .X(_07835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13485_ (.A1_N(_07835_),
    .A2_N(_07830_),
    .B1(\design_top.MEM[49][12] ),
    .B2(_07832_),
    .X(_06554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13486_ (.A(_07741_),
    .X(_07836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13487_ (.A1_N(_07836_),
    .A2_N(_07830_),
    .B1(\design_top.MEM[49][11] ),
    .B2(_07832_),
    .X(_06553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13488_ (.A(_07743_),
    .X(_07837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13489_ (.A1_N(_07837_),
    .A2_N(_07829_),
    .B1(\design_top.MEM[49][10] ),
    .B2(_07831_),
    .X(_06552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13490_ (.A(_07745_),
    .X(_07838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13491_ (.A1_N(_07838_),
    .A2_N(_07829_),
    .B1(\design_top.MEM[49][9] ),
    .B2(_07831_),
    .X(_06551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13492_ (.A(_07747_),
    .X(_07839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13493_ (.A1_N(_07839_),
    .A2_N(_07829_),
    .B1(\design_top.MEM[49][8] ),
    .B2(_07831_),
    .X(_06550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13494_ (.A(_07787_),
    .B(_07822_),
    .X(_07840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13495_ (.A(_07840_),
    .X(_07841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13496_ (.A1(_07668_),
    .A2(_07778_),
    .B1(_07840_),
    .X(_07842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13497_ (.A(_07842_),
    .X(_07843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13498_ (.A1_N(_07786_),
    .A2_N(_07841_),
    .B1(\design_top.MEM[41][23] ),
    .B2(_07843_),
    .X(_06549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13499_ (.A1_N(_07792_),
    .A2_N(_07841_),
    .B1(\design_top.MEM[41][22] ),
    .B2(_07843_),
    .X(_06548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13500_ (.A1_N(_07793_),
    .A2_N(_07841_),
    .B1(\design_top.MEM[41][21] ),
    .B2(_07843_),
    .X(_06547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13501_ (.A1_N(_07794_),
    .A2_N(_07841_),
    .B1(\design_top.MEM[41][20] ),
    .B2(_07843_),
    .X(_06546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13502_ (.A1_N(_07795_),
    .A2_N(_07841_),
    .B1(\design_top.MEM[41][19] ),
    .B2(_07843_),
    .X(_06545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13503_ (.A1_N(_07796_),
    .A2_N(_07840_),
    .B1(\design_top.MEM[41][18] ),
    .B2(_07842_),
    .X(_06544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13504_ (.A1_N(_07797_),
    .A2_N(_07840_),
    .B1(\design_top.MEM[41][17] ),
    .B2(_07842_),
    .X(_06543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13505_ (.A1_N(_07798_),
    .A2_N(_07840_),
    .B1(\design_top.MEM[41][16] ),
    .B2(_07842_),
    .X(_06542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13506_ (.A(_07800_),
    .B(_07822_),
    .X(_07844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13507_ (.A(_07844_),
    .X(_07845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13508_ (.A(_07508_),
    .X(_07846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13509_ (.A(_07777_),
    .X(_07847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13510_ (.A1(_07846_),
    .A2(_07847_),
    .B1(_07844_),
    .X(_07848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13511_ (.A(_07848_),
    .X(_07849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13512_ (.A1_N(_07799_),
    .A2_N(_07845_),
    .B1(\design_top.MEM[41][31] ),
    .B2(_07849_),
    .X(_06541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13513_ (.A1_N(_07805_),
    .A2_N(_07845_),
    .B1(\design_top.MEM[41][30] ),
    .B2(_07849_),
    .X(_06540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13514_ (.A1_N(_07806_),
    .A2_N(_07845_),
    .B1(\design_top.MEM[41][29] ),
    .B2(_07849_),
    .X(_06539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13515_ (.A1_N(_07807_),
    .A2_N(_07845_),
    .B1(\design_top.MEM[41][28] ),
    .B2(_07849_),
    .X(_06538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13516_ (.A1_N(_07808_),
    .A2_N(_07845_),
    .B1(\design_top.MEM[41][27] ),
    .B2(_07849_),
    .X(_06537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13517_ (.A1_N(_07809_),
    .A2_N(_07844_),
    .B1(\design_top.MEM[41][26] ),
    .B2(_07848_),
    .X(_06536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13518_ (.A1_N(_07810_),
    .A2_N(_07844_),
    .B1(\design_top.MEM[41][25] ),
    .B2(_07848_),
    .X(_06535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13519_ (.A1_N(_07811_),
    .A2_N(_07844_),
    .B1(\design_top.MEM[41][24] ),
    .B2(_07848_),
    .X(_06534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13520_ (.A(_07749_),
    .X(_07850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13521_ (.A(_10999_),
    .B(_07449_),
    .X(_07851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13522_ (.A(_07827_),
    .B(_07851_),
    .X(_07852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13523_ (.A(_07852_),
    .X(_07853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13524_ (.A1(_07715_),
    .A2(_07847_),
    .B1(_07852_),
    .X(_07854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13525_ (.A(_07854_),
    .X(_07855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13526_ (.A1_N(_07850_),
    .A2_N(_07853_),
    .B1(\design_top.MEM[42][15] ),
    .B2(_07855_),
    .X(_06533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13527_ (.A1_N(_07833_),
    .A2_N(_07853_),
    .B1(\design_top.MEM[42][14] ),
    .B2(_07855_),
    .X(_06532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13528_ (.A1_N(_07834_),
    .A2_N(_07853_),
    .B1(\design_top.MEM[42][13] ),
    .B2(_07855_),
    .X(_06531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13529_ (.A1_N(_07835_),
    .A2_N(_07853_),
    .B1(\design_top.MEM[42][12] ),
    .B2(_07855_),
    .X(_06530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13530_ (.A1_N(_07836_),
    .A2_N(_07853_),
    .B1(\design_top.MEM[42][11] ),
    .B2(_07855_),
    .X(_06529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13531_ (.A1_N(_07837_),
    .A2_N(_07852_),
    .B1(\design_top.MEM[42][10] ),
    .B2(_07854_),
    .X(_06528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13532_ (.A1_N(_07838_),
    .A2_N(_07852_),
    .B1(\design_top.MEM[42][9] ),
    .B2(_07854_),
    .X(_06527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13533_ (.A1_N(_07839_),
    .A2_N(_07852_),
    .B1(\design_top.MEM[42][8] ),
    .B2(_07854_),
    .X(_06526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13534_ (.A(_07787_),
    .B(_07828_),
    .X(_07856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13535_ (.A(_07856_),
    .X(_07857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13536_ (.A1(_07846_),
    .A2(_07814_),
    .B1(_07856_),
    .X(_07858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13537_ (.A(_07858_),
    .X(_07859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13538_ (.A1_N(_07786_),
    .A2_N(_07857_),
    .B1(\design_top.MEM[49][23] ),
    .B2(_07859_),
    .X(_06525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13539_ (.A1_N(_07792_),
    .A2_N(_07857_),
    .B1(\design_top.MEM[49][22] ),
    .B2(_07859_),
    .X(_06524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13540_ (.A1_N(_07793_),
    .A2_N(_07857_),
    .B1(\design_top.MEM[49][21] ),
    .B2(_07859_),
    .X(_06523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13541_ (.A1_N(_07794_),
    .A2_N(_07857_),
    .B1(\design_top.MEM[49][20] ),
    .B2(_07859_),
    .X(_06522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13542_ (.A1_N(_07795_),
    .A2_N(_07857_),
    .B1(\design_top.MEM[49][19] ),
    .B2(_07859_),
    .X(_06521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13543_ (.A1_N(_07796_),
    .A2_N(_07856_),
    .B1(\design_top.MEM[49][18] ),
    .B2(_07858_),
    .X(_06520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13544_ (.A1_N(_07797_),
    .A2_N(_07856_),
    .B1(\design_top.MEM[49][17] ),
    .B2(_07858_),
    .X(_06519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13545_ (.A1_N(_07798_),
    .A2_N(_07856_),
    .B1(\design_top.MEM[49][16] ),
    .B2(_07858_),
    .X(_06518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13546_ (.A(_07800_),
    .B(_07828_),
    .X(_07860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13547_ (.A(_07860_),
    .X(_07861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13548_ (.A1(_07846_),
    .A2(_07814_),
    .B1(_07860_),
    .X(_07862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13549_ (.A(_07862_),
    .X(_07863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13550_ (.A1_N(_07799_),
    .A2_N(_07861_),
    .B1(\design_top.MEM[49][31] ),
    .B2(_07863_),
    .X(_06517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13551_ (.A1_N(_07805_),
    .A2_N(_07861_),
    .B1(\design_top.MEM[49][30] ),
    .B2(_07863_),
    .X(_06516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13552_ (.A1_N(_07806_),
    .A2_N(_07861_),
    .B1(\design_top.MEM[49][29] ),
    .B2(_07863_),
    .X(_06515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13553_ (.A1_N(_07807_),
    .A2_N(_07861_),
    .B1(\design_top.MEM[49][28] ),
    .B2(_07863_),
    .X(_06514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13554_ (.A1_N(_07808_),
    .A2_N(_07861_),
    .B1(\design_top.MEM[49][27] ),
    .B2(_07863_),
    .X(_06513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13555_ (.A1_N(_07809_),
    .A2_N(_07860_),
    .B1(\design_top.MEM[49][26] ),
    .B2(_07862_),
    .X(_06512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13556_ (.A1_N(_07810_),
    .A2_N(_07860_),
    .B1(\design_top.MEM[49][25] ),
    .B2(_07862_),
    .X(_06511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13557_ (.A1_N(_07811_),
    .A2_N(_07860_),
    .B1(\design_top.MEM[49][24] ),
    .B2(_07862_),
    .X(_06510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13558_ (.A(_10783_),
    .B(_10958_),
    .X(_07864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13559_ (.A(_07827_),
    .B(_07864_),
    .X(_07865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13560_ (.A(_07865_),
    .X(_07866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _13561_ (.A(wbs_adr_i[3]),
    .B(wbs_adr_i[2]),
    .C(wbs_adr_i[1]),
    .D(_10963_),
    .X(_07867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13562_ (.A(_07867_),
    .X(_07868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13563_ (.A(_07868_),
    .X(_07869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13564_ (.A1(_07819_),
    .A2(_07869_),
    .B1(_07865_),
    .X(_07870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13565_ (.A(_07870_),
    .X(_07871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13566_ (.A1_N(_07850_),
    .A2_N(_07866_),
    .B1(\design_top.MEM[4][15] ),
    .B2(_07871_),
    .X(_06509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13567_ (.A1_N(_07833_),
    .A2_N(_07866_),
    .B1(\design_top.MEM[4][14] ),
    .B2(_07871_),
    .X(_06508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13568_ (.A1_N(_07834_),
    .A2_N(_07866_),
    .B1(\design_top.MEM[4][13] ),
    .B2(_07871_),
    .X(_06507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13569_ (.A1_N(_07835_),
    .A2_N(_07866_),
    .B1(\design_top.MEM[4][12] ),
    .B2(_07871_),
    .X(_06506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13570_ (.A1_N(_07836_),
    .A2_N(_07866_),
    .B1(\design_top.MEM[4][11] ),
    .B2(_07871_),
    .X(_06505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13571_ (.A1_N(_07837_),
    .A2_N(_07865_),
    .B1(\design_top.MEM[4][10] ),
    .B2(_07870_),
    .X(_06504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13572_ (.A1_N(_07838_),
    .A2_N(_07865_),
    .B1(\design_top.MEM[4][9] ),
    .B2(_07870_),
    .X(_06503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13573_ (.A1_N(_07839_),
    .A2_N(_07865_),
    .B1(\design_top.MEM[4][8] ),
    .B2(_07870_),
    .X(_06502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13574_ (.A(_07787_),
    .B(_07851_),
    .X(_07872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13575_ (.A(_07872_),
    .X(_07873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13576_ (.A1(_07715_),
    .A2(_07847_),
    .B1(_07872_),
    .X(_07874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13577_ (.A(_07874_),
    .X(_07875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13578_ (.A1_N(_07786_),
    .A2_N(_07873_),
    .B1(\design_top.MEM[42][23] ),
    .B2(_07875_),
    .X(_06501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13579_ (.A1_N(_07792_),
    .A2_N(_07873_),
    .B1(\design_top.MEM[42][22] ),
    .B2(_07875_),
    .X(_06500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13580_ (.A1_N(_07793_),
    .A2_N(_07873_),
    .B1(\design_top.MEM[42][21] ),
    .B2(_07875_),
    .X(_06499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13581_ (.A1_N(_07794_),
    .A2_N(_07873_),
    .B1(\design_top.MEM[42][20] ),
    .B2(_07875_),
    .X(_06498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13582_ (.A1_N(_07795_),
    .A2_N(_07873_),
    .B1(\design_top.MEM[42][19] ),
    .B2(_07875_),
    .X(_06497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13583_ (.A1_N(_07796_),
    .A2_N(_07872_),
    .B1(\design_top.MEM[42][18] ),
    .B2(_07874_),
    .X(_06496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13584_ (.A1_N(_07797_),
    .A2_N(_07872_),
    .B1(\design_top.MEM[42][17] ),
    .B2(_07874_),
    .X(_06495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13585_ (.A1_N(_07798_),
    .A2_N(_07872_),
    .B1(\design_top.MEM[42][16] ),
    .B2(_07874_),
    .X(_06494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13586_ (.A(_07800_),
    .B(_07851_),
    .X(_07876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13587_ (.A(_07876_),
    .X(_07877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13588_ (.A1(_07715_),
    .A2(_07847_),
    .B1(_07876_),
    .X(_07878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13589_ (.A(_07878_),
    .X(_07879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13590_ (.A1_N(_07799_),
    .A2_N(_07877_),
    .B1(\design_top.MEM[42][31] ),
    .B2(_07879_),
    .X(_06493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13591_ (.A1_N(_07805_),
    .A2_N(_07877_),
    .B1(\design_top.MEM[42][30] ),
    .B2(_07879_),
    .X(_06492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13592_ (.A1_N(_07806_),
    .A2_N(_07877_),
    .B1(\design_top.MEM[42][29] ),
    .B2(_07879_),
    .X(_06491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13593_ (.A1_N(_07807_),
    .A2_N(_07877_),
    .B1(\design_top.MEM[42][28] ),
    .B2(_07879_),
    .X(_06490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13594_ (.A1_N(_07808_),
    .A2_N(_07877_),
    .B1(\design_top.MEM[42][27] ),
    .B2(_07879_),
    .X(_06489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13595_ (.A1_N(_07809_),
    .A2_N(_07876_),
    .B1(\design_top.MEM[42][26] ),
    .B2(_07878_),
    .X(_06488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13596_ (.A1_N(_07810_),
    .A2_N(_07876_),
    .B1(\design_top.MEM[42][25] ),
    .B2(_07878_),
    .X(_06487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13597_ (.A1_N(_07811_),
    .A2_N(_07876_),
    .B1(\design_top.MEM[42][24] ),
    .B2(_07878_),
    .X(_06486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13598_ (.A(_07639_),
    .X(_07880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13599_ (.A(_07641_),
    .X(_07881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13600_ (.A(_07881_),
    .B(_07864_),
    .X(_07882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13601_ (.A(_07882_),
    .X(_07883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13602_ (.A1(_07819_),
    .A2(_07869_),
    .B1(_07882_),
    .X(_07884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13603_ (.A(_07884_),
    .X(_07885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13604_ (.A1_N(_07880_),
    .A2_N(_07883_),
    .B1(\design_top.MEM[4][23] ),
    .B2(_07885_),
    .X(_06485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13605_ (.A(_07648_),
    .X(_07886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13606_ (.A1_N(_07886_),
    .A2_N(_07883_),
    .B1(\design_top.MEM[4][22] ),
    .B2(_07885_),
    .X(_06484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13607_ (.A(_07650_),
    .X(_07887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13608_ (.A1_N(_07887_),
    .A2_N(_07883_),
    .B1(\design_top.MEM[4][21] ),
    .B2(_07885_),
    .X(_06483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13609_ (.A(_07652_),
    .X(_07888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13610_ (.A1_N(_07888_),
    .A2_N(_07883_),
    .B1(\design_top.MEM[4][20] ),
    .B2(_07885_),
    .X(_06482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13611_ (.A(_07654_),
    .X(_07889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13612_ (.A1_N(_07889_),
    .A2_N(_07883_),
    .B1(\design_top.MEM[4][19] ),
    .B2(_07885_),
    .X(_06481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13613_ (.A(_07656_),
    .X(_07890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13614_ (.A1_N(_07890_),
    .A2_N(_07882_),
    .B1(\design_top.MEM[4][18] ),
    .B2(_07884_),
    .X(_06480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13615_ (.A(_07658_),
    .X(_07891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13616_ (.A1_N(_07891_),
    .A2_N(_07882_),
    .B1(\design_top.MEM[4][17] ),
    .B2(_07884_),
    .X(_06479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13617_ (.A(_07660_),
    .X(_07892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13618_ (.A1_N(_07892_),
    .A2_N(_07882_),
    .B1(\design_top.MEM[4][16] ),
    .B2(_07884_),
    .X(_06478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13619_ (.A(_07676_),
    .X(_07893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13620_ (.A(_07678_),
    .X(_07894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13621_ (.A(_07894_),
    .B(_07864_),
    .X(_07895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13622_ (.A(_07895_),
    .X(_07896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13623_ (.A1(_07819_),
    .A2(_07869_),
    .B1(_07895_),
    .X(_07897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13624_ (.A(_07897_),
    .X(_07898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13625_ (.A1_N(_07893_),
    .A2_N(_07896_),
    .B1(\design_top.MEM[4][31] ),
    .B2(_07898_),
    .X(_06477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13626_ (.A(_07684_),
    .X(_07899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13627_ (.A1_N(_07899_),
    .A2_N(_07896_),
    .B1(\design_top.MEM[4][30] ),
    .B2(_07898_),
    .X(_06476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13628_ (.A(_07686_),
    .X(_07900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13629_ (.A1_N(_07900_),
    .A2_N(_07896_),
    .B1(\design_top.MEM[4][29] ),
    .B2(_07898_),
    .X(_06475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13630_ (.A(_07688_),
    .X(_07901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13631_ (.A1_N(_07901_),
    .A2_N(_07896_),
    .B1(\design_top.MEM[4][28] ),
    .B2(_07898_),
    .X(_06474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13632_ (.A(_07690_),
    .X(_07902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13633_ (.A1_N(_07902_),
    .A2_N(_07896_),
    .B1(\design_top.MEM[4][27] ),
    .B2(_07898_),
    .X(_06473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13634_ (.A(_07692_),
    .X(_07903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13635_ (.A1_N(_07903_),
    .A2_N(_07895_),
    .B1(\design_top.MEM[4][26] ),
    .B2(_07897_),
    .X(_06472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13636_ (.A(_07694_),
    .X(_07904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13637_ (.A1_N(_07904_),
    .A2_N(_07895_),
    .B1(\design_top.MEM[4][25] ),
    .B2(_07897_),
    .X(_06471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13638_ (.A(_07696_),
    .X(_07905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13639_ (.A1_N(_07905_),
    .A2_N(_07895_),
    .B1(\design_top.MEM[4][24] ),
    .B2(_07897_),
    .X(_06470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13640_ (.A(_10884_),
    .B(_07449_),
    .X(_07906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13641_ (.A(_07827_),
    .B(_07906_),
    .X(_07907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13642_ (.A(_07907_),
    .X(_07908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13643_ (.A1(_07731_),
    .A2(_07847_),
    .B1(_07907_),
    .X(_07909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13644_ (.A(_07909_),
    .X(_07910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13645_ (.A1_N(_07850_),
    .A2_N(_07908_),
    .B1(\design_top.MEM[43][15] ),
    .B2(_07910_),
    .X(_06469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13646_ (.A1_N(_07833_),
    .A2_N(_07908_),
    .B1(\design_top.MEM[43][14] ),
    .B2(_07910_),
    .X(_06468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13647_ (.A1_N(_07834_),
    .A2_N(_07908_),
    .B1(\design_top.MEM[43][13] ),
    .B2(_07910_),
    .X(_06467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13648_ (.A1_N(_07835_),
    .A2_N(_07908_),
    .B1(\design_top.MEM[43][12] ),
    .B2(_07910_),
    .X(_06466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13649_ (.A1_N(_07836_),
    .A2_N(_07908_),
    .B1(\design_top.MEM[43][11] ),
    .B2(_07910_),
    .X(_06465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13650_ (.A1_N(_07837_),
    .A2_N(_07907_),
    .B1(\design_top.MEM[43][10] ),
    .B2(_07909_),
    .X(_06464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13651_ (.A1_N(_07838_),
    .A2_N(_07907_),
    .B1(\design_top.MEM[43][9] ),
    .B2(_07909_),
    .X(_06463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13652_ (.A1_N(_07839_),
    .A2_N(_07907_),
    .B1(\design_top.MEM[43][8] ),
    .B2(_07909_),
    .X(_06462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13653_ (.A(_07827_),
    .B(_07559_),
    .X(_07911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13654_ (.A(_07911_),
    .X(_07912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13655_ (.A(_07434_),
    .X(_07913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13656_ (.A1(_07913_),
    .A2(_07563_),
    .B1(_07911_),
    .X(_07914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13657_ (.A(_07914_),
    .X(_07915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13658_ (.A1_N(_07850_),
    .A2_N(_07912_),
    .B1(\design_top.MEM[50][15] ),
    .B2(_07915_),
    .X(_06461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13659_ (.A1_N(_07833_),
    .A2_N(_07912_),
    .B1(\design_top.MEM[50][14] ),
    .B2(_07915_),
    .X(_06460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13660_ (.A1_N(_07834_),
    .A2_N(_07912_),
    .B1(\design_top.MEM[50][13] ),
    .B2(_07915_),
    .X(_06459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13661_ (.A1_N(_07835_),
    .A2_N(_07912_),
    .B1(\design_top.MEM[50][12] ),
    .B2(_07915_),
    .X(_06458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13662_ (.A1_N(_07836_),
    .A2_N(_07912_),
    .B1(\design_top.MEM[50][11] ),
    .B2(_07915_),
    .X(_06457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13663_ (.A1_N(_07837_),
    .A2_N(_07911_),
    .B1(\design_top.MEM[50][10] ),
    .B2(_07914_),
    .X(_06456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13664_ (.A1_N(_07838_),
    .A2_N(_07911_),
    .B1(\design_top.MEM[50][9] ),
    .B2(_07914_),
    .X(_06455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13665_ (.A1_N(_07839_),
    .A2_N(_07911_),
    .B1(\design_top.MEM[50][8] ),
    .B2(_07914_),
    .X(_06454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13666_ (.A(_07881_),
    .B(_07906_),
    .X(_07916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13667_ (.A(_07916_),
    .X(_07917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13668_ (.A1(_07731_),
    .A2(_07777_),
    .B1(_07916_),
    .X(_07918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13669_ (.A(_07918_),
    .X(_07919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13670_ (.A1_N(_07880_),
    .A2_N(_07917_),
    .B1(\design_top.MEM[43][23] ),
    .B2(_07919_),
    .X(_06453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13671_ (.A1_N(_07886_),
    .A2_N(_07917_),
    .B1(\design_top.MEM[43][22] ),
    .B2(_07919_),
    .X(_06452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13672_ (.A1_N(_07887_),
    .A2_N(_07917_),
    .B1(\design_top.MEM[43][21] ),
    .B2(_07919_),
    .X(_06451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13673_ (.A1_N(_07888_),
    .A2_N(_07917_),
    .B1(\design_top.MEM[43][20] ),
    .B2(_07919_),
    .X(_06450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13674_ (.A1_N(_07889_),
    .A2_N(_07917_),
    .B1(\design_top.MEM[43][19] ),
    .B2(_07919_),
    .X(_06449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13675_ (.A1_N(_07890_),
    .A2_N(_07916_),
    .B1(\design_top.MEM[43][18] ),
    .B2(_07918_),
    .X(_06448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13676_ (.A1_N(_07891_),
    .A2_N(_07916_),
    .B1(\design_top.MEM[43][17] ),
    .B2(_07918_),
    .X(_06447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13677_ (.A1_N(_07892_),
    .A2_N(_07916_),
    .B1(\design_top.MEM[43][16] ),
    .B2(_07918_),
    .X(_06446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13678_ (.A(_07894_),
    .B(_07906_),
    .X(_07920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13679_ (.A(_07920_),
    .X(_07921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13680_ (.A(_11251_),
    .X(_07922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13681_ (.A1(_07922_),
    .A2(_07777_),
    .B1(_07920_),
    .X(_07923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13682_ (.A(_07923_),
    .X(_07924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13683_ (.A1_N(_07893_),
    .A2_N(_07921_),
    .B1(\design_top.MEM[43][31] ),
    .B2(_07924_),
    .X(_06445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13684_ (.A1_N(_07899_),
    .A2_N(_07921_),
    .B1(\design_top.MEM[43][30] ),
    .B2(_07924_),
    .X(_06444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13685_ (.A1_N(_07900_),
    .A2_N(_07921_),
    .B1(\design_top.MEM[43][29] ),
    .B2(_07924_),
    .X(_06443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13686_ (.A1_N(_07901_),
    .A2_N(_07921_),
    .B1(\design_top.MEM[43][28] ),
    .B2(_07924_),
    .X(_06442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13687_ (.A1_N(_07902_),
    .A2_N(_07921_),
    .B1(\design_top.MEM[43][27] ),
    .B2(_07924_),
    .X(_06441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13688_ (.A1_N(_07903_),
    .A2_N(_07920_),
    .B1(\design_top.MEM[43][26] ),
    .B2(_07923_),
    .X(_06440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13689_ (.A1_N(_07904_),
    .A2_N(_07920_),
    .B1(\design_top.MEM[43][25] ),
    .B2(_07923_),
    .X(_06439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13690_ (.A1_N(_07905_),
    .A2_N(_07920_),
    .B1(\design_top.MEM[43][24] ),
    .B2(_07923_),
    .X(_06438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13691_ (.A(_07881_),
    .B(_07559_),
    .X(_07925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13692_ (.A(_07925_),
    .X(_07926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13693_ (.A1(_07913_),
    .A2(_07563_),
    .B1(_07925_),
    .X(_07927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13694_ (.A(_07927_),
    .X(_07928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13695_ (.A1_N(_07880_),
    .A2_N(_07926_),
    .B1(\design_top.MEM[50][23] ),
    .B2(_07928_),
    .X(_06437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13696_ (.A1_N(_07886_),
    .A2_N(_07926_),
    .B1(\design_top.MEM[50][22] ),
    .B2(_07928_),
    .X(_06436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13697_ (.A1_N(_07887_),
    .A2_N(_07926_),
    .B1(\design_top.MEM[50][21] ),
    .B2(_07928_),
    .X(_06435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13698_ (.A1_N(_07888_),
    .A2_N(_07926_),
    .B1(\design_top.MEM[50][20] ),
    .B2(_07928_),
    .X(_06434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13699_ (.A1_N(_07889_),
    .A2_N(_07926_),
    .B1(\design_top.MEM[50][19] ),
    .B2(_07928_),
    .X(_06433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13700_ (.A1_N(_07890_),
    .A2_N(_07925_),
    .B1(\design_top.MEM[50][18] ),
    .B2(_07927_),
    .X(_06432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13701_ (.A1_N(_07891_),
    .A2_N(_07925_),
    .B1(\design_top.MEM[50][17] ),
    .B2(_07927_),
    .X(_06431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13702_ (.A1_N(_07892_),
    .A2_N(_07925_),
    .B1(\design_top.MEM[50][16] ),
    .B2(_07927_),
    .X(_06430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13703_ (.A(_07726_),
    .X(_07929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13704_ (.A(_10957_),
    .B(_07449_),
    .X(_07930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13705_ (.A(_07929_),
    .B(_07930_),
    .X(_07931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13706_ (.A(_07931_),
    .X(_07932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13707_ (.A1(_07819_),
    .A2(_07732_),
    .B1(_07931_),
    .X(_07933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13708_ (.A(_07933_),
    .X(_07934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13709_ (.A1_N(_07850_),
    .A2_N(_07932_),
    .B1(\design_top.MEM[44][15] ),
    .B2(_07934_),
    .X(_06429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13710_ (.A(_07735_),
    .X(_07935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13711_ (.A1_N(_07935_),
    .A2_N(_07932_),
    .B1(\design_top.MEM[44][14] ),
    .B2(_07934_),
    .X(_06428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13712_ (.A(_07737_),
    .X(_07936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13713_ (.A1_N(_07936_),
    .A2_N(_07932_),
    .B1(\design_top.MEM[44][13] ),
    .B2(_07934_),
    .X(_06427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13714_ (.A(_07739_),
    .X(_07937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13715_ (.A1_N(_07937_),
    .A2_N(_07932_),
    .B1(\design_top.MEM[44][12] ),
    .B2(_07934_),
    .X(_06426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13716_ (.A(_07741_),
    .X(_07938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13717_ (.A1_N(_07938_),
    .A2_N(_07932_),
    .B1(\design_top.MEM[44][11] ),
    .B2(_07934_),
    .X(_06425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13718_ (.A(_07743_),
    .X(_07939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13719_ (.A1_N(_07939_),
    .A2_N(_07931_),
    .B1(\design_top.MEM[44][10] ),
    .B2(_07933_),
    .X(_06424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13720_ (.A(_07745_),
    .X(_07940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13721_ (.A1_N(_07940_),
    .A2_N(_07931_),
    .B1(\design_top.MEM[44][9] ),
    .B2(_07933_),
    .X(_06423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13722_ (.A(_07747_),
    .X(_07941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13723_ (.A1_N(_07941_),
    .A2_N(_07931_),
    .B1(\design_top.MEM[44][8] ),
    .B2(_07933_),
    .X(_06422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13724_ (.A(_07881_),
    .B(_07930_),
    .X(_07942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13725_ (.A(_07942_),
    .X(_07943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13726_ (.A(_11271_),
    .X(_07944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13727_ (.A1(_07944_),
    .A2(_07732_),
    .B1(_07942_),
    .X(_07945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13728_ (.A(_07945_),
    .X(_07946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13729_ (.A1_N(_07880_),
    .A2_N(_07943_),
    .B1(\design_top.MEM[44][23] ),
    .B2(_07946_),
    .X(_06421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13730_ (.A1_N(_07886_),
    .A2_N(_07943_),
    .B1(\design_top.MEM[44][22] ),
    .B2(_07946_),
    .X(_06420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13731_ (.A1_N(_07887_),
    .A2_N(_07943_),
    .B1(\design_top.MEM[44][21] ),
    .B2(_07946_),
    .X(_06419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13732_ (.A1_N(_07888_),
    .A2_N(_07943_),
    .B1(\design_top.MEM[44][20] ),
    .B2(_07946_),
    .X(_06418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13733_ (.A1_N(_07889_),
    .A2_N(_07943_),
    .B1(\design_top.MEM[44][19] ),
    .B2(_07946_),
    .X(_06417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13734_ (.A1_N(_07890_),
    .A2_N(_07942_),
    .B1(\design_top.MEM[44][18] ),
    .B2(_07945_),
    .X(_06416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13735_ (.A1_N(_07891_),
    .A2_N(_07942_),
    .B1(\design_top.MEM[44][17] ),
    .B2(_07945_),
    .X(_06415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13736_ (.A1_N(_07892_),
    .A2_N(_07942_),
    .B1(\design_top.MEM[44][16] ),
    .B2(_07945_),
    .X(_06414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13737_ (.A(_07894_),
    .B(_07930_),
    .X(_07947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13738_ (.A(_07947_),
    .X(_07948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13739_ (.A1(_07944_),
    .A2(_07455_),
    .B1(_07947_),
    .X(_07949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13740_ (.A(_07949_),
    .X(_07950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13741_ (.A1_N(_07893_),
    .A2_N(_07948_),
    .B1(\design_top.MEM[44][31] ),
    .B2(_07950_),
    .X(_06413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13742_ (.A1_N(_07899_),
    .A2_N(_07948_),
    .B1(\design_top.MEM[44][30] ),
    .B2(_07950_),
    .X(_06412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13743_ (.A1_N(_07900_),
    .A2_N(_07948_),
    .B1(\design_top.MEM[44][29] ),
    .B2(_07950_),
    .X(_06411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13744_ (.A1_N(_07901_),
    .A2_N(_07948_),
    .B1(\design_top.MEM[44][28] ),
    .B2(_07950_),
    .X(_06410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13745_ (.A1_N(_07902_),
    .A2_N(_07948_),
    .B1(\design_top.MEM[44][27] ),
    .B2(_07950_),
    .X(_06409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13746_ (.A1_N(_07903_),
    .A2_N(_07947_),
    .B1(\design_top.MEM[44][26] ),
    .B2(_07949_),
    .X(_06408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13747_ (.A1_N(_07904_),
    .A2_N(_07947_),
    .B1(\design_top.MEM[44][25] ),
    .B2(_07949_),
    .X(_06407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13748_ (.A1_N(_07905_),
    .A2_N(_07947_),
    .B1(\design_top.MEM[44][24] ),
    .B2(_07949_),
    .X(_06406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13749_ (.A(_07749_),
    .X(_07951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13750_ (.A(_07929_),
    .B(_07451_),
    .X(_07952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13751_ (.A(_07952_),
    .X(_07953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13752_ (.A1(_07846_),
    .A2(_07455_),
    .B1(_07952_),
    .X(_07954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13753_ (.A(_07954_),
    .X(_07955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13754_ (.A1_N(_07951_),
    .A2_N(_07953_),
    .B1(\design_top.MEM[45][15] ),
    .B2(_07955_),
    .X(_06405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13755_ (.A1_N(_07935_),
    .A2_N(_07953_),
    .B1(\design_top.MEM[45][14] ),
    .B2(_07955_),
    .X(_06404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13756_ (.A1_N(_07936_),
    .A2_N(_07953_),
    .B1(\design_top.MEM[45][13] ),
    .B2(_07955_),
    .X(_06403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13757_ (.A1_N(_07937_),
    .A2_N(_07953_),
    .B1(\design_top.MEM[45][12] ),
    .B2(_07955_),
    .X(_06402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13758_ (.A1_N(_07938_),
    .A2_N(_07953_),
    .B1(\design_top.MEM[45][11] ),
    .B2(_07955_),
    .X(_06401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13759_ (.A1_N(_07939_),
    .A2_N(_07952_),
    .B1(\design_top.MEM[45][10] ),
    .B2(_07954_),
    .X(_06400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13760_ (.A1_N(_07940_),
    .A2_N(_07952_),
    .B1(\design_top.MEM[45][9] ),
    .B2(_07954_),
    .X(_06399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13761_ (.A1_N(_07941_),
    .A2_N(_07952_),
    .B1(\design_top.MEM[45][8] ),
    .B2(_07954_),
    .X(_06398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13762_ (.A(_10783_),
    .B(_11276_),
    .X(_07956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13763_ (.A(_07894_),
    .B(_07956_),
    .X(_07957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13764_ (.A(_07957_),
    .X(_07958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13765_ (.A1(_11126_),
    .A2(_10992_),
    .B1(_07957_),
    .X(_07959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13766_ (.A(_07959_),
    .X(_07960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13767_ (.A1_N(_07893_),
    .A2_N(_07958_),
    .B1(\design_top.MEM[1][31] ),
    .B2(_07960_),
    .X(_06397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13768_ (.A1_N(_07899_),
    .A2_N(_07958_),
    .B1(\design_top.MEM[1][30] ),
    .B2(_07960_),
    .X(_06396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13769_ (.A1_N(_07900_),
    .A2_N(_07958_),
    .B1(\design_top.MEM[1][29] ),
    .B2(_07960_),
    .X(_06395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13770_ (.A1_N(_07901_),
    .A2_N(_07958_),
    .B1(\design_top.MEM[1][28] ),
    .B2(_07960_),
    .X(_06394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13771_ (.A1_N(_07902_),
    .A2_N(_07958_),
    .B1(\design_top.MEM[1][27] ),
    .B2(_07960_),
    .X(_06393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13772_ (.A1_N(_07903_),
    .A2_N(_07957_),
    .B1(\design_top.MEM[1][26] ),
    .B2(_07959_),
    .X(_06392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13773_ (.A1_N(_07904_),
    .A2_N(_07957_),
    .B1(\design_top.MEM[1][25] ),
    .B2(_07959_),
    .X(_06391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13774_ (.A1_N(_07905_),
    .A2_N(_07957_),
    .B1(\design_top.MEM[1][24] ),
    .B2(_07959_),
    .X(_06390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13775_ (.A(_07881_),
    .B(_07956_),
    .X(_07961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13776_ (.A(_07961_),
    .X(_07962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13777_ (.A1(_10792_),
    .A2(_10992_),
    .B1(_07961_),
    .X(_07963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13778_ (.A(_07963_),
    .X(_07964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13779_ (.A1_N(_07880_),
    .A2_N(_07962_),
    .B1(\design_top.MEM[1][23] ),
    .B2(_07964_),
    .X(_06389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13780_ (.A1_N(_07886_),
    .A2_N(_07962_),
    .B1(\design_top.MEM[1][22] ),
    .B2(_07964_),
    .X(_06388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13781_ (.A1_N(_07887_),
    .A2_N(_07962_),
    .B1(\design_top.MEM[1][21] ),
    .B2(_07964_),
    .X(_06387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13782_ (.A1_N(_07888_),
    .A2_N(_07962_),
    .B1(\design_top.MEM[1][20] ),
    .B2(_07964_),
    .X(_06386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13783_ (.A1_N(_07889_),
    .A2_N(_07962_),
    .B1(\design_top.MEM[1][19] ),
    .B2(_07964_),
    .X(_06385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13784_ (.A1_N(_07890_),
    .A2_N(_07961_),
    .B1(\design_top.MEM[1][18] ),
    .B2(_07963_),
    .X(_06384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13785_ (.A1_N(_07891_),
    .A2_N(_07961_),
    .B1(\design_top.MEM[1][17] ),
    .B2(_07963_),
    .X(_06383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13786_ (.A1_N(_07892_),
    .A2_N(_07961_),
    .B1(\design_top.MEM[1][16] ),
    .B2(_07963_),
    .X(_06382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13787_ (.A(_07929_),
    .B(_07956_),
    .X(_07965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13788_ (.A(_07965_),
    .X(_07966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13789_ (.A1(_10792_),
    .A2(_10992_),
    .B1(_07965_),
    .X(_07967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13790_ (.A(_07967_),
    .X(_07968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13791_ (.A1_N(_07951_),
    .A2_N(_07966_),
    .B1(\design_top.MEM[1][15] ),
    .B2(_07968_),
    .X(_06381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13792_ (.A1_N(_07935_),
    .A2_N(_07966_),
    .B1(\design_top.MEM[1][14] ),
    .B2(_07968_),
    .X(_06380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13793_ (.A1_N(_07936_),
    .A2_N(_07966_),
    .B1(\design_top.MEM[1][13] ),
    .B2(_07968_),
    .X(_06379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13794_ (.A1_N(_07937_),
    .A2_N(_07966_),
    .B1(\design_top.MEM[1][12] ),
    .B2(_07968_),
    .X(_06378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13795_ (.A1_N(_07938_),
    .A2_N(_07966_),
    .B1(\design_top.MEM[1][11] ),
    .B2(_07968_),
    .X(_06377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13796_ (.A1_N(_07939_),
    .A2_N(_07965_),
    .B1(\design_top.MEM[1][10] ),
    .B2(_07967_),
    .X(_06376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13797_ (.A1_N(_07940_),
    .A2_N(_07965_),
    .B1(\design_top.MEM[1][9] ),
    .B2(_07967_),
    .X(_06375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13798_ (.A1_N(_07941_),
    .A2_N(_07965_),
    .B1(\design_top.MEM[1][8] ),
    .B2(_07967_),
    .X(_06374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13799_ (.A(_07894_),
    .B(_07528_),
    .X(_07969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13800_ (.A(_07969_),
    .X(_07970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13801_ (.A1(_07913_),
    .A2(_07531_),
    .B1(_07969_),
    .X(_07971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13802_ (.A(_07971_),
    .X(_07972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13803_ (.A1_N(_07893_),
    .A2_N(_07970_),
    .B1(\design_top.MEM[22][31] ),
    .B2(_07972_),
    .X(_06373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13804_ (.A1_N(_07899_),
    .A2_N(_07970_),
    .B1(\design_top.MEM[22][30] ),
    .B2(_07972_),
    .X(_06372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13805_ (.A1_N(_07900_),
    .A2_N(_07970_),
    .B1(\design_top.MEM[22][29] ),
    .B2(_07972_),
    .X(_06371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13806_ (.A1_N(_07901_),
    .A2_N(_07970_),
    .B1(\design_top.MEM[22][28] ),
    .B2(_07972_),
    .X(_06370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13807_ (.A1_N(_07902_),
    .A2_N(_07970_),
    .B1(\design_top.MEM[22][27] ),
    .B2(_07972_),
    .X(_06369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13808_ (.A1_N(_07903_),
    .A2_N(_07969_),
    .B1(\design_top.MEM[22][26] ),
    .B2(_07971_),
    .X(_06368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13809_ (.A1_N(_07904_),
    .A2_N(_07969_),
    .B1(\design_top.MEM[22][25] ),
    .B2(_07971_),
    .X(_06367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13810_ (.A1_N(_07905_),
    .A2_N(_07969_),
    .B1(\design_top.MEM[22][24] ),
    .B2(_07971_),
    .X(_06366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13811_ (.A(_11039_),
    .B(_11255_),
    .X(_07973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13812_ (.A(_07929_),
    .B(_07973_),
    .X(_07974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13813_ (.A(_07974_),
    .X(_07975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13814_ (.A1(_07922_),
    .A2(_07531_),
    .B1(_07974_),
    .X(_07976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13815_ (.A(_07976_),
    .X(_07977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13816_ (.A1_N(_07951_),
    .A2_N(_07975_),
    .B1(\design_top.MEM[23][15] ),
    .B2(_07977_),
    .X(_06365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13817_ (.A1_N(_07935_),
    .A2_N(_07975_),
    .B1(\design_top.MEM[23][14] ),
    .B2(_07977_),
    .X(_06364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13818_ (.A1_N(_07936_),
    .A2_N(_07975_),
    .B1(\design_top.MEM[23][13] ),
    .B2(_07977_),
    .X(_06363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13819_ (.A1_N(_07937_),
    .A2_N(_07975_),
    .B1(\design_top.MEM[23][12] ),
    .B2(_07977_),
    .X(_06362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13820_ (.A1_N(_07938_),
    .A2_N(_07975_),
    .B1(\design_top.MEM[23][11] ),
    .B2(_07977_),
    .X(_06361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13821_ (.A1_N(_07939_),
    .A2_N(_07974_),
    .B1(\design_top.MEM[23][10] ),
    .B2(_07976_),
    .X(_06360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13822_ (.A1_N(_07940_),
    .A2_N(_07974_),
    .B1(\design_top.MEM[23][9] ),
    .B2(_07976_),
    .X(_06359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13823_ (.A1_N(_07941_),
    .A2_N(_07974_),
    .B1(\design_top.MEM[23][8] ),
    .B2(_07976_),
    .X(_06358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13824_ (.A(_10979_),
    .B(_11104_),
    .X(_07978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13825_ (.A(_07929_),
    .B(_07978_),
    .X(_07979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13826_ (.A(_07979_),
    .X(_07980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13827_ (.A1(_07846_),
    .A2(_07710_),
    .B1(_07979_),
    .X(_07981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13828_ (.A(_07981_),
    .X(_07982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13829_ (.A1_N(_07951_),
    .A2_N(_07980_),
    .B1(\design_top.MEM[37][15] ),
    .B2(_07982_),
    .X(_06357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13830_ (.A1_N(_07935_),
    .A2_N(_07980_),
    .B1(\design_top.MEM[37][14] ),
    .B2(_07982_),
    .X(_06356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13831_ (.A1_N(_07936_),
    .A2_N(_07980_),
    .B1(\design_top.MEM[37][13] ),
    .B2(_07982_),
    .X(_06355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13832_ (.A1_N(_07937_),
    .A2_N(_07980_),
    .B1(\design_top.MEM[37][12] ),
    .B2(_07982_),
    .X(_06354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13833_ (.A1_N(_07938_),
    .A2_N(_07980_),
    .B1(\design_top.MEM[37][11] ),
    .B2(_07982_),
    .X(_06353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13834_ (.A1_N(_07939_),
    .A2_N(_07979_),
    .B1(\design_top.MEM[37][10] ),
    .B2(_07981_),
    .X(_06352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13835_ (.A1_N(_07940_),
    .A2_N(_07979_),
    .B1(\design_top.MEM[37][9] ),
    .B2(_07981_),
    .X(_06351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13836_ (.A1_N(_07941_),
    .A2_N(_07979_),
    .B1(\design_top.MEM[37][8] ),
    .B2(_07981_),
    .X(_06350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13837_ (.A(_07639_),
    .X(_07983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13838_ (.A(_07641_),
    .X(_07984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13839_ (.A(_07984_),
    .B(_07973_),
    .X(_07985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13840_ (.A(_07985_),
    .X(_07986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13841_ (.A1(_07922_),
    .A2(_07531_),
    .B1(_07985_),
    .X(_07987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13842_ (.A(_07987_),
    .X(_07988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13843_ (.A1_N(_07983_),
    .A2_N(_07986_),
    .B1(\design_top.MEM[23][23] ),
    .B2(_07988_),
    .X(_06349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13844_ (.A(_07648_),
    .X(_07989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13845_ (.A1_N(_07989_),
    .A2_N(_07986_),
    .B1(\design_top.MEM[23][22] ),
    .B2(_07988_),
    .X(_06348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13846_ (.A(_07650_),
    .X(_07990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13847_ (.A1_N(_07990_),
    .A2_N(_07986_),
    .B1(\design_top.MEM[23][21] ),
    .B2(_07988_),
    .X(_06347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13848_ (.A(_07652_),
    .X(_07991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13849_ (.A1_N(_07991_),
    .A2_N(_07986_),
    .B1(\design_top.MEM[23][20] ),
    .B2(_07988_),
    .X(_06346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13850_ (.A(_07654_),
    .X(_07992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13851_ (.A1_N(_07992_),
    .A2_N(_07986_),
    .B1(\design_top.MEM[23][19] ),
    .B2(_07988_),
    .X(_06345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13852_ (.A(_07656_),
    .X(_07993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13853_ (.A1_N(_07993_),
    .A2_N(_07985_),
    .B1(\design_top.MEM[23][18] ),
    .B2(_07987_),
    .X(_06344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13854_ (.A(_07658_),
    .X(_07994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13855_ (.A1_N(_07994_),
    .A2_N(_07985_),
    .B1(\design_top.MEM[23][17] ),
    .B2(_07987_),
    .X(_06343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13856_ (.A(_07660_),
    .X(_07995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13857_ (.A1_N(_07995_),
    .A2_N(_07985_),
    .B1(\design_top.MEM[23][16] ),
    .B2(_07987_),
    .X(_06342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13858_ (.A(_07984_),
    .B(_07978_),
    .X(_07996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13859_ (.A(_07996_),
    .X(_07997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13860_ (.A(_07508_),
    .X(_07998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13861_ (.A1(_07998_),
    .A2(_07710_),
    .B1(_07996_),
    .X(_07999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13862_ (.A(_07999_),
    .X(_08000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13863_ (.A1_N(_07983_),
    .A2_N(_07997_),
    .B1(\design_top.MEM[37][23] ),
    .B2(_08000_),
    .X(_06341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13864_ (.A1_N(_07989_),
    .A2_N(_07997_),
    .B1(\design_top.MEM[37][22] ),
    .B2(_08000_),
    .X(_06340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13865_ (.A1_N(_07990_),
    .A2_N(_07997_),
    .B1(\design_top.MEM[37][21] ),
    .B2(_08000_),
    .X(_06339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13866_ (.A1_N(_07991_),
    .A2_N(_07997_),
    .B1(\design_top.MEM[37][20] ),
    .B2(_08000_),
    .X(_06338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13867_ (.A1_N(_07992_),
    .A2_N(_07997_),
    .B1(\design_top.MEM[37][19] ),
    .B2(_08000_),
    .X(_06337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13868_ (.A1_N(_07993_),
    .A2_N(_07996_),
    .B1(\design_top.MEM[37][18] ),
    .B2(_07999_),
    .X(_06336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13869_ (.A1_N(_07994_),
    .A2_N(_07996_),
    .B1(\design_top.MEM[37][17] ),
    .B2(_07999_),
    .X(_06335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13870_ (.A1_N(_07995_),
    .A2_N(_07996_),
    .B1(\design_top.MEM[37][16] ),
    .B2(_07999_),
    .X(_06334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13871_ (.A(_07676_),
    .X(_08001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13872_ (.A(_07678_),
    .X(_08002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13873_ (.A(_08002_),
    .B(_07978_),
    .X(_08003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13874_ (.A(_08003_),
    .X(_08004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13875_ (.A1(_07998_),
    .A2(_07710_),
    .B1(_08003_),
    .X(_08005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13876_ (.A(_08005_),
    .X(_08006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13877_ (.A1_N(_08001_),
    .A2_N(_08004_),
    .B1(\design_top.MEM[37][31] ),
    .B2(_08006_),
    .X(_06333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13878_ (.A(_07684_),
    .X(_08007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13879_ (.A1_N(_08007_),
    .A2_N(_08004_),
    .B1(\design_top.MEM[37][30] ),
    .B2(_08006_),
    .X(_06332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13880_ (.A(_07686_),
    .X(_08008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13881_ (.A1_N(_08008_),
    .A2_N(_08004_),
    .B1(\design_top.MEM[37][29] ),
    .B2(_08006_),
    .X(_06331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13882_ (.A(_07688_),
    .X(_08009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13883_ (.A1_N(_08009_),
    .A2_N(_08004_),
    .B1(\design_top.MEM[37][28] ),
    .B2(_08006_),
    .X(_06330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13884_ (.A(_07690_),
    .X(_08010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13885_ (.A1_N(_08010_),
    .A2_N(_08004_),
    .B1(\design_top.MEM[37][27] ),
    .B2(_08006_),
    .X(_06329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13886_ (.A(_07692_),
    .X(_08011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13887_ (.A1_N(_08011_),
    .A2_N(_08003_),
    .B1(\design_top.MEM[37][26] ),
    .B2(_08005_),
    .X(_06328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13888_ (.A(_07694_),
    .X(_08012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13889_ (.A1_N(_08012_),
    .A2_N(_08003_),
    .B1(\design_top.MEM[37][25] ),
    .B2(_08005_),
    .X(_06327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13890_ (.A(_07696_),
    .X(_08013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13891_ (.A1_N(_08013_),
    .A2_N(_08003_),
    .B1(\design_top.MEM[37][24] ),
    .B2(_08005_),
    .X(_06326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13892_ (.A(_08002_),
    .B(_07973_),
    .X(_08014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13893_ (.A(_08014_),
    .X(_08015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13894_ (.A1(_07922_),
    .A2(_07476_),
    .B1(_08014_),
    .X(_08016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13895_ (.A(_08016_),
    .X(_08017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13896_ (.A1_N(_08001_),
    .A2_N(_08015_),
    .B1(\design_top.MEM[23][31] ),
    .B2(_08017_),
    .X(_06325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13897_ (.A1_N(_08007_),
    .A2_N(_08015_),
    .B1(\design_top.MEM[23][30] ),
    .B2(_08017_),
    .X(_06324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13898_ (.A1_N(_08008_),
    .A2_N(_08015_),
    .B1(\design_top.MEM[23][29] ),
    .B2(_08017_),
    .X(_06323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13899_ (.A1_N(_08009_),
    .A2_N(_08015_),
    .B1(\design_top.MEM[23][28] ),
    .B2(_08017_),
    .X(_06322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13900_ (.A1_N(_08010_),
    .A2_N(_08015_),
    .B1(\design_top.MEM[23][27] ),
    .B2(_08017_),
    .X(_06321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13901_ (.A1_N(_08011_),
    .A2_N(_08014_),
    .B1(\design_top.MEM[23][26] ),
    .B2(_08016_),
    .X(_06320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13902_ (.A1_N(_08012_),
    .A2_N(_08014_),
    .B1(\design_top.MEM[23][25] ),
    .B2(_08016_),
    .X(_06319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13903_ (.A1_N(_08013_),
    .A2_N(_08014_),
    .B1(\design_top.MEM[23][24] ),
    .B2(_08016_),
    .X(_06318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13904_ (.A(_07726_),
    .X(_08018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13905_ (.A(_11102_),
    .B(_10956_),
    .X(_08019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13906_ (.A(_08018_),
    .B(_08019_),
    .X(_08020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13907_ (.A(_08020_),
    .X(_08021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13908_ (.A1(_07944_),
    .A2(_10899_),
    .B1(_08020_),
    .X(_08022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13909_ (.A(_08022_),
    .X(_08023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13910_ (.A1_N(_07951_),
    .A2_N(_08021_),
    .B1(\design_top.MEM[24][15] ),
    .B2(_08023_),
    .X(_06317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13911_ (.A(_07735_),
    .X(_08024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13912_ (.A1_N(_08024_),
    .A2_N(_08021_),
    .B1(\design_top.MEM[24][14] ),
    .B2(_08023_),
    .X(_06316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13913_ (.A(_07737_),
    .X(_08025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13914_ (.A1_N(_08025_),
    .A2_N(_08021_),
    .B1(\design_top.MEM[24][13] ),
    .B2(_08023_),
    .X(_06315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13915_ (.A(_07739_),
    .X(_08026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13916_ (.A1_N(_08026_),
    .A2_N(_08021_),
    .B1(\design_top.MEM[24][12] ),
    .B2(_08023_),
    .X(_06314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13917_ (.A(_07741_),
    .X(_08027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13918_ (.A1_N(_08027_),
    .A2_N(_08021_),
    .B1(\design_top.MEM[24][11] ),
    .B2(_08023_),
    .X(_06313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13919_ (.A(_07743_),
    .X(_08028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13920_ (.A1_N(_08028_),
    .A2_N(_08020_),
    .B1(\design_top.MEM[24][10] ),
    .B2(_08022_),
    .X(_06312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13921_ (.A(_07745_),
    .X(_08029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13922_ (.A1_N(_08029_),
    .A2_N(_08020_),
    .B1(\design_top.MEM[24][9] ),
    .B2(_08022_),
    .X(_06311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13923_ (.A(_07747_),
    .X(_08030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13924_ (.A1_N(_08030_),
    .A2_N(_08020_),
    .B1(\design_top.MEM[24][8] ),
    .B2(_08022_),
    .X(_06310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13925_ (.A(_07749_),
    .X(_08031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13926_ (.A(_08018_),
    .B(_07671_),
    .X(_08032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13927_ (.A(_08032_),
    .X(_08033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13928_ (.A1(_07913_),
    .A2(_07520_),
    .B1(_08032_),
    .X(_08034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13929_ (.A(_08034_),
    .X(_08035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13930_ (.A1_N(_08031_),
    .A2_N(_08033_),
    .B1(\design_top.MEM[38][15] ),
    .B2(_08035_),
    .X(_06309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13931_ (.A1_N(_08024_),
    .A2_N(_08033_),
    .B1(\design_top.MEM[38][14] ),
    .B2(_08035_),
    .X(_06308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13932_ (.A1_N(_08025_),
    .A2_N(_08033_),
    .B1(\design_top.MEM[38][13] ),
    .B2(_08035_),
    .X(_06307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13933_ (.A1_N(_08026_),
    .A2_N(_08033_),
    .B1(\design_top.MEM[38][12] ),
    .B2(_08035_),
    .X(_06306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13934_ (.A1_N(_08027_),
    .A2_N(_08033_),
    .B1(\design_top.MEM[38][11] ),
    .B2(_08035_),
    .X(_06305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13935_ (.A1_N(_08028_),
    .A2_N(_08032_),
    .B1(\design_top.MEM[38][10] ),
    .B2(_08034_),
    .X(_06304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13936_ (.A1_N(_08029_),
    .A2_N(_08032_),
    .B1(\design_top.MEM[38][9] ),
    .B2(_08034_),
    .X(_06303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13937_ (.A1_N(_08030_),
    .A2_N(_08032_),
    .B1(\design_top.MEM[38][8] ),
    .B2(_08034_),
    .X(_06302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13938_ (.A(_07984_),
    .B(_08019_),
    .X(_08036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13939_ (.A(_08036_),
    .X(_08037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13940_ (.A1(_07944_),
    .A2(_10899_),
    .B1(_08036_),
    .X(_08038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13941_ (.A(_08038_),
    .X(_08039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13942_ (.A1_N(_07983_),
    .A2_N(_08037_),
    .B1(\design_top.MEM[24][23] ),
    .B2(_08039_),
    .X(_06301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13943_ (.A1_N(_07989_),
    .A2_N(_08037_),
    .B1(\design_top.MEM[24][22] ),
    .B2(_08039_),
    .X(_06300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13944_ (.A1_N(_07990_),
    .A2_N(_08037_),
    .B1(\design_top.MEM[24][21] ),
    .B2(_08039_),
    .X(_06299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13945_ (.A1_N(_07991_),
    .A2_N(_08037_),
    .B1(\design_top.MEM[24][20] ),
    .B2(_08039_),
    .X(_06298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13946_ (.A1_N(_07992_),
    .A2_N(_08037_),
    .B1(\design_top.MEM[24][19] ),
    .B2(_08039_),
    .X(_06297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13947_ (.A1_N(_07993_),
    .A2_N(_08036_),
    .B1(\design_top.MEM[24][18] ),
    .B2(_08038_),
    .X(_06296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13948_ (.A1_N(_07994_),
    .A2_N(_08036_),
    .B1(\design_top.MEM[24][17] ),
    .B2(_08038_),
    .X(_06295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13949_ (.A1_N(_07995_),
    .A2_N(_08036_),
    .B1(\design_top.MEM[24][16] ),
    .B2(_08038_),
    .X(_06294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13950_ (.A(_08002_),
    .B(_08019_),
    .X(_08040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13951_ (.A(_08040_),
    .X(_08041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13952_ (.A1(_07944_),
    .A2(_10898_),
    .B1(_08040_),
    .X(_08042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13953_ (.A(_08042_),
    .X(_08043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13954_ (.A1_N(_08001_),
    .A2_N(_08041_),
    .B1(\design_top.MEM[24][31] ),
    .B2(_08043_),
    .X(_06293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13955_ (.A1_N(_08007_),
    .A2_N(_08041_),
    .B1(\design_top.MEM[24][30] ),
    .B2(_08043_),
    .X(_06292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13956_ (.A1_N(_08008_),
    .A2_N(_08041_),
    .B1(\design_top.MEM[24][29] ),
    .B2(_08043_),
    .X(_06291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13957_ (.A1_N(_08009_),
    .A2_N(_08041_),
    .B1(\design_top.MEM[24][28] ),
    .B2(_08043_),
    .X(_06290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13958_ (.A1_N(_08010_),
    .A2_N(_08041_),
    .B1(\design_top.MEM[24][27] ),
    .B2(_08043_),
    .X(_06289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13959_ (.A1_N(_08011_),
    .A2_N(_08040_),
    .B1(\design_top.MEM[24][26] ),
    .B2(_08042_),
    .X(_06288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13960_ (.A1_N(_08012_),
    .A2_N(_08040_),
    .B1(\design_top.MEM[24][25] ),
    .B2(_08042_),
    .X(_06287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13961_ (.A1_N(_08013_),
    .A2_N(_08040_),
    .B1(\design_top.MEM[24][24] ),
    .B2(_08042_),
    .X(_06286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13962_ (.A(_10881_),
    .B(_11276_),
    .X(_08044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13963_ (.A(_08018_),
    .B(_08044_),
    .X(_08045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13964_ (.A(_08045_),
    .X(_08046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13965_ (.A(_10898_),
    .X(_08047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13966_ (.A1(_08047_),
    .A2(_11196_),
    .B1(_08045_),
    .X(_08048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13967_ (.A(_08048_),
    .X(_08049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13968_ (.A1_N(_08031_),
    .A2_N(_08046_),
    .B1(\design_top.MEM[25][15] ),
    .B2(_08049_),
    .X(_06285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13969_ (.A1_N(_08024_),
    .A2_N(_08046_),
    .B1(\design_top.MEM[25][14] ),
    .B2(_08049_),
    .X(_06284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13970_ (.A1_N(_08025_),
    .A2_N(_08046_),
    .B1(\design_top.MEM[25][13] ),
    .B2(_08049_),
    .X(_06283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13971_ (.A1_N(_08026_),
    .A2_N(_08046_),
    .B1(\design_top.MEM[25][12] ),
    .B2(_08049_),
    .X(_06282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13972_ (.A1_N(_08027_),
    .A2_N(_08046_),
    .B1(\design_top.MEM[25][11] ),
    .B2(_08049_),
    .X(_06281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13973_ (.A1_N(_08028_),
    .A2_N(_08045_),
    .B1(\design_top.MEM[25][10] ),
    .B2(_08048_),
    .X(_06280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13974_ (.A1_N(_08029_),
    .A2_N(_08045_),
    .B1(\design_top.MEM[25][9] ),
    .B2(_08048_),
    .X(_06279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13975_ (.A1_N(_08030_),
    .A2_N(_08045_),
    .B1(\design_top.MEM[25][8] ),
    .B2(_08048_),
    .X(_06278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13976_ (.A(_07984_),
    .B(_07671_),
    .X(_08050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13977_ (.A(_08050_),
    .X(_08051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13978_ (.A1(_07913_),
    .A2(_07520_),
    .B1(_08050_),
    .X(_08052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13979_ (.A(_08052_),
    .X(_08053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13980_ (.A1_N(_07983_),
    .A2_N(_08051_),
    .B1(\design_top.MEM[38][23] ),
    .B2(_08053_),
    .X(_06277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13981_ (.A1_N(_07989_),
    .A2_N(_08051_),
    .B1(\design_top.MEM[38][22] ),
    .B2(_08053_),
    .X(_06276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13982_ (.A1_N(_07990_),
    .A2_N(_08051_),
    .B1(\design_top.MEM[38][21] ),
    .B2(_08053_),
    .X(_06275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13983_ (.A1_N(_07991_),
    .A2_N(_08051_),
    .B1(\design_top.MEM[38][20] ),
    .B2(_08053_),
    .X(_06274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13984_ (.A1_N(_07992_),
    .A2_N(_08051_),
    .B1(\design_top.MEM[38][19] ),
    .B2(_08053_),
    .X(_06273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13985_ (.A1_N(_07993_),
    .A2_N(_08050_),
    .B1(\design_top.MEM[38][18] ),
    .B2(_08052_),
    .X(_06272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13986_ (.A1_N(_07994_),
    .A2_N(_08050_),
    .B1(\design_top.MEM[38][17] ),
    .B2(_08052_),
    .X(_06271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13987_ (.A1_N(_07995_),
    .A2_N(_08050_),
    .B1(\design_top.MEM[38][16] ),
    .B2(_08052_),
    .X(_06270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13988_ (.A(_08002_),
    .B(_07472_),
    .X(_08054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13989_ (.A(_08054_),
    .X(_08055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13990_ (.A(_10797_),
    .X(_08056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13991_ (.A(_08056_),
    .X(_08057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13992_ (.A1(_08057_),
    .A2(_07476_),
    .B1(_08054_),
    .X(_08058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13993_ (.A(_08058_),
    .X(_08059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13994_ (.A1_N(_08001_),
    .A2_N(_08055_),
    .B1(\design_top.MEM[20][31] ),
    .B2(_08059_),
    .X(_06269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13995_ (.A1_N(_08007_),
    .A2_N(_08055_),
    .B1(\design_top.MEM[20][30] ),
    .B2(_08059_),
    .X(_06268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13996_ (.A1_N(_08008_),
    .A2_N(_08055_),
    .B1(\design_top.MEM[20][29] ),
    .B2(_08059_),
    .X(_06267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13997_ (.A1_N(_08009_),
    .A2_N(_08055_),
    .B1(\design_top.MEM[20][28] ),
    .B2(_08059_),
    .X(_06266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13998_ (.A1_N(_08010_),
    .A2_N(_08055_),
    .B1(\design_top.MEM[20][27] ),
    .B2(_08059_),
    .X(_06265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13999_ (.A1_N(_08011_),
    .A2_N(_08054_),
    .B1(\design_top.MEM[20][26] ),
    .B2(_08058_),
    .X(_06264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14000_ (.A1_N(_08012_),
    .A2_N(_08054_),
    .B1(\design_top.MEM[20][25] ),
    .B2(_08058_),
    .X(_06263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14001_ (.A1_N(_08013_),
    .A2_N(_08054_),
    .B1(\design_top.MEM[20][24] ),
    .B2(_08058_),
    .X(_06262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14002_ (.A(_07984_),
    .B(_08044_),
    .X(_08060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14003_ (.A(_08060_),
    .X(_08061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14004_ (.A1(_08047_),
    .A2(_11196_),
    .B1(_08060_),
    .X(_08062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14005_ (.A(_08062_),
    .X(_08063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14006_ (.A1_N(_07983_),
    .A2_N(_08061_),
    .B1(\design_top.MEM[25][23] ),
    .B2(_08063_),
    .X(_06261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14007_ (.A1_N(_07989_),
    .A2_N(_08061_),
    .B1(\design_top.MEM[25][22] ),
    .B2(_08063_),
    .X(_06260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14008_ (.A1_N(_07990_),
    .A2_N(_08061_),
    .B1(\design_top.MEM[25][21] ),
    .B2(_08063_),
    .X(_06259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14009_ (.A1_N(_07991_),
    .A2_N(_08061_),
    .B1(\design_top.MEM[25][20] ),
    .B2(_08063_),
    .X(_06258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14010_ (.A1_N(_07992_),
    .A2_N(_08061_),
    .B1(\design_top.MEM[25][19] ),
    .B2(_08063_),
    .X(_06257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14011_ (.A1_N(_07993_),
    .A2_N(_08060_),
    .B1(\design_top.MEM[25][18] ),
    .B2(_08062_),
    .X(_06256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14012_ (.A1_N(_07994_),
    .A2_N(_08060_),
    .B1(\design_top.MEM[25][17] ),
    .B2(_08062_),
    .X(_06255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14013_ (.A1_N(_07995_),
    .A2_N(_08060_),
    .B1(\design_top.MEM[25][16] ),
    .B2(_08062_),
    .X(_06254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14014_ (.A(_08002_),
    .B(_08044_),
    .X(_08064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14015_ (.A(_08064_),
    .X(_08065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14016_ (.A1(_08047_),
    .A2(_11196_),
    .B1(_08064_),
    .X(_08066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14017_ (.A(_08066_),
    .X(_08067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14018_ (.A1_N(_08001_),
    .A2_N(_08065_),
    .B1(\design_top.MEM[25][31] ),
    .B2(_08067_),
    .X(_06253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14019_ (.A1_N(_08007_),
    .A2_N(_08065_),
    .B1(\design_top.MEM[25][30] ),
    .B2(_08067_),
    .X(_06252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14020_ (.A1_N(_08008_),
    .A2_N(_08065_),
    .B1(\design_top.MEM[25][29] ),
    .B2(_08067_),
    .X(_06251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14021_ (.A1_N(_08009_),
    .A2_N(_08065_),
    .B1(\design_top.MEM[25][28] ),
    .B2(_08067_),
    .X(_06250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14022_ (.A1_N(_08010_),
    .A2_N(_08065_),
    .B1(\design_top.MEM[25][27] ),
    .B2(_08067_),
    .X(_06249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14023_ (.A1_N(_08011_),
    .A2_N(_08064_),
    .B1(\design_top.MEM[25][26] ),
    .B2(_08066_),
    .X(_06248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14024_ (.A1_N(_08012_),
    .A2_N(_08064_),
    .B1(\design_top.MEM[25][25] ),
    .B2(_08066_),
    .X(_06247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14025_ (.A1_N(_08013_),
    .A2_N(_08064_),
    .B1(\design_top.MEM[25][24] ),
    .B2(_08066_),
    .X(_06246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14026_ (.A(_10881_),
    .B(_11000_),
    .X(_08068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14027_ (.A(_08018_),
    .B(_08068_),
    .X(_08069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14028_ (.A(_08069_),
    .X(_08070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14029_ (.A1(_08047_),
    .A2(_11135_),
    .B1(_08069_),
    .X(_08071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14030_ (.A(_08071_),
    .X(_08072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14031_ (.A1_N(_08031_),
    .A2_N(_08070_),
    .B1(\design_top.MEM[26][15] ),
    .B2(_08072_),
    .X(_06245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14032_ (.A1_N(_08024_),
    .A2_N(_08070_),
    .B1(\design_top.MEM[26][14] ),
    .B2(_08072_),
    .X(_06244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14033_ (.A1_N(_08025_),
    .A2_N(_08070_),
    .B1(\design_top.MEM[26][13] ),
    .B2(_08072_),
    .X(_06243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14034_ (.A1_N(_08026_),
    .A2_N(_08070_),
    .B1(\design_top.MEM[26][12] ),
    .B2(_08072_),
    .X(_06242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14035_ (.A1_N(_08027_),
    .A2_N(_08070_),
    .B1(\design_top.MEM[26][11] ),
    .B2(_08072_),
    .X(_06241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14036_ (.A1_N(_08028_),
    .A2_N(_08069_),
    .B1(\design_top.MEM[26][10] ),
    .B2(_08071_),
    .X(_06240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14037_ (.A1_N(_08029_),
    .A2_N(_08069_),
    .B1(\design_top.MEM[26][9] ),
    .B2(_08071_),
    .X(_06239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14038_ (.A1_N(_08030_),
    .A2_N(_08069_),
    .B1(\design_top.MEM[26][8] ),
    .B2(_08071_),
    .X(_06238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14039_ (.A(_07639_),
    .X(_08073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14040_ (.A(_07641_),
    .X(_08074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14041_ (.A(_08074_),
    .B(_08068_),
    .X(_08075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14042_ (.A(_08075_),
    .X(_08076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14043_ (.A1(_08047_),
    .A2(_11135_),
    .B1(_08075_),
    .X(_08077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14044_ (.A(_08077_),
    .X(_08078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14045_ (.A1_N(_08073_),
    .A2_N(_08076_),
    .B1(\design_top.MEM[26][23] ),
    .B2(_08078_),
    .X(_06237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14046_ (.A(_07648_),
    .X(_08079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14047_ (.A1_N(_08079_),
    .A2_N(_08076_),
    .B1(\design_top.MEM[26][22] ),
    .B2(_08078_),
    .X(_06236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14048_ (.A(_07650_),
    .X(_08080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14049_ (.A1_N(_08080_),
    .A2_N(_08076_),
    .B1(\design_top.MEM[26][21] ),
    .B2(_08078_),
    .X(_06235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14050_ (.A(_07652_),
    .X(_08081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14051_ (.A1_N(_08081_),
    .A2_N(_08076_),
    .B1(\design_top.MEM[26][20] ),
    .B2(_08078_),
    .X(_06234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14052_ (.A(_07654_),
    .X(_08082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14053_ (.A1_N(_08082_),
    .A2_N(_08076_),
    .B1(\design_top.MEM[26][19] ),
    .B2(_08078_),
    .X(_06233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14054_ (.A(_07656_),
    .X(_08083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14055_ (.A1_N(_08083_),
    .A2_N(_08075_),
    .B1(\design_top.MEM[26][18] ),
    .B2(_08077_),
    .X(_06232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14056_ (.A(_07658_),
    .X(_08084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14057_ (.A1_N(_08084_),
    .A2_N(_08075_),
    .B1(\design_top.MEM[26][17] ),
    .B2(_08077_),
    .X(_06231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14058_ (.A(_07660_),
    .X(_08085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14059_ (.A1_N(_08085_),
    .A2_N(_08075_),
    .B1(\design_top.MEM[26][16] ),
    .B2(_08077_),
    .X(_06230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14060_ (.A(_07676_),
    .X(_08086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14061_ (.A(_07678_),
    .X(_08087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14062_ (.A(_08087_),
    .B(_08068_),
    .X(_08088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14063_ (.A(_08088_),
    .X(_08089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14064_ (.A1(_10899_),
    .A2(_11135_),
    .B1(_08088_),
    .X(_08090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14065_ (.A(_08090_),
    .X(_08091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14066_ (.A1_N(_08086_),
    .A2_N(_08089_),
    .B1(\design_top.MEM[26][31] ),
    .B2(_08091_),
    .X(_06229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14067_ (.A(_07684_),
    .X(_08092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14068_ (.A1_N(_08092_),
    .A2_N(_08089_),
    .B1(\design_top.MEM[26][30] ),
    .B2(_08091_),
    .X(_06228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14069_ (.A(_07686_),
    .X(_08093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14070_ (.A1_N(_08093_),
    .A2_N(_08089_),
    .B1(\design_top.MEM[26][29] ),
    .B2(_08091_),
    .X(_06227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14071_ (.A(_07688_),
    .X(_08094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14072_ (.A1_N(_08094_),
    .A2_N(_08089_),
    .B1(\design_top.MEM[26][28] ),
    .B2(_08091_),
    .X(_06226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14073_ (.A(_07690_),
    .X(_08095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14074_ (.A1_N(_08095_),
    .A2_N(_08089_),
    .B1(\design_top.MEM[26][27] ),
    .B2(_08091_),
    .X(_06225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14075_ (.A(_07692_),
    .X(_08096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14076_ (.A1_N(_08096_),
    .A2_N(_08088_),
    .B1(\design_top.MEM[26][26] ),
    .B2(_08090_),
    .X(_06224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14077_ (.A(_07694_),
    .X(_08097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14078_ (.A1_N(_08097_),
    .A2_N(_08088_),
    .B1(\design_top.MEM[26][25] ),
    .B2(_08090_),
    .X(_06223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14079_ (.A(_07696_),
    .X(_08098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14080_ (.A1_N(_08098_),
    .A2_N(_08088_),
    .B1(\design_top.MEM[26][24] ),
    .B2(_08090_),
    .X(_06222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14081_ (.A(_08018_),
    .B(_10886_),
    .X(_08099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14082_ (.A(_08099_),
    .X(_08100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14083_ (.A1(_07922_),
    .A2(_10898_),
    .B1(_08099_),
    .X(_08101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14084_ (.A(_08101_),
    .X(_08102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14085_ (.A1_N(_08031_),
    .A2_N(_08100_),
    .B1(\design_top.MEM[27][15] ),
    .B2(_08102_),
    .X(_06221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14086_ (.A1_N(_08024_),
    .A2_N(_08100_),
    .B1(\design_top.MEM[27][14] ),
    .B2(_08102_),
    .X(_06220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14087_ (.A1_N(_08025_),
    .A2_N(_08100_),
    .B1(\design_top.MEM[27][13] ),
    .B2(_08102_),
    .X(_06219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14088_ (.A1_N(_08026_),
    .A2_N(_08100_),
    .B1(\design_top.MEM[27][12] ),
    .B2(_08102_),
    .X(_06218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14089_ (.A1_N(_08027_),
    .A2_N(_08100_),
    .B1(\design_top.MEM[27][11] ),
    .B2(_08102_),
    .X(_06217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14090_ (.A1_N(_08028_),
    .A2_N(_08099_),
    .B1(\design_top.MEM[27][10] ),
    .B2(_08101_),
    .X(_06216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14091_ (.A1_N(_08029_),
    .A2_N(_08099_),
    .B1(\design_top.MEM[27][9] ),
    .B2(_08101_),
    .X(_06215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14092_ (.A1_N(_08030_),
    .A2_N(_08099_),
    .B1(\design_top.MEM[27][8] ),
    .B2(_08101_),
    .X(_06214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14093_ (.A(_11129_),
    .B(_11276_),
    .X(_08103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14094_ (.A(_08074_),
    .B(_08103_),
    .X(_08104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14095_ (.A(_08104_),
    .X(_08105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14096_ (.A1(_07998_),
    .A2(_11162_),
    .B1(_08104_),
    .X(_08106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14097_ (.A(_08106_),
    .X(_08107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14098_ (.A1_N(_08073_),
    .A2_N(_08105_),
    .B1(\design_top.MEM[9][23] ),
    .B2(_08107_),
    .X(_06213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14099_ (.A1_N(_08079_),
    .A2_N(_08105_),
    .B1(\design_top.MEM[9][22] ),
    .B2(_08107_),
    .X(_06212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14100_ (.A1_N(_08080_),
    .A2_N(_08105_),
    .B1(\design_top.MEM[9][21] ),
    .B2(_08107_),
    .X(_06211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14101_ (.A1_N(_08081_),
    .A2_N(_08105_),
    .B1(\design_top.MEM[9][20] ),
    .B2(_08107_),
    .X(_06210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14102_ (.A1_N(_08082_),
    .A2_N(_08105_),
    .B1(\design_top.MEM[9][19] ),
    .B2(_08107_),
    .X(_06209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14103_ (.A1_N(_08083_),
    .A2_N(_08104_),
    .B1(\design_top.MEM[9][18] ),
    .B2(_08106_),
    .X(_06208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14104_ (.A1_N(_08084_),
    .A2_N(_08104_),
    .B1(\design_top.MEM[9][17] ),
    .B2(_08106_),
    .X(_06207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14105_ (.A1_N(_08085_),
    .A2_N(_08104_),
    .B1(\design_top.MEM[9][16] ),
    .B2(_08106_),
    .X(_06206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14106_ (.A(_07726_),
    .X(_08108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14107_ (.A(_08108_),
    .B(_08103_),
    .X(_08109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14108_ (.A(_08109_),
    .X(_08110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14109_ (.A1(_07998_),
    .A2(_11162_),
    .B1(_08109_),
    .X(_08111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14110_ (.A(_08111_),
    .X(_08112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14111_ (.A1_N(_08031_),
    .A2_N(_08110_),
    .B1(\design_top.MEM[9][15] ),
    .B2(_08112_),
    .X(_06205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14112_ (.A(_07735_),
    .X(_08113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14113_ (.A1_N(_08113_),
    .A2_N(_08110_),
    .B1(\design_top.MEM[9][14] ),
    .B2(_08112_),
    .X(_06204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14114_ (.A(_07737_),
    .X(_08114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14115_ (.A1_N(_08114_),
    .A2_N(_08110_),
    .B1(\design_top.MEM[9][13] ),
    .B2(_08112_),
    .X(_06203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14116_ (.A(_07739_),
    .X(_08115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14117_ (.A1_N(_08115_),
    .A2_N(_08110_),
    .B1(\design_top.MEM[9][12] ),
    .B2(_08112_),
    .X(_06202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14118_ (.A(_07741_),
    .X(_08116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14119_ (.A1_N(_08116_),
    .A2_N(_08110_),
    .B1(\design_top.MEM[9][11] ),
    .B2(_08112_),
    .X(_06201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14120_ (.A(_07743_),
    .X(_08117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14121_ (.A1_N(_08117_),
    .A2_N(_08109_),
    .B1(\design_top.MEM[9][10] ),
    .B2(_08111_),
    .X(_06200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14122_ (.A(_07745_),
    .X(_08118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14123_ (.A1_N(_08118_),
    .A2_N(_08109_),
    .B1(\design_top.MEM[9][9] ),
    .B2(_08111_),
    .X(_06199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14124_ (.A(_07747_),
    .X(_08119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14125_ (.A1_N(_08119_),
    .A2_N(_08109_),
    .B1(\design_top.MEM[9][8] ),
    .B2(_08111_),
    .X(_06198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14126_ (.A(_10776_),
    .B(_11129_),
    .X(_08120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14127_ (.A(_08087_),
    .B(_08120_),
    .X(_08121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14128_ (.A(_08121_),
    .X(_08122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14129_ (.A1(_08057_),
    .A2(_11162_),
    .B1(_08121_),
    .X(_08123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14130_ (.A(_08123_),
    .X(_08124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14131_ (.A1_N(_08086_),
    .A2_N(_08122_),
    .B1(\design_top.MEM[8][31] ),
    .B2(_08124_),
    .X(_06197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14132_ (.A1_N(_08092_),
    .A2_N(_08122_),
    .B1(\design_top.MEM[8][30] ),
    .B2(_08124_),
    .X(_06196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14133_ (.A1_N(_08093_),
    .A2_N(_08122_),
    .B1(\design_top.MEM[8][29] ),
    .B2(_08124_),
    .X(_06195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14134_ (.A1_N(_08094_),
    .A2_N(_08122_),
    .B1(\design_top.MEM[8][28] ),
    .B2(_08124_),
    .X(_06194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14135_ (.A1_N(_08095_),
    .A2_N(_08122_),
    .B1(\design_top.MEM[8][27] ),
    .B2(_08124_),
    .X(_06193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14136_ (.A1_N(_08096_),
    .A2_N(_08121_),
    .B1(\design_top.MEM[8][26] ),
    .B2(_08123_),
    .X(_06192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14137_ (.A1_N(_08097_),
    .A2_N(_08121_),
    .B1(\design_top.MEM[8][25] ),
    .B2(_08123_),
    .X(_06191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14138_ (.A1_N(_08098_),
    .A2_N(_08121_),
    .B1(\design_top.MEM[8][24] ),
    .B2(_08123_),
    .X(_06190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14139_ (.A(_08074_),
    .B(_08120_),
    .X(_08125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14140_ (.A(_08125_),
    .X(_08126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14141_ (.A1(_08057_),
    .A2(_11162_),
    .B1(_08125_),
    .X(_08127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14142_ (.A(_08127_),
    .X(_08128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14143_ (.A1_N(_08073_),
    .A2_N(_08126_),
    .B1(\design_top.MEM[8][23] ),
    .B2(_08128_),
    .X(_06189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14144_ (.A1_N(_08079_),
    .A2_N(_08126_),
    .B1(\design_top.MEM[8][22] ),
    .B2(_08128_),
    .X(_06188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14145_ (.A1_N(_08080_),
    .A2_N(_08126_),
    .B1(\design_top.MEM[8][21] ),
    .B2(_08128_),
    .X(_06187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14146_ (.A1_N(_08081_),
    .A2_N(_08126_),
    .B1(\design_top.MEM[8][20] ),
    .B2(_08128_),
    .X(_06186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14147_ (.A1_N(_08082_),
    .A2_N(_08126_),
    .B1(\design_top.MEM[8][19] ),
    .B2(_08128_),
    .X(_06185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14148_ (.A1_N(_08083_),
    .A2_N(_08125_),
    .B1(\design_top.MEM[8][18] ),
    .B2(_08127_),
    .X(_06184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14149_ (.A1_N(_08084_),
    .A2_N(_08125_),
    .B1(\design_top.MEM[8][17] ),
    .B2(_08127_),
    .X(_06183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14150_ (.A1_N(_08085_),
    .A2_N(_08125_),
    .B1(\design_top.MEM[8][16] ),
    .B2(_08127_),
    .X(_06182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14151_ (.A(_07749_),
    .X(_08129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14152_ (.A(_08108_),
    .B(_08120_),
    .X(_08130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14153_ (.A(_08130_),
    .X(_08131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14154_ (.A1(_08057_),
    .A2(_11138_),
    .B1(_08130_),
    .X(_08132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14155_ (.A(_08132_),
    .X(_08133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14156_ (.A1_N(_08129_),
    .A2_N(_08131_),
    .B1(\design_top.MEM[8][15] ),
    .B2(_08133_),
    .X(_06181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14157_ (.A1_N(_08113_),
    .A2_N(_08131_),
    .B1(\design_top.MEM[8][14] ),
    .B2(_08133_),
    .X(_06180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14158_ (.A1_N(_08114_),
    .A2_N(_08131_),
    .B1(\design_top.MEM[8][13] ),
    .B2(_08133_),
    .X(_06179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14159_ (.A1_N(_08115_),
    .A2_N(_08131_),
    .B1(\design_top.MEM[8][12] ),
    .B2(_08133_),
    .X(_06178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14160_ (.A1_N(_08116_),
    .A2_N(_08131_),
    .B1(\design_top.MEM[8][11] ),
    .B2(_08133_),
    .X(_06177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14161_ (.A1_N(_08117_),
    .A2_N(_08130_),
    .B1(\design_top.MEM[8][10] ),
    .B2(_08132_),
    .X(_06176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14162_ (.A1_N(_08118_),
    .A2_N(_08130_),
    .B1(\design_top.MEM[8][9] ),
    .B2(_08132_),
    .X(_06175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14163_ (.A1_N(_08119_),
    .A2_N(_08130_),
    .B1(\design_top.MEM[8][8] ),
    .B2(_08132_),
    .X(_06174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14164_ (.A(_10782_),
    .B(_11040_),
    .X(_08134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14165_ (.A(_08087_),
    .B(_08134_),
    .X(_08135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14166_ (.A(_08135_),
    .X(_08136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14167_ (.A(_10889_),
    .X(_08137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14168_ (.A(_08137_),
    .X(_08138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14169_ (.A1(_08138_),
    .A2(_07869_),
    .B1(_08135_),
    .X(_08139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14170_ (.A(_08139_),
    .X(_08140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14171_ (.A1_N(_08086_),
    .A2_N(_08136_),
    .B1(\design_top.MEM[7][31] ),
    .B2(_08140_),
    .X(_06173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14172_ (.A1_N(_08092_),
    .A2_N(_08136_),
    .B1(\design_top.MEM[7][30] ),
    .B2(_08140_),
    .X(_06172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14173_ (.A1_N(_08093_),
    .A2_N(_08136_),
    .B1(\design_top.MEM[7][29] ),
    .B2(_08140_),
    .X(_06171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14174_ (.A1_N(_08094_),
    .A2_N(_08136_),
    .B1(\design_top.MEM[7][28] ),
    .B2(_08140_),
    .X(_06170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14175_ (.A1_N(_08095_),
    .A2_N(_08136_),
    .B1(\design_top.MEM[7][27] ),
    .B2(_08140_),
    .X(_06169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14176_ (.A1_N(_08096_),
    .A2_N(_08135_),
    .B1(\design_top.MEM[7][26] ),
    .B2(_08139_),
    .X(_06168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14177_ (.A1_N(_08097_),
    .A2_N(_08135_),
    .B1(\design_top.MEM[7][25] ),
    .B2(_08139_),
    .X(_06167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14178_ (.A1_N(_08098_),
    .A2_N(_08135_),
    .B1(\design_top.MEM[7][24] ),
    .B2(_08139_),
    .X(_06166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14179_ (.A(_08074_),
    .B(_08134_),
    .X(_08141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14180_ (.A(_08141_),
    .X(_08142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14181_ (.A1(_08138_),
    .A2(_07869_),
    .B1(_08141_),
    .X(_08143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14182_ (.A(_08143_),
    .X(_08144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14183_ (.A1_N(_08073_),
    .A2_N(_08142_),
    .B1(\design_top.MEM[7][23] ),
    .B2(_08144_),
    .X(_06165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14184_ (.A1_N(_08079_),
    .A2_N(_08142_),
    .B1(\design_top.MEM[7][22] ),
    .B2(_08144_),
    .X(_06164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14185_ (.A1_N(_08080_),
    .A2_N(_08142_),
    .B1(\design_top.MEM[7][21] ),
    .B2(_08144_),
    .X(_06163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14186_ (.A1_N(_08081_),
    .A2_N(_08142_),
    .B1(\design_top.MEM[7][20] ),
    .B2(_08144_),
    .X(_06162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14187_ (.A1_N(_08082_),
    .A2_N(_08142_),
    .B1(\design_top.MEM[7][19] ),
    .B2(_08144_),
    .X(_06161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14188_ (.A1_N(_08083_),
    .A2_N(_08141_),
    .B1(\design_top.MEM[7][18] ),
    .B2(_08143_),
    .X(_06160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14189_ (.A1_N(_08084_),
    .A2_N(_08141_),
    .B1(\design_top.MEM[7][17] ),
    .B2(_08143_),
    .X(_06159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14190_ (.A1_N(_08085_),
    .A2_N(_08141_),
    .B1(\design_top.MEM[7][16] ),
    .B2(_08143_),
    .X(_06158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14191_ (.A(_08108_),
    .B(_08134_),
    .X(_08145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14192_ (.A(_08145_),
    .X(_08146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14193_ (.A(_07868_),
    .X(_08147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14194_ (.A1(_08138_),
    .A2(_08147_),
    .B1(_08145_),
    .X(_08148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14195_ (.A(_08148_),
    .X(_08149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14196_ (.A1_N(_08129_),
    .A2_N(_08146_),
    .B1(\design_top.MEM[7][15] ),
    .B2(_08149_),
    .X(_06157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14197_ (.A1_N(_08113_),
    .A2_N(_08146_),
    .B1(\design_top.MEM[7][14] ),
    .B2(_08149_),
    .X(_06156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14198_ (.A1_N(_08114_),
    .A2_N(_08146_),
    .B1(\design_top.MEM[7][13] ),
    .B2(_08149_),
    .X(_06155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14199_ (.A1_N(_08115_),
    .A2_N(_08146_),
    .B1(\design_top.MEM[7][12] ),
    .B2(_08149_),
    .X(_06154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14200_ (.A1_N(_08116_),
    .A2_N(_08146_),
    .B1(\design_top.MEM[7][11] ),
    .B2(_08149_),
    .X(_06153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14201_ (.A1_N(_08117_),
    .A2_N(_08145_),
    .B1(\design_top.MEM[7][10] ),
    .B2(_08148_),
    .X(_06152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14202_ (.A1_N(_08118_),
    .A2_N(_08145_),
    .B1(\design_top.MEM[7][9] ),
    .B2(_08148_),
    .X(_06151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14203_ (.A1_N(_08119_),
    .A2_N(_08145_),
    .B1(\design_top.MEM[7][8] ),
    .B2(_08148_),
    .X(_06150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14204_ (.A(_10782_),
    .B(_11019_),
    .X(_08150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14205_ (.A(_08087_),
    .B(_08150_),
    .X(_08151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14206_ (.A(_08151_),
    .X(_08152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14207_ (.A(_07434_),
    .X(_08153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14208_ (.A1(_08153_),
    .A2(_08147_),
    .B1(_08151_),
    .X(_08154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14209_ (.A(_08154_),
    .X(_08155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14210_ (.A1_N(_08086_),
    .A2_N(_08152_),
    .B1(\design_top.MEM[6][31] ),
    .B2(_08155_),
    .X(_06149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14211_ (.A1_N(_08092_),
    .A2_N(_08152_),
    .B1(\design_top.MEM[6][30] ),
    .B2(_08155_),
    .X(_06148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14212_ (.A1_N(_08093_),
    .A2_N(_08152_),
    .B1(\design_top.MEM[6][29] ),
    .B2(_08155_),
    .X(_06147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14213_ (.A1_N(_08094_),
    .A2_N(_08152_),
    .B1(\design_top.MEM[6][28] ),
    .B2(_08155_),
    .X(_06146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14214_ (.A1_N(_08095_),
    .A2_N(_08152_),
    .B1(\design_top.MEM[6][27] ),
    .B2(_08155_),
    .X(_06145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14215_ (.A1_N(_08096_),
    .A2_N(_08151_),
    .B1(\design_top.MEM[6][26] ),
    .B2(_08154_),
    .X(_06144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14216_ (.A1_N(_08097_),
    .A2_N(_08151_),
    .B1(\design_top.MEM[6][25] ),
    .B2(_08154_),
    .X(_06143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14217_ (.A1_N(_08098_),
    .A2_N(_08151_),
    .B1(\design_top.MEM[6][24] ),
    .B2(_08154_),
    .X(_06142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14218_ (.A(_08074_),
    .B(_08150_),
    .X(_08156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14219_ (.A(_08156_),
    .X(_08157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14220_ (.A1(_08153_),
    .A2(_08147_),
    .B1(_08156_),
    .X(_08158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14221_ (.A(_08158_),
    .X(_08159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14222_ (.A1_N(_08073_),
    .A2_N(_08157_),
    .B1(\design_top.MEM[6][23] ),
    .B2(_08159_),
    .X(_06141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14223_ (.A1_N(_08079_),
    .A2_N(_08157_),
    .B1(\design_top.MEM[6][22] ),
    .B2(_08159_),
    .X(_06140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14224_ (.A1_N(_08080_),
    .A2_N(_08157_),
    .B1(\design_top.MEM[6][21] ),
    .B2(_08159_),
    .X(_06139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14225_ (.A1_N(_08081_),
    .A2_N(_08157_),
    .B1(\design_top.MEM[6][20] ),
    .B2(_08159_),
    .X(_06138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14226_ (.A1_N(_08082_),
    .A2_N(_08157_),
    .B1(\design_top.MEM[6][19] ),
    .B2(_08159_),
    .X(_06137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14227_ (.A1_N(_08083_),
    .A2_N(_08156_),
    .B1(\design_top.MEM[6][18] ),
    .B2(_08158_),
    .X(_06136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14228_ (.A1_N(_08084_),
    .A2_N(_08156_),
    .B1(\design_top.MEM[6][17] ),
    .B2(_08158_),
    .X(_06135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14229_ (.A1_N(_08085_),
    .A2_N(_08156_),
    .B1(\design_top.MEM[6][16] ),
    .B2(_08158_),
    .X(_06134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14230_ (.A(_08108_),
    .B(_08150_),
    .X(_08160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14231_ (.A(_08160_),
    .X(_08161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14232_ (.A1(_08153_),
    .A2(_08147_),
    .B1(_08160_),
    .X(_08162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14233_ (.A(_08162_),
    .X(_08163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14234_ (.A1_N(_08129_),
    .A2_N(_08161_),
    .B1(\design_top.MEM[6][15] ),
    .B2(_08163_),
    .X(_06133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14235_ (.A1_N(_08113_),
    .A2_N(_08161_),
    .B1(\design_top.MEM[6][14] ),
    .B2(_08163_),
    .X(_06132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14236_ (.A1_N(_08114_),
    .A2_N(_08161_),
    .B1(\design_top.MEM[6][13] ),
    .B2(_08163_),
    .X(_06131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14237_ (.A1_N(_08115_),
    .A2_N(_08161_),
    .B1(\design_top.MEM[6][12] ),
    .B2(_08163_),
    .X(_06130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14238_ (.A1_N(_08116_),
    .A2_N(_08161_),
    .B1(\design_top.MEM[6][11] ),
    .B2(_08163_),
    .X(_06129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14239_ (.A1_N(_08117_),
    .A2_N(_08160_),
    .B1(\design_top.MEM[6][10] ),
    .B2(_08162_),
    .X(_06128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14240_ (.A1_N(_08118_),
    .A2_N(_08160_),
    .B1(\design_top.MEM[6][9] ),
    .B2(_08162_),
    .X(_06127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14241_ (.A1_N(_08119_),
    .A2_N(_08160_),
    .B1(\design_top.MEM[6][8] ),
    .B2(_08162_),
    .X(_06126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14242_ (.A(_02860_),
    .B(_07556_),
    .X(_08164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14243_ (.A(_08164_),
    .X(_08165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14244_ (.A(_11039_),
    .B(_08165_),
    .X(_08166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14245_ (.A(_08108_),
    .B(_08166_),
    .X(_08167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14246_ (.A(_08167_),
    .X(_08168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _14247_ (.A(_11109_),
    .B(_10893_),
    .C(_10895_),
    .D(_10963_),
    .X(_08169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14248_ (.A(_08169_),
    .X(_08170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14249_ (.A(_08170_),
    .X(_08171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14250_ (.A1(_08138_),
    .A2(_08171_),
    .B1(_08167_),
    .X(_08172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14251_ (.A(_08172_),
    .X(_08173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14252_ (.A1_N(_08129_),
    .A2_N(_08168_),
    .B1(\design_top.MEM[63][15] ),
    .B2(_08173_),
    .X(_06125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14253_ (.A1_N(_08113_),
    .A2_N(_08168_),
    .B1(\design_top.MEM[63][14] ),
    .B2(_08173_),
    .X(_06124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14254_ (.A1_N(_08114_),
    .A2_N(_08168_),
    .B1(\design_top.MEM[63][13] ),
    .B2(_08173_),
    .X(_06123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14255_ (.A1_N(_08115_),
    .A2_N(_08168_),
    .B1(\design_top.MEM[63][12] ),
    .B2(_08173_),
    .X(_06122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14256_ (.A1_N(_08116_),
    .A2_N(_08168_),
    .B1(\design_top.MEM[63][11] ),
    .B2(_08173_),
    .X(_06121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14257_ (.A1_N(_08117_),
    .A2_N(_08167_),
    .B1(\design_top.MEM[63][10] ),
    .B2(_08172_),
    .X(_06120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14258_ (.A1_N(_08118_),
    .A2_N(_08167_),
    .B1(\design_top.MEM[63][9] ),
    .B2(_08172_),
    .X(_06119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14259_ (.A1_N(_08119_),
    .A2_N(_08167_),
    .B1(\design_top.MEM[63][8] ),
    .B2(_08172_),
    .X(_06118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14260_ (.A(_10874_),
    .X(_08174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14261_ (.A(_10877_),
    .X(_08175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14262_ (.A(_08175_),
    .B(_08166_),
    .X(_08176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14263_ (.A(_08176_),
    .X(_08177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14264_ (.A1(_08138_),
    .A2(_08171_),
    .B1(_08176_),
    .X(_08178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14265_ (.A(_08178_),
    .X(_08179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14266_ (.A1_N(_08174_),
    .A2_N(_08177_),
    .B1(\design_top.MEM[63][23] ),
    .B2(_08179_),
    .X(_06117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14267_ (.A(_10902_),
    .X(_08180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14268_ (.A1_N(_08180_),
    .A2_N(_08177_),
    .B1(\design_top.MEM[63][22] ),
    .B2(_08179_),
    .X(_06116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14269_ (.A(_10905_),
    .X(_08181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14270_ (.A1_N(_08181_),
    .A2_N(_08177_),
    .B1(\design_top.MEM[63][21] ),
    .B2(_08179_),
    .X(_06115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14271_ (.A(_10908_),
    .X(_08182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14272_ (.A1_N(_08182_),
    .A2_N(_08177_),
    .B1(\design_top.MEM[63][20] ),
    .B2(_08179_),
    .X(_06114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14273_ (.A(_10911_),
    .X(_08183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14274_ (.A1_N(_08183_),
    .A2_N(_08177_),
    .B1(\design_top.MEM[63][19] ),
    .B2(_08179_),
    .X(_06113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14275_ (.A(_10914_),
    .X(_08184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14276_ (.A1_N(_08184_),
    .A2_N(_08176_),
    .B1(\design_top.MEM[63][18] ),
    .B2(_08178_),
    .X(_06112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14277_ (.A(_10917_),
    .X(_08185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14278_ (.A1_N(_08185_),
    .A2_N(_08176_),
    .B1(\design_top.MEM[63][17] ),
    .B2(_08178_),
    .X(_06111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14279_ (.A(_10920_),
    .X(_08186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14280_ (.A1_N(_08186_),
    .A2_N(_08176_),
    .B1(\design_top.MEM[63][16] ),
    .B2(_08178_),
    .X(_06110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14281_ (.A(_08087_),
    .B(_08166_),
    .X(_08187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14282_ (.A(_08187_),
    .X(_08188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14283_ (.A(_08137_),
    .X(_08189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14284_ (.A1(_08189_),
    .A2(_08171_),
    .B1(_08187_),
    .X(_08190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14285_ (.A(_08190_),
    .X(_08191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14286_ (.A1_N(_08086_),
    .A2_N(_08188_),
    .B1(\design_top.MEM[63][31] ),
    .B2(_08191_),
    .X(_06109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14287_ (.A1_N(_08092_),
    .A2_N(_08188_),
    .B1(\design_top.MEM[63][30] ),
    .B2(_08191_),
    .X(_06108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14288_ (.A1_N(_08093_),
    .A2_N(_08188_),
    .B1(\design_top.MEM[63][29] ),
    .B2(_08191_),
    .X(_06107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14289_ (.A1_N(_08094_),
    .A2_N(_08188_),
    .B1(\design_top.MEM[63][28] ),
    .B2(_08191_),
    .X(_06106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14290_ (.A1_N(_08095_),
    .A2_N(_08188_),
    .B1(\design_top.MEM[63][27] ),
    .B2(_08191_),
    .X(_06105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14291_ (.A1_N(_08096_),
    .A2_N(_08187_),
    .B1(\design_top.MEM[63][26] ),
    .B2(_08190_),
    .X(_06104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14292_ (.A1_N(_08097_),
    .A2_N(_08187_),
    .B1(\design_top.MEM[63][25] ),
    .B2(_08190_),
    .X(_06103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14293_ (.A1_N(_08098_),
    .A2_N(_08187_),
    .B1(\design_top.MEM[63][24] ),
    .B2(_08190_),
    .X(_06102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14294_ (.A(_10767_),
    .X(_08192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14295_ (.A(_11018_),
    .B(_08165_),
    .X(_08193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14296_ (.A(_08192_),
    .B(_08193_),
    .X(_08194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14297_ (.A(_08194_),
    .X(_08195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14298_ (.A1(_08153_),
    .A2(_08171_),
    .B1(_08194_),
    .X(_08196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14299_ (.A(_08196_),
    .X(_08197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14300_ (.A1_N(_08129_),
    .A2_N(_08195_),
    .B1(\design_top.MEM[62][15] ),
    .B2(_08197_),
    .X(_06101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14301_ (.A(_10587_),
    .X(_08198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14302_ (.A1_N(_08198_),
    .A2_N(_08195_),
    .B1(\design_top.MEM[62][14] ),
    .B2(_08197_),
    .X(_06100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14303_ (.A(_10802_),
    .X(_08199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14304_ (.A1_N(_08199_),
    .A2_N(_08195_),
    .B1(\design_top.MEM[62][13] ),
    .B2(_08197_),
    .X(_06099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14305_ (.A(_10805_),
    .X(_08200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14306_ (.A1_N(_08200_),
    .A2_N(_08195_),
    .B1(\design_top.MEM[62][12] ),
    .B2(_08197_),
    .X(_06098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14307_ (.A(_10808_),
    .X(_08201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14308_ (.A1_N(_08201_),
    .A2_N(_08195_),
    .B1(\design_top.MEM[62][11] ),
    .B2(_08197_),
    .X(_06097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14309_ (.A(_10811_),
    .X(_08202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14310_ (.A1_N(_08202_),
    .A2_N(_08194_),
    .B1(\design_top.MEM[62][10] ),
    .B2(_08196_),
    .X(_06096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14311_ (.A(_10814_),
    .X(_08203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14312_ (.A1_N(_08203_),
    .A2_N(_08194_),
    .B1(\design_top.MEM[62][9] ),
    .B2(_08196_),
    .X(_06095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14313_ (.A(_10817_),
    .X(_08204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14314_ (.A1_N(_08204_),
    .A2_N(_08194_),
    .B1(\design_top.MEM[62][8] ),
    .B2(_08196_),
    .X(_06094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14315_ (.A(_08175_),
    .B(_08193_),
    .X(_08205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14316_ (.A(_08205_),
    .X(_08206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14317_ (.A1(_08153_),
    .A2(_08171_),
    .B1(_08205_),
    .X(_08207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14318_ (.A(_08207_),
    .X(_08208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14319_ (.A1_N(_08174_),
    .A2_N(_08206_),
    .B1(\design_top.MEM[62][23] ),
    .B2(_08208_),
    .X(_06093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14320_ (.A1_N(_08180_),
    .A2_N(_08206_),
    .B1(\design_top.MEM[62][22] ),
    .B2(_08208_),
    .X(_06092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14321_ (.A1_N(_08181_),
    .A2_N(_08206_),
    .B1(\design_top.MEM[62][21] ),
    .B2(_08208_),
    .X(_06091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14322_ (.A1_N(_08182_),
    .A2_N(_08206_),
    .B1(\design_top.MEM[62][20] ),
    .B2(_08208_),
    .X(_06090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14323_ (.A1_N(_08183_),
    .A2_N(_08206_),
    .B1(\design_top.MEM[62][19] ),
    .B2(_08208_),
    .X(_06089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14324_ (.A1_N(_08184_),
    .A2_N(_08205_),
    .B1(\design_top.MEM[62][18] ),
    .B2(_08207_),
    .X(_06088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14325_ (.A1_N(_08185_),
    .A2_N(_08205_),
    .B1(\design_top.MEM[62][17] ),
    .B2(_08207_),
    .X(_06087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14326_ (.A1_N(_08186_),
    .A2_N(_08205_),
    .B1(\design_top.MEM[62][16] ),
    .B2(_08207_),
    .X(_06086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14327_ (.A(_10820_),
    .X(_08209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14328_ (.A(_10925_),
    .X(_08210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14329_ (.A(_08210_),
    .B(_08193_),
    .X(_08211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14330_ (.A(_08211_),
    .X(_08212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14331_ (.A(_08170_),
    .X(_08213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14332_ (.A1(_11006_),
    .A2(_08213_),
    .B1(_08211_),
    .X(_08214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14333_ (.A(_08214_),
    .X(_08215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14334_ (.A1_N(_08209_),
    .A2_N(_08212_),
    .B1(\design_top.MEM[62][31] ),
    .B2(_08215_),
    .X(_06085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14335_ (.A(_10932_),
    .X(_08216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14336_ (.A1_N(_08216_),
    .A2_N(_08212_),
    .B1(\design_top.MEM[62][30] ),
    .B2(_08215_),
    .X(_06084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14337_ (.A(_10935_),
    .X(_08217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14338_ (.A1_N(_08217_),
    .A2_N(_08212_),
    .B1(\design_top.MEM[62][29] ),
    .B2(_08215_),
    .X(_06083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14339_ (.A(_10938_),
    .X(_08218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14340_ (.A1_N(_08218_),
    .A2_N(_08212_),
    .B1(\design_top.MEM[62][28] ),
    .B2(_08215_),
    .X(_06082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14341_ (.A(_10941_),
    .X(_08219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14342_ (.A1_N(_08219_),
    .A2_N(_08212_),
    .B1(\design_top.MEM[62][27] ),
    .B2(_08215_),
    .X(_06081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14343_ (.A(_10944_),
    .X(_08220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14344_ (.A1_N(_08220_),
    .A2_N(_08211_),
    .B1(\design_top.MEM[62][26] ),
    .B2(_08214_),
    .X(_06080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14345_ (.A(_10947_),
    .X(_08221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14346_ (.A1_N(_08221_),
    .A2_N(_08211_),
    .B1(\design_top.MEM[62][25] ),
    .B2(_08214_),
    .X(_06079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14347_ (.A(_10950_),
    .X(_08222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14348_ (.A1_N(_08222_),
    .A2_N(_08211_),
    .B1(\design_top.MEM[62][24] ),
    .B2(_08214_),
    .X(_06078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14349_ (.A(_10953_),
    .X(_08223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14350_ (.A(_10979_),
    .B(_08165_),
    .X(_08224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14351_ (.A(_08192_),
    .B(_08224_),
    .X(_08225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14352_ (.A(_08225_),
    .X(_08226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14353_ (.A1(_07998_),
    .A2(_08213_),
    .B1(_08225_),
    .X(_08227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14354_ (.A(_08227_),
    .X(_08228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14355_ (.A1_N(_08223_),
    .A2_N(_08226_),
    .B1(\design_top.MEM[61][15] ),
    .B2(_08228_),
    .X(_06077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14356_ (.A1_N(_08198_),
    .A2_N(_08226_),
    .B1(\design_top.MEM[61][14] ),
    .B2(_08228_),
    .X(_06076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14357_ (.A1_N(_08199_),
    .A2_N(_08226_),
    .B1(\design_top.MEM[61][13] ),
    .B2(_08228_),
    .X(_06075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14358_ (.A1_N(_08200_),
    .A2_N(_08226_),
    .B1(\design_top.MEM[61][12] ),
    .B2(_08228_),
    .X(_06074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14359_ (.A1_N(_08201_),
    .A2_N(_08226_),
    .B1(\design_top.MEM[61][11] ),
    .B2(_08228_),
    .X(_06073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14360_ (.A1_N(_08202_),
    .A2_N(_08225_),
    .B1(\design_top.MEM[61][10] ),
    .B2(_08227_),
    .X(_06072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14361_ (.A1_N(_08203_),
    .A2_N(_08225_),
    .B1(\design_top.MEM[61][9] ),
    .B2(_08227_),
    .X(_06071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14362_ (.A1_N(_08204_),
    .A2_N(_08225_),
    .B1(\design_top.MEM[61][8] ),
    .B2(_08227_),
    .X(_06070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14363_ (.A(_08175_),
    .B(_08224_),
    .X(_08229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14364_ (.A(_08229_),
    .X(_08230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14365_ (.A(_07508_),
    .X(_08231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14366_ (.A1(_08231_),
    .A2(_08213_),
    .B1(_08229_),
    .X(_08232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14367_ (.A(_08232_),
    .X(_08233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14368_ (.A1_N(_08174_),
    .A2_N(_08230_),
    .B1(\design_top.MEM[61][23] ),
    .B2(_08233_),
    .X(_06069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14369_ (.A1_N(_08180_),
    .A2_N(_08230_),
    .B1(\design_top.MEM[61][22] ),
    .B2(_08233_),
    .X(_06068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14370_ (.A1_N(_08181_),
    .A2_N(_08230_),
    .B1(\design_top.MEM[61][21] ),
    .B2(_08233_),
    .X(_06067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14371_ (.A1_N(_08182_),
    .A2_N(_08230_),
    .B1(\design_top.MEM[61][20] ),
    .B2(_08233_),
    .X(_06066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14372_ (.A1_N(_08183_),
    .A2_N(_08230_),
    .B1(\design_top.MEM[61][19] ),
    .B2(_08233_),
    .X(_06065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14373_ (.A1_N(_08184_),
    .A2_N(_08229_),
    .B1(\design_top.MEM[61][18] ),
    .B2(_08232_),
    .X(_06064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14374_ (.A1_N(_08185_),
    .A2_N(_08229_),
    .B1(\design_top.MEM[61][17] ),
    .B2(_08232_),
    .X(_06063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14375_ (.A1_N(_08186_),
    .A2_N(_08229_),
    .B1(\design_top.MEM[61][16] ),
    .B2(_08232_),
    .X(_06062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14376_ (.A(_08210_),
    .B(_08224_),
    .X(_08234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14377_ (.A(_08234_),
    .X(_08235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14378_ (.A1(_08231_),
    .A2(_08213_),
    .B1(_08234_),
    .X(_08236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14379_ (.A(_08236_),
    .X(_08237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14380_ (.A1_N(_08209_),
    .A2_N(_08235_),
    .B1(\design_top.MEM[61][31] ),
    .B2(_08237_),
    .X(_06061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14381_ (.A1_N(_08216_),
    .A2_N(_08235_),
    .B1(\design_top.MEM[61][30] ),
    .B2(_08237_),
    .X(_06060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14382_ (.A1_N(_08217_),
    .A2_N(_08235_),
    .B1(\design_top.MEM[61][29] ),
    .B2(_08237_),
    .X(_06059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14383_ (.A1_N(_08218_),
    .A2_N(_08235_),
    .B1(\design_top.MEM[61][28] ),
    .B2(_08237_),
    .X(_06058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14384_ (.A1_N(_08219_),
    .A2_N(_08235_),
    .B1(\design_top.MEM[61][27] ),
    .B2(_08237_),
    .X(_06057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14385_ (.A1_N(_08220_),
    .A2_N(_08234_),
    .B1(\design_top.MEM[61][26] ),
    .B2(_08236_),
    .X(_06056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14386_ (.A1_N(_08221_),
    .A2_N(_08234_),
    .B1(\design_top.MEM[61][25] ),
    .B2(_08236_),
    .X(_06055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14387_ (.A1_N(_08222_),
    .A2_N(_08234_),
    .B1(\design_top.MEM[61][24] ),
    .B2(_08236_),
    .X(_06054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14388_ (.A(_10957_),
    .B(_08165_),
    .X(_08238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14389_ (.A(_08192_),
    .B(_08238_),
    .X(_08239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14390_ (.A(_08239_),
    .X(_08240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14391_ (.A1(_08057_),
    .A2(_08213_),
    .B1(_08239_),
    .X(_08241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14392_ (.A(_08241_),
    .X(_08242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14393_ (.A1_N(_08223_),
    .A2_N(_08240_),
    .B1(\design_top.MEM[60][15] ),
    .B2(_08242_),
    .X(_06053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14394_ (.A1_N(_08198_),
    .A2_N(_08240_),
    .B1(\design_top.MEM[60][14] ),
    .B2(_08242_),
    .X(_06052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14395_ (.A1_N(_08199_),
    .A2_N(_08240_),
    .B1(\design_top.MEM[60][13] ),
    .B2(_08242_),
    .X(_06051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14396_ (.A1_N(_08200_),
    .A2_N(_08240_),
    .B1(\design_top.MEM[60][12] ),
    .B2(_08242_),
    .X(_06050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14397_ (.A1_N(_08201_),
    .A2_N(_08240_),
    .B1(\design_top.MEM[60][11] ),
    .B2(_08242_),
    .X(_06049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14398_ (.A1_N(_08202_),
    .A2_N(_08239_),
    .B1(\design_top.MEM[60][10] ),
    .B2(_08241_),
    .X(_06048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14399_ (.A1_N(_08203_),
    .A2_N(_08239_),
    .B1(\design_top.MEM[60][9] ),
    .B2(_08241_),
    .X(_06047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14400_ (.A1_N(_08204_),
    .A2_N(_08239_),
    .B1(\design_top.MEM[60][8] ),
    .B2(_08241_),
    .X(_06046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14401_ (.A(_08175_),
    .B(_08238_),
    .X(_08243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14402_ (.A(_08243_),
    .X(_08244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14403_ (.A(_08056_),
    .X(_08245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14404_ (.A1(_08245_),
    .A2(_08170_),
    .B1(_08243_),
    .X(_08246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14405_ (.A(_08246_),
    .X(_08247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14406_ (.A1_N(_08174_),
    .A2_N(_08244_),
    .B1(\design_top.MEM[60][23] ),
    .B2(_08247_),
    .X(_06045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14407_ (.A1_N(_08180_),
    .A2_N(_08244_),
    .B1(\design_top.MEM[60][22] ),
    .B2(_08247_),
    .X(_06044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14408_ (.A1_N(_08181_),
    .A2_N(_08244_),
    .B1(\design_top.MEM[60][21] ),
    .B2(_08247_),
    .X(_06043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14409_ (.A1_N(_08182_),
    .A2_N(_08244_),
    .B1(\design_top.MEM[60][20] ),
    .B2(_08247_),
    .X(_06042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14410_ (.A1_N(_08183_),
    .A2_N(_08244_),
    .B1(\design_top.MEM[60][19] ),
    .B2(_08247_),
    .X(_06041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14411_ (.A1_N(_08184_),
    .A2_N(_08243_),
    .B1(\design_top.MEM[60][18] ),
    .B2(_08246_),
    .X(_06040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14412_ (.A1_N(_08185_),
    .A2_N(_08243_),
    .B1(\design_top.MEM[60][17] ),
    .B2(_08246_),
    .X(_06039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14413_ (.A1_N(_08186_),
    .A2_N(_08243_),
    .B1(\design_top.MEM[60][16] ),
    .B2(_08246_),
    .X(_06038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14414_ (.A(_08210_),
    .B(_08238_),
    .X(_08248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14415_ (.A(_08248_),
    .X(_08249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14416_ (.A1(_08245_),
    .A2(_08170_),
    .B1(_08248_),
    .X(_08250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14417_ (.A(_08250_),
    .X(_08251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14418_ (.A1_N(_08209_),
    .A2_N(_08249_),
    .B1(\design_top.MEM[60][31] ),
    .B2(_08251_),
    .X(_06037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14419_ (.A1_N(_08216_),
    .A2_N(_08249_),
    .B1(\design_top.MEM[60][30] ),
    .B2(_08251_),
    .X(_06036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14420_ (.A1_N(_08217_),
    .A2_N(_08249_),
    .B1(\design_top.MEM[60][29] ),
    .B2(_08251_),
    .X(_06035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14421_ (.A1_N(_08218_),
    .A2_N(_08249_),
    .B1(\design_top.MEM[60][28] ),
    .B2(_08251_),
    .X(_06034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14422_ (.A1_N(_08219_),
    .A2_N(_08249_),
    .B1(\design_top.MEM[60][27] ),
    .B2(_08251_),
    .X(_06033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14423_ (.A1_N(_08220_),
    .A2_N(_08248_),
    .B1(\design_top.MEM[60][26] ),
    .B2(_08250_),
    .X(_06032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14424_ (.A1_N(_08221_),
    .A2_N(_08248_),
    .B1(\design_top.MEM[60][25] ),
    .B2(_08250_),
    .X(_06031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14425_ (.A1_N(_08222_),
    .A2_N(_08248_),
    .B1(\design_top.MEM[60][24] ),
    .B2(_08250_),
    .X(_06030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14426_ (.A(_10782_),
    .B(_10980_),
    .X(_08252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14427_ (.A(_08210_),
    .B(_08252_),
    .X(_08253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14428_ (.A(_08253_),
    .X(_08254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14429_ (.A1(_08231_),
    .A2(_08147_),
    .B1(_08253_),
    .X(_08255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14430_ (.A(_08255_),
    .X(_08256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14431_ (.A1_N(_08209_),
    .A2_N(_08254_),
    .B1(\design_top.MEM[5][31] ),
    .B2(_08256_),
    .X(_06029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14432_ (.A1_N(_08216_),
    .A2_N(_08254_),
    .B1(\design_top.MEM[5][30] ),
    .B2(_08256_),
    .X(_06028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14433_ (.A1_N(_08217_),
    .A2_N(_08254_),
    .B1(\design_top.MEM[5][29] ),
    .B2(_08256_),
    .X(_06027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14434_ (.A1_N(_08218_),
    .A2_N(_08254_),
    .B1(\design_top.MEM[5][28] ),
    .B2(_08256_),
    .X(_06026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14435_ (.A1_N(_08219_),
    .A2_N(_08254_),
    .B1(\design_top.MEM[5][27] ),
    .B2(_08256_),
    .X(_06025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14436_ (.A1_N(_08220_),
    .A2_N(_08253_),
    .B1(\design_top.MEM[5][26] ),
    .B2(_08255_),
    .X(_06024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14437_ (.A1_N(_08221_),
    .A2_N(_08253_),
    .B1(\design_top.MEM[5][25] ),
    .B2(_08255_),
    .X(_06023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14438_ (.A1_N(_08222_),
    .A2_N(_08253_),
    .B1(\design_top.MEM[5][24] ),
    .B2(_08255_),
    .X(_06022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14439_ (.A(_08175_),
    .B(_08252_),
    .X(_08257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14440_ (.A(_08257_),
    .X(_08258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14441_ (.A1(_08231_),
    .A2(_07868_),
    .B1(_08257_),
    .X(_08259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14442_ (.A(_08259_),
    .X(_08260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14443_ (.A1_N(_08174_),
    .A2_N(_08258_),
    .B1(\design_top.MEM[5][23] ),
    .B2(_08260_),
    .X(_06021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14444_ (.A1_N(_08180_),
    .A2_N(_08258_),
    .B1(\design_top.MEM[5][22] ),
    .B2(_08260_),
    .X(_06020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14445_ (.A1_N(_08181_),
    .A2_N(_08258_),
    .B1(\design_top.MEM[5][21] ),
    .B2(_08260_),
    .X(_06019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14446_ (.A1_N(_08182_),
    .A2_N(_08258_),
    .B1(\design_top.MEM[5][20] ),
    .B2(_08260_),
    .X(_06018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14447_ (.A1_N(_08183_),
    .A2_N(_08258_),
    .B1(\design_top.MEM[5][19] ),
    .B2(_08260_),
    .X(_06017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14448_ (.A1_N(_08184_),
    .A2_N(_08257_),
    .B1(\design_top.MEM[5][18] ),
    .B2(_08259_),
    .X(_06016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14449_ (.A1_N(_08185_),
    .A2_N(_08257_),
    .B1(\design_top.MEM[5][17] ),
    .B2(_08259_),
    .X(_06015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14450_ (.A1_N(_08186_),
    .A2_N(_08257_),
    .B1(\design_top.MEM[5][16] ),
    .B2(_08259_),
    .X(_06014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14451_ (.A(_08192_),
    .B(_08252_),
    .X(_08261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14452_ (.A(_08261_),
    .X(_08262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14453_ (.A1(_08231_),
    .A2(_07868_),
    .B1(_08261_),
    .X(_08263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14454_ (.A(_08263_),
    .X(_08264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14455_ (.A1_N(_08223_),
    .A2_N(_08262_),
    .B1(\design_top.MEM[5][15] ),
    .B2(_08264_),
    .X(_06013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14456_ (.A1_N(_08198_),
    .A2_N(_08262_),
    .B1(\design_top.MEM[5][14] ),
    .B2(_08264_),
    .X(_06012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14457_ (.A1_N(_08199_),
    .A2_N(_08262_),
    .B1(\design_top.MEM[5][13] ),
    .B2(_08264_),
    .X(_06011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14458_ (.A1_N(_08200_),
    .A2_N(_08262_),
    .B1(\design_top.MEM[5][12] ),
    .B2(_08264_),
    .X(_06010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14459_ (.A1_N(_08201_),
    .A2_N(_08262_),
    .B1(\design_top.MEM[5][11] ),
    .B2(_08264_),
    .X(_06009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14460_ (.A1_N(_08202_),
    .A2_N(_08261_),
    .B1(\design_top.MEM[5][10] ),
    .B2(_08263_),
    .X(_06008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14461_ (.A1_N(_08203_),
    .A2_N(_08261_),
    .B1(\design_top.MEM[5][9] ),
    .B2(_08263_),
    .X(_06007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14462_ (.A1_N(_08204_),
    .A2_N(_08261_),
    .B1(\design_top.MEM[5][8] ),
    .B2(_08263_),
    .X(_06006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14463_ (.A(_10884_),
    .B(_08165_),
    .X(_08265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14464_ (.A(_08192_),
    .B(_08265_),
    .X(_08266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14465_ (.A(_08266_),
    .X(_08267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _14466_ (.A(_11109_),
    .B(_10893_),
    .C(_10895_),
    .D(wbs_adr_i[0]),
    .X(_08268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14467_ (.A(_08268_),
    .X(_08269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14468_ (.A(_08269_),
    .X(_08270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14469_ (.A1(_08189_),
    .A2(_08270_),
    .B1(_08266_),
    .X(_08271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14470_ (.A(_08271_),
    .X(_08272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14471_ (.A1_N(_08223_),
    .A2_N(_08267_),
    .B1(\design_top.MEM[59][15] ),
    .B2(_08272_),
    .X(_06005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14472_ (.A1_N(_08198_),
    .A2_N(_08267_),
    .B1(\design_top.MEM[59][14] ),
    .B2(_08272_),
    .X(_06004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14473_ (.A1_N(_08199_),
    .A2_N(_08267_),
    .B1(\design_top.MEM[59][13] ),
    .B2(_08272_),
    .X(_06003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14474_ (.A1_N(_08200_),
    .A2_N(_08267_),
    .B1(\design_top.MEM[59][12] ),
    .B2(_08272_),
    .X(_06002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14475_ (.A1_N(_08201_),
    .A2_N(_08267_),
    .B1(\design_top.MEM[59][11] ),
    .B2(_08272_),
    .X(_06001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14476_ (.A1_N(_08202_),
    .A2_N(_08266_),
    .B1(\design_top.MEM[59][10] ),
    .B2(_08271_),
    .X(_06000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14477_ (.A1_N(_08203_),
    .A2_N(_08266_),
    .B1(\design_top.MEM[59][9] ),
    .B2(_08271_),
    .X(_05999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14478_ (.A1_N(_08204_),
    .A2_N(_08266_),
    .B1(\design_top.MEM[59][8] ),
    .B2(_08271_),
    .X(_05998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14479_ (.A(_10878_),
    .B(_08265_),
    .X(_08273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14480_ (.A(_08273_),
    .X(_08274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14481_ (.A1(_08189_),
    .A2(_08270_),
    .B1(_08273_),
    .X(_08275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14482_ (.A(_08275_),
    .X(_08276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14483_ (.A1_N(_10875_),
    .A2_N(_08274_),
    .B1(\design_top.MEM[59][23] ),
    .B2(_08276_),
    .X(_05997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14484_ (.A1_N(_10903_),
    .A2_N(_08274_),
    .B1(\design_top.MEM[59][22] ),
    .B2(_08276_),
    .X(_05996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14485_ (.A1_N(_10906_),
    .A2_N(_08274_),
    .B1(\design_top.MEM[59][21] ),
    .B2(_08276_),
    .X(_05995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14486_ (.A1_N(_10909_),
    .A2_N(_08274_),
    .B1(\design_top.MEM[59][20] ),
    .B2(_08276_),
    .X(_05994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14487_ (.A1_N(_10912_),
    .A2_N(_08274_),
    .B1(\design_top.MEM[59][19] ),
    .B2(_08276_),
    .X(_05993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14488_ (.A1_N(_10915_),
    .A2_N(_08273_),
    .B1(\design_top.MEM[59][18] ),
    .B2(_08275_),
    .X(_05992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14489_ (.A1_N(_10918_),
    .A2_N(_08273_),
    .B1(\design_top.MEM[59][17] ),
    .B2(_08275_),
    .X(_05991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14490_ (.A1_N(_10921_),
    .A2_N(_08273_),
    .B1(\design_top.MEM[59][16] ),
    .B2(_08275_),
    .X(_05990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14491_ (.A(_08210_),
    .B(_08265_),
    .X(_08277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14492_ (.A(_08277_),
    .X(_08278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14493_ (.A1(_08189_),
    .A2(_08270_),
    .B1(_08277_),
    .X(_08279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14494_ (.A(_08279_),
    .X(_08280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14495_ (.A1_N(_08209_),
    .A2_N(_08278_),
    .B1(\design_top.MEM[59][31] ),
    .B2(_08280_),
    .X(_05989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14496_ (.A1_N(_08216_),
    .A2_N(_08278_),
    .B1(\design_top.MEM[59][30] ),
    .B2(_08280_),
    .X(_05988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14497_ (.A1_N(_08217_),
    .A2_N(_08278_),
    .B1(\design_top.MEM[59][29] ),
    .B2(_08280_),
    .X(_05987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14498_ (.A1_N(_08218_),
    .A2_N(_08278_),
    .B1(\design_top.MEM[59][28] ),
    .B2(_08280_),
    .X(_05986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14499_ (.A1_N(_08219_),
    .A2_N(_08278_),
    .B1(\design_top.MEM[59][27] ),
    .B2(_08280_),
    .X(_05985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14500_ (.A1_N(_08220_),
    .A2_N(_08277_),
    .B1(\design_top.MEM[59][26] ),
    .B2(_08279_),
    .X(_05984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14501_ (.A1_N(_08221_),
    .A2_N(_08277_),
    .B1(\design_top.MEM[59][25] ),
    .B2(_08279_),
    .X(_05983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14502_ (.A1_N(_08222_),
    .A2_N(_08277_),
    .B1(\design_top.MEM[59][24] ),
    .B2(_08279_),
    .X(_05982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14503_ (.A(_10999_),
    .B(_08164_),
    .X(_08281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14504_ (.A(_10768_),
    .B(_08281_),
    .X(_08282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14505_ (.A(_08282_),
    .X(_08283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14506_ (.A1(_11006_),
    .A2(_08270_),
    .B1(_08282_),
    .X(_08284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14507_ (.A(_08284_),
    .X(_08285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14508_ (.A1_N(_08223_),
    .A2_N(_08283_),
    .B1(\design_top.MEM[58][15] ),
    .B2(_08285_),
    .X(_05981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14509_ (.A1_N(_10588_),
    .A2_N(_08283_),
    .B1(\design_top.MEM[58][14] ),
    .B2(_08285_),
    .X(_05980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14510_ (.A1_N(_10803_),
    .A2_N(_08283_),
    .B1(\design_top.MEM[58][13] ),
    .B2(_08285_),
    .X(_05979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14511_ (.A1_N(_10806_),
    .A2_N(_08283_),
    .B1(\design_top.MEM[58][12] ),
    .B2(_08285_),
    .X(_05978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14512_ (.A1_N(_10809_),
    .A2_N(_08283_),
    .B1(\design_top.MEM[58][11] ),
    .B2(_08285_),
    .X(_05977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14513_ (.A1_N(_10812_),
    .A2_N(_08282_),
    .B1(\design_top.MEM[58][10] ),
    .B2(_08284_),
    .X(_05976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14514_ (.A1_N(_10815_),
    .A2_N(_08282_),
    .B1(\design_top.MEM[58][9] ),
    .B2(_08284_),
    .X(_05975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14515_ (.A1_N(_10818_),
    .A2_N(_08282_),
    .B1(\design_top.MEM[58][8] ),
    .B2(_08284_),
    .X(_05974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14516_ (.A(_10878_),
    .B(_08281_),
    .X(_08286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14517_ (.A(_08286_),
    .X(_08287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14518_ (.A1(_11006_),
    .A2(_08270_),
    .B1(_08286_),
    .X(_08288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14519_ (.A(_08288_),
    .X(_08289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14520_ (.A1_N(_10875_),
    .A2_N(_08287_),
    .B1(\design_top.MEM[58][23] ),
    .B2(_08289_),
    .X(_05973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14521_ (.A1_N(_10903_),
    .A2_N(_08287_),
    .B1(\design_top.MEM[58][22] ),
    .B2(_08289_),
    .X(_05972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14522_ (.A1_N(_10906_),
    .A2_N(_08287_),
    .B1(\design_top.MEM[58][21] ),
    .B2(_08289_),
    .X(_05971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14523_ (.A1_N(_10909_),
    .A2_N(_08287_),
    .B1(\design_top.MEM[58][20] ),
    .B2(_08289_),
    .X(_05970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14524_ (.A1_N(_10912_),
    .A2_N(_08287_),
    .B1(\design_top.MEM[58][19] ),
    .B2(_08289_),
    .X(_05969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14525_ (.A1_N(_10915_),
    .A2_N(_08286_),
    .B1(\design_top.MEM[58][18] ),
    .B2(_08288_),
    .X(_05968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14526_ (.A1_N(_10918_),
    .A2_N(_08286_),
    .B1(\design_top.MEM[58][17] ),
    .B2(_08288_),
    .X(_05967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14527_ (.A1_N(_10921_),
    .A2_N(_08286_),
    .B1(\design_top.MEM[58][16] ),
    .B2(_08288_),
    .X(_05966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14528_ (.A(_10926_),
    .B(_08281_),
    .X(_08290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14529_ (.A(_08290_),
    .X(_08291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14530_ (.A(_08269_),
    .X(_08292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14531_ (.A1(_11006_),
    .A2(_08292_),
    .B1(_08290_),
    .X(_08293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14532_ (.A(_08293_),
    .X(_08294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14533_ (.A1_N(_10923_),
    .A2_N(_08291_),
    .B1(\design_top.MEM[58][31] ),
    .B2(_08294_),
    .X(_05965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14534_ (.A1_N(_10933_),
    .A2_N(_08291_),
    .B1(\design_top.MEM[58][30] ),
    .B2(_08294_),
    .X(_05964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14535_ (.A1_N(_10936_),
    .A2_N(_08291_),
    .B1(\design_top.MEM[58][29] ),
    .B2(_08294_),
    .X(_05963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14536_ (.A1_N(_10939_),
    .A2_N(_08291_),
    .B1(\design_top.MEM[58][28] ),
    .B2(_08294_),
    .X(_05962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14537_ (.A1_N(_10942_),
    .A2_N(_08291_),
    .B1(\design_top.MEM[58][27] ),
    .B2(_08294_),
    .X(_05961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14538_ (.A1_N(_10945_),
    .A2_N(_08290_),
    .B1(\design_top.MEM[58][26] ),
    .B2(_08293_),
    .X(_05960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14539_ (.A1_N(_10948_),
    .A2_N(_08290_),
    .B1(\design_top.MEM[58][25] ),
    .B2(_08293_),
    .X(_05959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14540_ (.A1_N(_10951_),
    .A2_N(_08290_),
    .B1(\design_top.MEM[58][24] ),
    .B2(_08293_),
    .X(_05958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14541_ (.A(_11275_),
    .B(_08164_),
    .X(_08295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14542_ (.A(_10768_),
    .B(_08295_),
    .X(_08296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14543_ (.A(_08296_),
    .X(_08297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14544_ (.A1(_10987_),
    .A2(_08292_),
    .B1(_08296_),
    .X(_08298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14545_ (.A(_08298_),
    .X(_08299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14546_ (.A1_N(_10954_),
    .A2_N(_08297_),
    .B1(\design_top.MEM[57][15] ),
    .B2(_08299_),
    .X(_05957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14547_ (.A1_N(_10588_),
    .A2_N(_08297_),
    .B1(\design_top.MEM[57][14] ),
    .B2(_08299_),
    .X(_05956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14548_ (.A1_N(_10803_),
    .A2_N(_08297_),
    .B1(\design_top.MEM[57][13] ),
    .B2(_08299_),
    .X(_05955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14549_ (.A1_N(_10806_),
    .A2_N(_08297_),
    .B1(\design_top.MEM[57][12] ),
    .B2(_08299_),
    .X(_05954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14550_ (.A1_N(_10809_),
    .A2_N(_08297_),
    .B1(\design_top.MEM[57][11] ),
    .B2(_08299_),
    .X(_05953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14551_ (.A1_N(_10812_),
    .A2_N(_08296_),
    .B1(\design_top.MEM[57][10] ),
    .B2(_08298_),
    .X(_05952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14552_ (.A1_N(_10815_),
    .A2_N(_08296_),
    .B1(\design_top.MEM[57][9] ),
    .B2(_08298_),
    .X(_05951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14553_ (.A1_N(_10818_),
    .A2_N(_08296_),
    .B1(\design_top.MEM[57][8] ),
    .B2(_08298_),
    .X(_05950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14554_ (.A(_10878_),
    .B(_08295_),
    .X(_08300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14555_ (.A(_08300_),
    .X(_08301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14556_ (.A1(_10987_),
    .A2(_08292_),
    .B1(_08300_),
    .X(_08302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14557_ (.A(_08302_),
    .X(_08303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14558_ (.A1_N(_10875_),
    .A2_N(_08301_),
    .B1(\design_top.MEM[57][23] ),
    .B2(_08303_),
    .X(_05949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14559_ (.A1_N(_10903_),
    .A2_N(_08301_),
    .B1(\design_top.MEM[57][22] ),
    .B2(_08303_),
    .X(_05948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14560_ (.A1_N(_10906_),
    .A2_N(_08301_),
    .B1(\design_top.MEM[57][21] ),
    .B2(_08303_),
    .X(_05947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14561_ (.A1_N(_10909_),
    .A2_N(_08301_),
    .B1(\design_top.MEM[57][20] ),
    .B2(_08303_),
    .X(_05946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14562_ (.A1_N(_10912_),
    .A2_N(_08301_),
    .B1(\design_top.MEM[57][19] ),
    .B2(_08303_),
    .X(_05945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14563_ (.A1_N(_10915_),
    .A2_N(_08300_),
    .B1(\design_top.MEM[57][18] ),
    .B2(_08302_),
    .X(_05944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14564_ (.A1_N(_10918_),
    .A2_N(_08300_),
    .B1(\design_top.MEM[57][17] ),
    .B2(_08302_),
    .X(_05943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14565_ (.A1_N(_10921_),
    .A2_N(_08300_),
    .B1(\design_top.MEM[57][16] ),
    .B2(_08302_),
    .X(_05942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14566_ (.A(_10926_),
    .B(_08295_),
    .X(_08304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14567_ (.A(_08304_),
    .X(_08305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14568_ (.A1(_10987_),
    .A2(_08292_),
    .B1(_08304_),
    .X(_08306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14569_ (.A(_08306_),
    .X(_08307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14570_ (.A1_N(_10923_),
    .A2_N(_08305_),
    .B1(\design_top.MEM[57][31] ),
    .B2(_08307_),
    .X(_05941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14571_ (.A1_N(_10933_),
    .A2_N(_08305_),
    .B1(\design_top.MEM[57][30] ),
    .B2(_08307_),
    .X(_05940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14572_ (.A1_N(_10936_),
    .A2_N(_08305_),
    .B1(\design_top.MEM[57][29] ),
    .B2(_08307_),
    .X(_05939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14573_ (.A1_N(_10939_),
    .A2_N(_08305_),
    .B1(\design_top.MEM[57][28] ),
    .B2(_08307_),
    .X(_05938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14574_ (.A1_N(_10942_),
    .A2_N(_08305_),
    .B1(\design_top.MEM[57][27] ),
    .B2(_08307_),
    .X(_05937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14575_ (.A1_N(_10945_),
    .A2_N(_08304_),
    .B1(\design_top.MEM[57][26] ),
    .B2(_08306_),
    .X(_05936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14576_ (.A1_N(_10948_),
    .A2_N(_08304_),
    .B1(\design_top.MEM[57][25] ),
    .B2(_08306_),
    .X(_05935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14577_ (.A1_N(_10951_),
    .A2_N(_08304_),
    .B1(\design_top.MEM[57][24] ),
    .B2(_08306_),
    .X(_05934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14578_ (.A(_10776_),
    .B(_08164_),
    .X(_08308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14579_ (.A(_10768_),
    .B(_08308_),
    .X(_08309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14580_ (.A(_08309_),
    .X(_08310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14581_ (.A1(_08245_),
    .A2(_08292_),
    .B1(_08309_),
    .X(_08311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14582_ (.A(_08311_),
    .X(_08312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14583_ (.A1_N(_10954_),
    .A2_N(_08310_),
    .B1(\design_top.MEM[56][15] ),
    .B2(_08312_),
    .X(_05933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14584_ (.A1_N(_10588_),
    .A2_N(_08310_),
    .B1(\design_top.MEM[56][14] ),
    .B2(_08312_),
    .X(_05932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14585_ (.A1_N(_10803_),
    .A2_N(_08310_),
    .B1(\design_top.MEM[56][13] ),
    .B2(_08312_),
    .X(_05931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14586_ (.A1_N(_10806_),
    .A2_N(_08310_),
    .B1(\design_top.MEM[56][12] ),
    .B2(_08312_),
    .X(_05930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14587_ (.A1_N(_10809_),
    .A2_N(_08310_),
    .B1(\design_top.MEM[56][11] ),
    .B2(_08312_),
    .X(_05929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14588_ (.A1_N(_10812_),
    .A2_N(_08309_),
    .B1(\design_top.MEM[56][10] ),
    .B2(_08311_),
    .X(_05928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14589_ (.A1_N(_10815_),
    .A2_N(_08309_),
    .B1(\design_top.MEM[56][9] ),
    .B2(_08311_),
    .X(_05927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14590_ (.A1_N(_10818_),
    .A2_N(_08309_),
    .B1(\design_top.MEM[56][8] ),
    .B2(_08311_),
    .X(_05926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14591_ (.A(_10878_),
    .B(_08308_),
    .X(_08313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14592_ (.A(_08313_),
    .X(_08314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14593_ (.A1(_08245_),
    .A2(_08269_),
    .B1(_08313_),
    .X(_08315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14594_ (.A(_08315_),
    .X(_08316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14595_ (.A1_N(_10875_),
    .A2_N(_08314_),
    .B1(\design_top.MEM[56][23] ),
    .B2(_08316_),
    .X(_05925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14596_ (.A1_N(_10903_),
    .A2_N(_08314_),
    .B1(\design_top.MEM[56][22] ),
    .B2(_08316_),
    .X(_05924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14597_ (.A1_N(_10906_),
    .A2_N(_08314_),
    .B1(\design_top.MEM[56][21] ),
    .B2(_08316_),
    .X(_05923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14598_ (.A1_N(_10909_),
    .A2_N(_08314_),
    .B1(\design_top.MEM[56][20] ),
    .B2(_08316_),
    .X(_05922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14599_ (.A1_N(_10912_),
    .A2_N(_08314_),
    .B1(\design_top.MEM[56][19] ),
    .B2(_08316_),
    .X(_05921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14600_ (.A1_N(_10915_),
    .A2_N(_08313_),
    .B1(\design_top.MEM[56][18] ),
    .B2(_08315_),
    .X(_05920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14601_ (.A1_N(_10918_),
    .A2_N(_08313_),
    .B1(\design_top.MEM[56][17] ),
    .B2(_08315_),
    .X(_05919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14602_ (.A1_N(_10921_),
    .A2_N(_08313_),
    .B1(\design_top.MEM[56][16] ),
    .B2(_08315_),
    .X(_05918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14603_ (.A(_10926_),
    .B(_08308_),
    .X(_08317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14604_ (.A(_08317_),
    .X(_08318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14605_ (.A1(_08245_),
    .A2(_08269_),
    .B1(_08317_),
    .X(_08319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14606_ (.A(_08319_),
    .X(_08320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14607_ (.A1_N(_10923_),
    .A2_N(_08318_),
    .B1(\design_top.MEM[56][31] ),
    .B2(_08320_),
    .X(_05917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14608_ (.A1_N(_10933_),
    .A2_N(_08318_),
    .B1(\design_top.MEM[56][30] ),
    .B2(_08320_),
    .X(_05916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14609_ (.A1_N(_10936_),
    .A2_N(_08318_),
    .B1(\design_top.MEM[56][29] ),
    .B2(_08320_),
    .X(_05915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14610_ (.A1_N(_10939_),
    .A2_N(_08318_),
    .B1(\design_top.MEM[56][28] ),
    .B2(_08320_),
    .X(_05914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14611_ (.A1_N(_10942_),
    .A2_N(_08318_),
    .B1(\design_top.MEM[56][27] ),
    .B2(_08320_),
    .X(_05913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14612_ (.A1_N(_10945_),
    .A2_N(_08317_),
    .B1(\design_top.MEM[56][26] ),
    .B2(_08319_),
    .X(_05912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14613_ (.A1_N(_10948_),
    .A2_N(_08317_),
    .B1(\design_top.MEM[56][25] ),
    .B2(_08319_),
    .X(_05911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14614_ (.A1_N(_10951_),
    .A2_N(_08317_),
    .B1(\design_top.MEM[56][24] ),
    .B2(_08319_),
    .X(_05910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14615_ (.A(_10768_),
    .B(_07624_),
    .X(_08321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14616_ (.A(_08321_),
    .X(_08322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14617_ (.A1(_08189_),
    .A2(_07572_),
    .B1(_08321_),
    .X(_08323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14618_ (.A(_08323_),
    .X(_08324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14619_ (.A1_N(_10954_),
    .A2_N(_08322_),
    .B1(\design_top.MEM[55][15] ),
    .B2(_08324_),
    .X(_05909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14620_ (.A1_N(_10588_),
    .A2_N(_08322_),
    .B1(\design_top.MEM[55][14] ),
    .B2(_08324_),
    .X(_05908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14621_ (.A1_N(_10803_),
    .A2_N(_08322_),
    .B1(\design_top.MEM[55][13] ),
    .B2(_08324_),
    .X(_05907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14622_ (.A1_N(_10806_),
    .A2_N(_08322_),
    .B1(\design_top.MEM[55][12] ),
    .B2(_08324_),
    .X(_05906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14623_ (.A1_N(_10809_),
    .A2_N(_08322_),
    .B1(\design_top.MEM[55][11] ),
    .B2(_08324_),
    .X(_05905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14624_ (.A1_N(_10812_),
    .A2_N(_08321_),
    .B1(\design_top.MEM[55][10] ),
    .B2(_08323_),
    .X(_05904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14625_ (.A1_N(_10815_),
    .A2_N(_08321_),
    .B1(\design_top.MEM[55][9] ),
    .B2(_08323_),
    .X(_05903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14626_ (.A1_N(_10818_),
    .A2_N(_08321_),
    .B1(\design_top.MEM[55][8] ),
    .B2(_08323_),
    .X(_05902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _14627_ (.A1(_02643_),
    .A2(_10822_),
    .A3(_10821_),
    .B1(_10712_),
    .B2(_10714_),
    .X(_08325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14628_ (.A(_10823_),
    .B(_08325_),
    .X(_03200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _14629_ (.A(_02651_),
    .B(_03200_),
    .C(_02660_),
    .D(_10828_),
    .X(_08326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14630_ (.A(_08326_),
    .Y(_08327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14631_ (.A(_08327_),
    .X(_08328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14632_ (.A(_08328_),
    .X(_08329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14633_ (.A(_08326_),
    .X(_08330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14634_ (.A1(\design_top.IOMUX[3][31] ),
    .A2(_08329_),
    .B1(\design_top.DATAO[31] ),
    .B2(_08330_),
    .C1(_10873_),
    .X(_05901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14635_ (.A(_08328_),
    .X(_08331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14636_ (.A(_08326_),
    .X(_08332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14637_ (.A(_08332_),
    .X(_08333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14638_ (.A1(\design_top.IOMUX[3][30] ),
    .A2(_08331_),
    .B1(\design_top.DATAO[30] ),
    .B2(_08333_),
    .C1(_10873_),
    .X(_05900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14639_ (.A1(\design_top.IOMUX[3][29] ),
    .A2(_08331_),
    .B1(\design_top.DATAO[29] ),
    .B2(_08333_),
    .C1(_10873_),
    .X(_05899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14640_ (.A1(\design_top.IOMUX[3][28] ),
    .A2(_08331_),
    .B1(\design_top.DATAO[28] ),
    .B2(_08333_),
    .C1(_10873_),
    .X(_05898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14641_ (.A(_10872_),
    .X(_08334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14642_ (.A1(\design_top.IOMUX[3][27] ),
    .A2(_08331_),
    .B1(\design_top.DATAO[27] ),
    .B2(_08333_),
    .C1(_08334_),
    .X(_05897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14643_ (.A1(\design_top.IOMUX[3][26] ),
    .A2(_08331_),
    .B1(\design_top.DATAO[26] ),
    .B2(_08333_),
    .C1(_08334_),
    .X(_05896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14644_ (.A(_08328_),
    .X(_08335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14645_ (.A(_08332_),
    .X(_08336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14646_ (.A1(\design_top.IOMUX[3][25] ),
    .A2(_08335_),
    .B1(\design_top.DATAO[25] ),
    .B2(_08336_),
    .C1(_08334_),
    .X(_05895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14647_ (.A1(\design_top.IOMUX[3][24] ),
    .A2(_08335_),
    .B1(\design_top.DATAO[24] ),
    .B2(_08336_),
    .C1(_08334_),
    .X(_05894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14648_ (.A1(\design_top.IOMUX[3][23] ),
    .A2(_08335_),
    .B1(\design_top.DATAO[23] ),
    .B2(_08336_),
    .C1(_08334_),
    .X(_05893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14649_ (.A(_10872_),
    .X(_08337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14650_ (.A1(\design_top.IOMUX[3][22] ),
    .A2(_08335_),
    .B1(\design_top.DATAO[22] ),
    .B2(_08336_),
    .C1(_08337_),
    .X(_05892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14651_ (.A1(\design_top.IOMUX[3][21] ),
    .A2(_08335_),
    .B1(\design_top.DATAO[21] ),
    .B2(_08336_),
    .C1(_08337_),
    .X(_05891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14652_ (.A(_08327_),
    .X(_08338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14653_ (.A(_08332_),
    .X(_08339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14654_ (.A1(\design_top.IOMUX[3][20] ),
    .A2(_08338_),
    .B1(\design_top.DATAO[20] ),
    .B2(_08339_),
    .C1(_08337_),
    .X(_05890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14655_ (.A1(\design_top.IOMUX[3][19] ),
    .A2(_08338_),
    .B1(\design_top.DATAO[19] ),
    .B2(_08339_),
    .C1(_08337_),
    .X(_05889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14656_ (.A1(\design_top.IOMUX[3][18] ),
    .A2(_08338_),
    .B1(\design_top.DATAO[18] ),
    .B2(_08339_),
    .C1(_08337_),
    .X(_05888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14657_ (.A(_10832_),
    .X(_08340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14658_ (.A1(\design_top.IOMUX[3][17] ),
    .A2(_08338_),
    .B1(\design_top.DATAO[17] ),
    .B2(_08339_),
    .C1(_08340_),
    .X(_05887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14659_ (.A1(\design_top.IOMUX[3][16] ),
    .A2(_08338_),
    .B1(\design_top.DATAO[16] ),
    .B2(_08339_),
    .C1(_08340_),
    .X(_05886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14660_ (.A(_08327_),
    .X(_08341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14661_ (.A(_08326_),
    .X(_08342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14662_ (.A1(\design_top.IOMUX[3][15] ),
    .A2(_08341_),
    .B1(\design_top.DATAO[15] ),
    .B2(_08342_),
    .C1(_08340_),
    .X(_05885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14663_ (.A1(\design_top.IOMUX[3][14] ),
    .A2(_08341_),
    .B1(\design_top.DATAO[14] ),
    .B2(_08342_),
    .C1(_08340_),
    .X(_05884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14664_ (.A1(\design_top.IOMUX[3][13] ),
    .A2(_08341_),
    .B1(\design_top.DATAO[13] ),
    .B2(_08342_),
    .C1(_08340_),
    .X(_05883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14665_ (.A(_10832_),
    .X(_08343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14666_ (.A1(\design_top.IOMUX[3][12] ),
    .A2(_08341_),
    .B1(\design_top.DATAO[12] ),
    .B2(_08342_),
    .C1(_08343_),
    .X(_05882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14667_ (.A1(\design_top.IOMUX[3][11] ),
    .A2(_08341_),
    .B1(\design_top.DATAO[11] ),
    .B2(_08342_),
    .C1(_08343_),
    .X(_05881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14668_ (.A(_08327_),
    .X(_08344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14669_ (.A(_08326_),
    .X(_08345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14670_ (.A1(\design_top.IOMUX[3][10] ),
    .A2(_08344_),
    .B1(\design_top.DATAO[10] ),
    .B2(_08345_),
    .C1(_08343_),
    .X(_05880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14671_ (.A1(\design_top.IOMUX[3][9] ),
    .A2(_08344_),
    .B1(\design_top.DATAO[9] ),
    .B2(_08345_),
    .C1(_08343_),
    .X(_05879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14672_ (.A1(\design_top.IOMUX[3][8] ),
    .A2(_08344_),
    .B1(\design_top.DATAO[8] ),
    .B2(_08345_),
    .C1(_08343_),
    .X(_05878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14673_ (.A(_10832_),
    .X(_08346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14674_ (.A1(\design_top.IOMUX[3][7] ),
    .A2(_08344_),
    .B1(\design_top.DATAO[7] ),
    .B2(_08345_),
    .C1(_08346_),
    .X(_05877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14675_ (.A(\design_top.IRES[7] ),
    .X(_08347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14676_ (.A(_08347_),
    .X(_08348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a221o_2 _14677_ (.A1(\design_top.DATAO[6] ),
    .A2(_08329_),
    .B1(\design_top.IOMUX[3][6] ),
    .B2(_08330_),
    .C1(_08348_),
    .X(_05876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a221o_2 _14678_ (.A1(\design_top.DATAO[5] ),
    .A2(_08329_),
    .B1(\design_top.IOMUX[3][5] ),
    .B2(_08330_),
    .C1(_08348_),
    .X(_05875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14679_ (.A1(\design_top.IOMUX[3][4] ),
    .A2(_08344_),
    .B1(\design_top.DATAO[4] ),
    .B2(_08345_),
    .C1(_08346_),
    .X(_05874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14680_ (.A1(\design_top.IOMUX[3][3] ),
    .A2(_08328_),
    .B1(\design_top.DATAO[3] ),
    .B2(_08332_),
    .C1(_08346_),
    .X(_05873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14681_ (.A1(\design_top.IOMUX[3][2] ),
    .A2(_08328_),
    .B1(\design_top.DATAO[2] ),
    .B2(_08332_),
    .C1(_08346_),
    .X(_05872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a221o_2 _14682_ (.A1(\design_top.DATAO[1] ),
    .A2(_08329_),
    .B1(\design_top.IOMUX[3][1] ),
    .B2(_08330_),
    .C1(_08347_),
    .X(_05871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a221o_2 _14683_ (.A1(\design_top.DATAO[0] ),
    .A2(_08329_),
    .B1(\design_top.IOMUX[3][0] ),
    .B2(_08330_),
    .C1(_08347_),
    .X(_05870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14684_ (.A(\design_top.core0.XRES ),
    .X(_08349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14685_ (.A(_08349_),
    .X(_08350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14686_ (.A(\design_top.IDATA[31] ),
    .Y(_08351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14687_ (.A(_10594_),
    .X(_08352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14688_ (.A(_08352_),
    .X(_08353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14689_ (.A(_03270_),
    .Y(_08354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14690_ (.A(_08354_),
    .B(_03271_),
    .C(_03272_),
    .X(_08355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14691_ (.A(io_out[21]),
    .B(io_out[20]),
    .Y(_08356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _14692_ (.A(io_out[23]),
    .B(_08356_),
    .C_N(io_out[22]),
    .X(_08357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14693_ (.A(_08355_),
    .B(_08357_),
    .Y(_08358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14694_ (.A(_03271_),
    .Y(_08359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14695_ (.A(_08354_),
    .B(_08359_),
    .C(_03272_),
    .X(_08360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14696_ (.A(_08357_),
    .B(_08360_),
    .Y(_08361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14697_ (.A(_08358_),
    .B(_08361_),
    .X(_08362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14698_ (.A(_08362_),
    .Y(_08363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14699_ (.A(_08363_),
    .X(_03914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14700_ (.A(\design_top.core0.UIMM[31] ),
    .Y(_08364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14701_ (.A(_10593_),
    .X(_08365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14702_ (.A(_08365_),
    .X(_08366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14703_ (.A(_08366_),
    .X(_08367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _14704_ (.A1(_08351_),
    .A2(_08353_),
    .A3(_03914_),
    .B1(_08364_),
    .B2(_08367_),
    .X(_08368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14705_ (.A(_08350_),
    .B(_08368_),
    .Y(_05869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14706_ (.A(_10594_),
    .X(_08369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14707_ (.A(_08369_),
    .X(_08370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14708_ (.A(_08370_),
    .X(_08371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14709_ (.A(_08371_),
    .X(\design_top.HLT ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14710_ (.A(\design_top.IDATA[30] ),
    .Y(_08372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14711_ (.A(\design_top.core0.UIMM[30] ),
    .Y(_08373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14712_ (.A(_08366_),
    .X(_08374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _14713_ (.A1(_08372_),
    .A2(_08353_),
    .A3(_03914_),
    .B1(_08373_),
    .B2(_08374_),
    .X(_08375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14714_ (.A(_08350_),
    .B(_08375_),
    .Y(_05868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14715_ (.A(_08370_),
    .X(_08376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14716_ (.A(_00693_),
    .Y(_08377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14717_ (.A(_10594_),
    .B(_08363_),
    .X(_08378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14718_ (.A(_08378_),
    .X(_08379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14719_ (.A1_N(\design_top.core0.UIMM[29] ),
    .A2_N(_08376_),
    .B1(_08377_),
    .B2(_08379_),
    .X(_08380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14720_ (.A(_08350_),
    .B(_08380_),
    .Y(_05867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14721_ (.A(_03968_),
    .Y(_08381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14722_ (.A1_N(\design_top.core0.UIMM[28] ),
    .A2_N(_08376_),
    .B1(_08381_),
    .B2(_08379_),
    .X(_08382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14723_ (.A(_08350_),
    .B(_08382_),
    .Y(_05866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14724_ (.A(_03964_),
    .Y(_08383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14725_ (.A1_N(\design_top.core0.UIMM[27] ),
    .A2_N(_08376_),
    .B1(_08383_),
    .B2(_08379_),
    .X(_08384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14726_ (.A(_08350_),
    .B(_08384_),
    .Y(_05865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14727_ (.A(_08349_),
    .X(_08385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14728_ (.A(_08369_),
    .X(_08386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14729_ (.A(_08386_),
    .X(_08387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14730_ (.A(_03960_),
    .Y(_08388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14731_ (.A1_N(\design_top.core0.UIMM[26] ),
    .A2_N(_08387_),
    .B1(_08388_),
    .B2(_08379_),
    .X(_08389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14732_ (.A(_08385_),
    .B(_08389_),
    .Y(_05864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14733_ (.A(_03956_),
    .Y(_08390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14734_ (.A1_N(\design_top.core0.UIMM[25] ),
    .A2_N(_08387_),
    .B1(_08390_),
    .B2(_08379_),
    .X(_08391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14735_ (.A(_08385_),
    .B(_08391_),
    .Y(_05863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14736_ (.A(_03952_),
    .Y(_08392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14737_ (.A1_N(\design_top.core0.UIMM[24] ),
    .A2_N(_08387_),
    .B1(_08392_),
    .B2(_08378_),
    .X(_08393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14738_ (.A(_08385_),
    .B(_08393_),
    .Y(_05862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14739_ (.A(\design_top.IDATA[23] ),
    .Y(_08394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14740_ (.A(\design_top.core0.UIMM[23] ),
    .Y(_08395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _14741_ (.A1(_08394_),
    .A2(_08353_),
    .A3(_03914_),
    .B1(_08395_),
    .B2(_08374_),
    .X(_08396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14742_ (.A(_08385_),
    .B(_08396_),
    .Y(_05861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14743_ (.A(\design_top.IDATA[22] ),
    .Y(_08397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14744_ (.A(_08352_),
    .X(_08398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14745_ (.A(\design_top.core0.UIMM[22] ),
    .Y(_08399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _14746_ (.A1(_08397_),
    .A2(_08398_),
    .A3(_08363_),
    .B1(_08399_),
    .B2(_08374_),
    .X(_08400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14747_ (.A(_08385_),
    .B(_08400_),
    .Y(_05860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14748_ (.A(_08349_),
    .X(_08401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14749_ (.A(\design_top.IDATA[21] ),
    .Y(_08402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14750_ (.A(\design_top.core0.UIMM[21] ),
    .Y(_08403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _14751_ (.A1(_08402_),
    .A2(_08398_),
    .A3(_08363_),
    .B1(_08403_),
    .B2(_08374_),
    .X(_08404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14752_ (.A(_08401_),
    .B(_08404_),
    .Y(_05859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14753_ (.A(_00753_),
    .Y(_08405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14754_ (.A(io_out[22]),
    .B(io_out[23]),
    .C(_08356_),
    .X(_08406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31ai_2 _14755_ (.A1(_03270_),
    .A2(_08359_),
    .A3(_08406_),
    .B1(_08365_),
    .Y(_08407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14756_ (.A(_08407_),
    .X(_08408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14757_ (.A1_N(\design_top.core0.UIMM[20] ),
    .A2_N(_08387_),
    .B1(_08405_),
    .B2(_08408_),
    .X(_08409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14758_ (.A(_08401_),
    .B(_08409_),
    .Y(_05858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14759_ (.A(_00751_),
    .Y(_08410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14760_ (.A1_N(\design_top.core0.UIMM[19] ),
    .A2_N(_08387_),
    .B1(_08410_),
    .B2(_08408_),
    .X(_08411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14761_ (.A(_08401_),
    .B(_08411_),
    .Y(_05857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14762_ (.A(_08386_),
    .X(_08412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14763_ (.A(_00749_),
    .Y(_08413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14764_ (.A1_N(\design_top.core0.UIMM[18] ),
    .A2_N(_08412_),
    .B1(_08413_),
    .B2(_08408_),
    .X(_08414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14765_ (.A(_08401_),
    .B(_08414_),
    .Y(_05856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14766_ (.A(_00747_),
    .Y(_08415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14767_ (.A1_N(\design_top.core0.UIMM[17] ),
    .A2_N(_08412_),
    .B1(_08415_),
    .B2(_08408_),
    .X(_08416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14768_ (.A(_08401_),
    .B(_08416_),
    .Y(_05855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14769_ (.A(_08349_),
    .X(_08417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14770_ (.A(_00745_),
    .Y(_08418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14771_ (.A1_N(\design_top.core0.UIMM[16] ),
    .A2_N(_08412_),
    .B1(_08418_),
    .B2(_08408_),
    .X(_08419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14772_ (.A(_08417_),
    .B(_08419_),
    .Y(_05854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14773_ (.A(_00743_),
    .Y(_08420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14774_ (.A1_N(\design_top.core0.UIMM[15] ),
    .A2_N(_08412_),
    .B1(_08420_),
    .B2(_08407_),
    .X(_08421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14775_ (.A(_08417_),
    .B(_08421_),
    .Y(_05853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14776_ (.A(_00741_),
    .Y(_08422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14777_ (.A1_N(\design_top.core0.UIMM[14] ),
    .A2_N(_08412_),
    .B1(_08422_),
    .B2(_08407_),
    .X(_08423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14778_ (.A(_08417_),
    .B(_08423_),
    .Y(_05852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14779_ (.A(_00739_),
    .Y(_08424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14780_ (.A1_N(\design_top.core0.UIMM[13] ),
    .A2_N(_08371_),
    .B1(_08424_),
    .B2(_08407_),
    .X(_08425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14781_ (.A(_08417_),
    .B(_08425_),
    .Y(_05851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14782_ (.A(_00737_),
    .Y(_08426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14783_ (.A(_03272_),
    .Y(_08427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and4b_2 _14784_ (.A_N(_08406_),
    .B(_03271_),
    .C(_08427_),
    .D(_08354_),
    .X(_00010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14785_ (.A(_08369_),
    .B(_00010_),
    .X(_08428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14786_ (.A1_N(\design_top.core0.UIMM[12] ),
    .A2_N(_08371_),
    .B1(_08426_),
    .B2(_08428_),
    .X(_08429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14787_ (.A(_08417_),
    .B(_08429_),
    .Y(_05850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14788_ (.A(_08398_),
    .X(_08430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14789_ (.A(_08366_),
    .X(_08431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14790_ (.A(\design_top.core0.XRES ),
    .Y(_08432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14791_ (.A(_08432_),
    .X(_08433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14792_ (.A(_08433_),
    .X(_08434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14793_ (.A1(_00049_),
    .A2(_08430_),
    .B1(_10688_),
    .B2(_08431_),
    .C1(_08434_),
    .X(_05849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14794_ (.A(_08433_),
    .X(_08435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14795_ (.A(_08435_),
    .X(_08436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14796_ (.A1(_00048_),
    .A2(_08430_),
    .B1(\design_top.core0.SIMM[10] ),
    .B2(_08431_),
    .C1(_08436_),
    .X(_05848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14797_ (.A(\design_top.core0.SIMM[9] ),
    .X(_08437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14798_ (.A(_08365_),
    .X(_08438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14799_ (.A(_08438_),
    .X(_08439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14800_ (.A(_08439_),
    .X(_08440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14801_ (.A1(_00077_),
    .A2(_08430_),
    .B1(_08437_),
    .B2(_08440_),
    .C1(_08436_),
    .X(_05847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14802_ (.A(\design_top.core0.SIMM[8] ),
    .X(_08441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14803_ (.A1(_00076_),
    .A2(_08430_),
    .B1(_08441_),
    .B2(_08440_),
    .C1(_08436_),
    .X(_05846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14804_ (.A(_08398_),
    .X(_08442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14805_ (.A(\design_top.core0.SIMM[7] ),
    .X(_08443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14806_ (.A1(_00075_),
    .A2(_08442_),
    .B1(_08443_),
    .B2(_08440_),
    .C1(_08436_),
    .X(_05845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14807_ (.A(\design_top.core0.SIMM[6] ),
    .X(_08444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14808_ (.A1(_00074_),
    .A2(_08442_),
    .B1(_08444_),
    .B2(_08440_),
    .C1(_08436_),
    .X(_05844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14809_ (.A(\design_top.core0.SIMM[5] ),
    .X(_08445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14810_ (.A(_08435_),
    .X(_08446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14811_ (.A1(_00073_),
    .A2(_08442_),
    .B1(_08445_),
    .B2(_08440_),
    .C1(_08446_),
    .X(_05843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14812_ (.A(\design_top.core0.SIMM[4] ),
    .X(_08447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14813_ (.A(_08439_),
    .X(_08448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14814_ (.A1(_00072_),
    .A2(_08442_),
    .B1(_08447_),
    .B2(_08448_),
    .C1(_08446_),
    .X(_05842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14815_ (.A1(_00071_),
    .A2(_08442_),
    .B1(_10702_),
    .B2(_08448_),
    .C1(_08446_),
    .X(_05841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14816_ (.A(_08352_),
    .X(_08449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14817_ (.A(_08449_),
    .X(_08450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14818_ (.A1(_00069_),
    .A2(_08450_),
    .B1(_10706_),
    .B2(_08448_),
    .C1(_08446_),
    .X(_05840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14819_ (.A1(_00058_),
    .A2(_08450_),
    .B1(_10709_),
    .B2(_08448_),
    .C1(_08446_),
    .X(_05839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14820_ (.A(_08435_),
    .X(_08451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14821_ (.A1(_00047_),
    .A2(_08450_),
    .B1(\design_top.core0.SIMM[0] ),
    .B2(_08448_),
    .C1(_08451_),
    .X(_05838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14822_ (.A(_08349_),
    .X(_08452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14823_ (.A1(_08351_),
    .A2(_08371_),
    .B1(_00780_),
    .B2(_08367_),
    .X(_08453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14824_ (.A(_08452_),
    .B(_08453_),
    .Y(_05837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14825_ (.A(_08439_),
    .X(_08454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14826_ (.A1(_00070_),
    .A2(_08450_),
    .B1(\design_top.core0.SIMM[30] ),
    .B2(_08454_),
    .C1(_08451_),
    .X(_05836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14827_ (.A1(_00068_),
    .A2(_08450_),
    .B1(_10600_),
    .B2(_08454_),
    .C1(_08451_),
    .X(_05835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14828_ (.A(_08449_),
    .X(_08455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14829_ (.A1(_00067_),
    .A2(_08455_),
    .B1(_10605_),
    .B2(_08454_),
    .C1(_08451_),
    .X(_05834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14830_ (.A1(_00066_),
    .A2(_08455_),
    .B1(\design_top.core0.SIMM[27] ),
    .B2(_08454_),
    .C1(_08451_),
    .X(_05833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14831_ (.A(_08435_),
    .X(_08456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14832_ (.A1(_00065_),
    .A2(_08455_),
    .B1(\design_top.core0.SIMM[26] ),
    .B2(_08454_),
    .C1(_08456_),
    .X(_05832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14833_ (.A(\design_top.core0.SIMM[25] ),
    .X(_08457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14834_ (.A(_08365_),
    .X(_08458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14835_ (.A(_08458_),
    .X(_08459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14836_ (.A1(_00064_),
    .A2(_08455_),
    .B1(_08457_),
    .B2(_08459_),
    .C1(_08456_),
    .X(_05831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14837_ (.A(\design_top.core0.SIMM[24] ),
    .X(_08460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14838_ (.A1(_00063_),
    .A2(_08455_),
    .B1(_08460_),
    .B2(_08459_),
    .C1(_08456_),
    .X(_05830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14839_ (.A(_08449_),
    .X(_08461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14840_ (.A1(_00062_),
    .A2(_08461_),
    .B1(_10750_),
    .B2(_08459_),
    .C1(_08456_),
    .X(_05829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14841_ (.A1(_00061_),
    .A2(_08461_),
    .B1(_10634_),
    .B2(_08459_),
    .C1(_08456_),
    .X(_05828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14842_ (.A(\design_top.core0.SIMM[21] ),
    .X(_08462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14843_ (.A(_08435_),
    .X(_08463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14844_ (.A1(_00060_),
    .A2(_08461_),
    .B1(_08462_),
    .B2(_08459_),
    .C1(_08463_),
    .X(_05827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14845_ (.A(_08458_),
    .X(_08464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14846_ (.A1(_00059_),
    .A2(_08461_),
    .B1(_10625_),
    .B2(_08464_),
    .C1(_08463_),
    .X(_05826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14847_ (.A1(_00057_),
    .A2(_08461_),
    .B1(_10653_),
    .B2(_08464_),
    .C1(_08463_),
    .X(_05825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14848_ (.A(_08449_),
    .X(_08465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14849_ (.A1(_00056_),
    .A2(_08465_),
    .B1(\design_top.core0.SIMM[18] ),
    .B2(_08464_),
    .C1(_08463_),
    .X(_05824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14850_ (.A(\design_top.core0.SIMM[17] ),
    .X(_08466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14851_ (.A1(_00055_),
    .A2(_08465_),
    .B1(_08466_),
    .B2(_08464_),
    .C1(_08463_),
    .X(_05823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14852_ (.A(\design_top.core0.SIMM[16] ),
    .X(_08467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14853_ (.A(_08433_),
    .X(_08468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14854_ (.A(_08468_),
    .X(_08469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14855_ (.A1(_00054_),
    .A2(_08465_),
    .B1(_08467_),
    .B2(_08464_),
    .C1(_08469_),
    .X(_05822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14856_ (.A(_08458_),
    .X(_08470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14857_ (.A1(_00053_),
    .A2(_08465_),
    .B1(_10735_),
    .B2(_08470_),
    .C1(_08469_),
    .X(_05821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14858_ (.A1(_00052_),
    .A2(_08465_),
    .B1(_10663_),
    .B2(_08470_),
    .C1(_08469_),
    .X(_05820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14859_ (.A(_08449_),
    .X(_08471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14860_ (.A(\design_top.core0.SIMM[13] ),
    .X(_08472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14861_ (.A1(_00051_),
    .A2(_08471_),
    .B1(_08472_),
    .B2(_08470_),
    .C1(_08469_),
    .X(_05819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14862_ (.A1(_00050_),
    .A2(_08471_),
    .B1(_10671_),
    .B2(_08470_),
    .C1(_08469_),
    .X(_05818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14863_ (.A(_08352_),
    .X(_08473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14864_ (.A(_08406_),
    .X(_08474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14865_ (.A(\design_top.core0.XRCC ),
    .Y(_08475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _14866_ (.A1(_08473_),
    .A2(_08474_),
    .A3(_08360_),
    .B1(_08475_),
    .B2(_08374_),
    .X(_08476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14867_ (.A(_08452_),
    .B(_08476_),
    .Y(_05817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14868_ (.A(\design_top.core0.XMCC ),
    .Y(_08477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14869_ (.A(_08438_),
    .X(_08478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _14870_ (.A1(_08473_),
    .A2(_08474_),
    .A3(_08355_),
    .B1(_08477_),
    .B2(_08478_),
    .X(_08479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14871_ (.A(_08452_),
    .B(_08479_),
    .Y(_05816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14872_ (.A(_08433_),
    .X(_08480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _14873_ (.A1(\design_top.core0.XSCC ),
    .A2(_08431_),
    .B1(_08480_),
    .C1(_08428_),
    .X(_05815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and4b_2 _14874_ (.A_N(_08474_),
    .B(_08427_),
    .C(_08354_),
    .D(_08359_),
    .X(_08481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14875_ (.A(_08480_),
    .X(_08482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14876_ (.A1(\design_top.HLT ),
    .A2(_08481_),
    .B1(_08482_),
    .X(_05814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14877_ (.A(_03270_),
    .B(_08359_),
    .C(_08427_),
    .X(_08483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14878_ (.A(\design_top.core0.XBCC ),
    .Y(_08484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _14879_ (.A1(_08473_),
    .A2(_08474_),
    .A3(_08483_),
    .B1(_08484_),
    .B2(_08478_),
    .X(_08485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14880_ (.A(_08452_),
    .B(_08485_),
    .Y(_05813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14881_ (.A(_08474_),
    .B(_08483_),
    .Y(_00009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14882_ (.A(\design_top.core0.XJALR ),
    .Y(_08486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _14883_ (.A1(_08473_),
    .A2(_08483_),
    .A3(_08357_),
    .B1(_08486_),
    .B2(_08478_),
    .X(_08487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14884_ (.A(_08452_),
    .B(_08487_),
    .Y(_05812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14885_ (.A(_08366_),
    .X(_08488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14886_ (.A(_08398_),
    .X(_08489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and4bb_2 _14887_ (.A_N(_08483_),
    .B_N(_08356_),
    .C(io_out[23]),
    .D(io_out[22]),
    .X(_00008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14888_ (.A(_08468_),
    .X(_08490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14889_ (.A1(\design_top.core0.XJAL ),
    .A2(_08488_),
    .B1(_08489_),
    .B2(_00008_),
    .C1(_08490_),
    .X(_05811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14890_ (.A1(\design_top.core0.XAUIPC ),
    .A2(_08488_),
    .B1(_08489_),
    .B2(_08358_),
    .C1(_08490_),
    .X(_05810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14891_ (.A1(\design_top.core0.XLUI ),
    .A2(_08488_),
    .B1(_08430_),
    .B2(_08361_),
    .C1(_08490_),
    .X(_05809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14892_ (.A(\design_top.core0.XRES ),
    .X(_08491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14893_ (.A(\design_top.core0.FCT7[5] ),
    .Y(_08492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14894_ (.A1(_08372_),
    .A2(_08371_),
    .B1(_08492_),
    .B2(_08367_),
    .X(_08493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14895_ (.A(_08491_),
    .B(_08493_),
    .Y(_05808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14896_ (.A(_08386_),
    .X(_08494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22oi_2 _14897_ (.A1(\design_top.IDATA[23] ),
    .A2(_08488_),
    .B1(\design_top.core0.S2PTR[3] ),
    .B2(_08494_),
    .Y(_08495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14898_ (.A(_08491_),
    .B(_08495_),
    .Y(_05807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22oi_2 _14899_ (.A1(\design_top.IDATA[22] ),
    .A2(_08367_),
    .B1(\design_top.core0.S2PTR[2] ),
    .B2(_08376_),
    .Y(_08496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14900_ (.A(_08491_),
    .B(_08496_),
    .Y(_05806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22oi_2 _14901_ (.A1(\design_top.IDATA[21] ),
    .A2(_08367_),
    .B1(\design_top.core0.S2PTR[1] ),
    .B2(_08376_),
    .Y(_08497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14902_ (.A(_08491_),
    .B(_08497_),
    .Y(_05805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14903_ (.A1(\design_top.IDATA[20] ),
    .A2(_08471_),
    .B1(\design_top.core0.S2PTR[0] ),
    .B2(_08470_),
    .C1(_08490_),
    .X(_05804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14904_ (.A(_08458_),
    .X(_08498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14905_ (.A1(\design_top.IDATA[18] ),
    .A2(_08471_),
    .B1(\design_top.core0.S1PTR[3] ),
    .B2(_08498_),
    .C1(_08490_),
    .X(_05803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14906_ (.A(_08468_),
    .X(_08499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14907_ (.A1(\design_top.IDATA[17] ),
    .A2(_08471_),
    .B1(\design_top.core0.S1PTR[2] ),
    .B2(_08498_),
    .C1(_08499_),
    .X(_05802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14908_ (.A(_08352_),
    .X(_08500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14909_ (.A(_08500_),
    .X(_08501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14910_ (.A1(\design_top.IDATA[16] ),
    .A2(_08501_),
    .B1(\design_top.core0.S1PTR[1] ),
    .B2(_08498_),
    .C1(_08499_),
    .X(_05801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14911_ (.A1(\design_top.IDATA[15] ),
    .A2(_08501_),
    .B1(\design_top.core0.S1PTR[0] ),
    .B2(_08498_),
    .C1(_08499_),
    .X(_05800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14912_ (.A1(\design_top.IDATA[14] ),
    .A2(_08501_),
    .B1(\design_top.core0.FCT3[2] ),
    .B2(_08498_),
    .C1(_08499_),
    .X(_05799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14913_ (.A(\design_top.core0.FCT3[1] ),
    .X(_08502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14914_ (.A(_08458_),
    .X(_08503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14915_ (.A1(\design_top.IDATA[13] ),
    .A2(_08501_),
    .B1(_08502_),
    .B2(_08503_),
    .C1(_08499_),
    .X(_05798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14916_ (.A(_08468_),
    .X(_08504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14917_ (.A1(\design_top.IDATA[12] ),
    .A2(_08501_),
    .B1(\design_top.core0.FCT3[0] ),
    .B2(_08503_),
    .C1(_08504_),
    .X(_05797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14918_ (.A(_08500_),
    .X(_08505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14919_ (.A1(\design_top.IDATA[10] ),
    .A2(_08505_),
    .B1(\design_top.core0.XIDATA[10] ),
    .B2(_08503_),
    .C1(_08504_),
    .X(_05796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14920_ (.A1(\design_top.IDATA[9] ),
    .A2(_08505_),
    .B1(\design_top.core0.XIDATA[9] ),
    .B2(_08503_),
    .C1(_08504_),
    .X(_05795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14921_ (.A1(\design_top.IDATA[8] ),
    .A2(_08505_),
    .B1(\design_top.core0.XIDATA[8] ),
    .B2(_08503_),
    .C1(_08504_),
    .X(_05794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14922_ (.A(_08365_),
    .X(_08506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14923_ (.A(_08506_),
    .X(_08507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14924_ (.A1(\design_top.IDATA[7] ),
    .A2(_08505_),
    .B1(\design_top.core0.XIDATA[7] ),
    .B2(_08507_),
    .C1(_08504_),
    .X(_05793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14925_ (.A(_08468_),
    .X(_08508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14926_ (.A1(_00101_),
    .A2(_08505_),
    .B1(\design_top.IADDR[31] ),
    .B2(_08507_),
    .C1(_08508_),
    .X(_05792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14927_ (.A(_08500_),
    .X(_08509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14928_ (.A1(_00100_),
    .A2(_08509_),
    .B1(\design_top.IADDR[30] ),
    .B2(_08507_),
    .C1(_08508_),
    .X(_05791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14929_ (.A1(_00098_),
    .A2(_08509_),
    .B1(\design_top.IADDR[29] ),
    .B2(_08507_),
    .C1(_08508_),
    .X(_05790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14930_ (.A1(_00097_),
    .A2(_08509_),
    .B1(\design_top.IADDR[28] ),
    .B2(_08507_),
    .C1(_08508_),
    .X(_05789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14931_ (.A(_08506_),
    .X(_08510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14932_ (.A1(_00096_),
    .A2(_08509_),
    .B1(\design_top.IADDR[27] ),
    .B2(_08510_),
    .C1(_08508_),
    .X(_05788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14933_ (.A(_08433_),
    .X(_08511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14934_ (.A(_08511_),
    .X(_08512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14935_ (.A1(_00095_),
    .A2(_08509_),
    .B1(\design_top.IADDR[26] ),
    .B2(_08510_),
    .C1(_08512_),
    .X(_05787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14936_ (.A(_08500_),
    .X(_08513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14937_ (.A1(_00094_),
    .A2(_08513_),
    .B1(\design_top.IADDR[25] ),
    .B2(_08510_),
    .C1(_08512_),
    .X(_05786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14938_ (.A1(_00093_),
    .A2(_08513_),
    .B1(\design_top.IADDR[24] ),
    .B2(_08510_),
    .C1(_08512_),
    .X(_05785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14939_ (.A1(_00092_),
    .A2(_08513_),
    .B1(\design_top.IADDR[23] ),
    .B2(_08510_),
    .C1(_08512_),
    .X(_05784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14940_ (.A(_08506_),
    .X(_08514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14941_ (.A1(_00091_),
    .A2(_08513_),
    .B1(\design_top.IADDR[22] ),
    .B2(_08514_),
    .C1(_08512_),
    .X(_05783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14942_ (.A(_08511_),
    .X(_08515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14943_ (.A1(_00090_),
    .A2(_08513_),
    .B1(\design_top.IADDR[21] ),
    .B2(_08514_),
    .C1(_08515_),
    .X(_05782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14944_ (.A(_08500_),
    .X(_08516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14945_ (.A1(_00089_),
    .A2(_08516_),
    .B1(\design_top.IADDR[20] ),
    .B2(_08514_),
    .C1(_08515_),
    .X(_05781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14946_ (.A1(_00088_),
    .A2(_08516_),
    .B1(\design_top.IADDR[19] ),
    .B2(_08514_),
    .C1(_08515_),
    .X(_05780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14947_ (.A1(_00087_),
    .A2(_08516_),
    .B1(\design_top.IADDR[18] ),
    .B2(_08514_),
    .C1(_08515_),
    .X(_05779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14948_ (.A(_08506_),
    .X(_08517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14949_ (.A1(_00086_),
    .A2(_08516_),
    .B1(\design_top.IADDR[17] ),
    .B2(_08517_),
    .C1(_08515_),
    .X(_05778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14950_ (.A(_08511_),
    .X(_08518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14951_ (.A1(_00085_),
    .A2(_08516_),
    .B1(\design_top.IADDR[16] ),
    .B2(_08517_),
    .C1(_08518_),
    .X(_05777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14952_ (.A(_08386_),
    .X(_08519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14953_ (.A1(_00084_),
    .A2(_08519_),
    .B1(\design_top.IADDR[15] ),
    .B2(_08517_),
    .C1(_08518_),
    .X(_05776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14954_ (.A1(_00083_),
    .A2(_08519_),
    .B1(\design_top.IADDR[14] ),
    .B2(_08517_),
    .C1(_08518_),
    .X(_05775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14955_ (.A1(_00082_),
    .A2(_08519_),
    .B1(\design_top.IADDR[13] ),
    .B2(_08517_),
    .C1(_08518_),
    .X(_05774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14956_ (.A(_08506_),
    .X(_08520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14957_ (.A1(_00081_),
    .A2(_08519_),
    .B1(\design_top.IADDR[12] ),
    .B2(_08520_),
    .C1(_08518_),
    .X(_05773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14958_ (.A(_08511_),
    .X(_08521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14959_ (.A1(_00080_),
    .A2(_08519_),
    .B1(\design_top.IADDR[11] ),
    .B2(_08520_),
    .C1(_08521_),
    .X(_05772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14960_ (.A(_08386_),
    .X(_08522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14961_ (.A1(_00079_),
    .A2(_08522_),
    .B1(\design_top.IADDR[10] ),
    .B2(_08520_),
    .C1(_08521_),
    .X(_05771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14962_ (.A1(_00108_),
    .A2(_08522_),
    .B1(\design_top.IADDR[9] ),
    .B2(_08520_),
    .C1(_08521_),
    .X(_05770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14963_ (.A1(_00107_),
    .A2(_08522_),
    .B1(\design_top.IADDR[8] ),
    .B2(_08520_),
    .C1(_08521_),
    .X(_05769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14964_ (.A(_08366_),
    .X(_08523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14965_ (.A1(_00106_),
    .A2(_08522_),
    .B1(\design_top.IADDR[7] ),
    .B2(_08523_),
    .C1(_08521_),
    .X(_05768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14966_ (.A(_08511_),
    .X(_08524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14967_ (.A1(_00105_),
    .A2(_08522_),
    .B1(\design_top.IADDR[6] ),
    .B2(_08523_),
    .C1(_08524_),
    .X(_05767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14968_ (.A1(_00104_),
    .A2(_08494_),
    .B1(\design_top.IADDR[5] ),
    .B2(_08523_),
    .C1(_08524_),
    .X(_05766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14969_ (.A(\design_top.IADDR[4] ),
    .X(_08525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14970_ (.A1(_00103_),
    .A2(_08494_),
    .B1(_08525_),
    .B2(_08523_),
    .C1(_08524_),
    .X(_05765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14971_ (.A1(_00102_),
    .A2(_08494_),
    .B1(io_out[19]),
    .B2(_08523_),
    .C1(_08524_),
    .X(_05764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14972_ (.A1(_00099_),
    .A2(_08494_),
    .B1(io_out[18]),
    .B2(_08488_),
    .C1(_08524_),
    .X(_05763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14973_ (.A(_08478_),
    .X(_08526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _14974_ (.A1(_00011_),
    .A2(_08526_),
    .B1(_08491_),
    .X(_05762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _14975_ (.A(_08480_),
    .B(\design_top.core0.FLUSH[1] ),
    .C(_10591_),
    .X(_05761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14976_ (.A(\design_top.core0.XJAL ),
    .Y(_08527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14977_ (.A(_03194_),
    .Y(_08528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14978_ (.A(_02945_),
    .B(_10638_),
    .Y(_02947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14979_ (.A(_02945_),
    .B(_10638_),
    .X(_08529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14980_ (.A(_02947_),
    .B(_08529_),
    .Y(_03180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14981_ (.A(_03180_),
    .Y(_08530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14982_ (.A(_10629_),
    .X(_08531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14983_ (.A(_02962_),
    .B(_10629_),
    .Y(_02964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14984_ (.A1(_02962_),
    .A2(_08531_),
    .B1(_02964_),
    .Y(_03178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14985_ (.A(_03178_),
    .Y(_08532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14986_ (.A(_02749_),
    .X(_08533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14987_ (.A(_02971_),
    .B(_08533_),
    .Y(_01601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14988_ (.A1(_02971_),
    .A2(_08533_),
    .B1(_01601_),
    .Y(_08534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14989_ (.A(_08534_),
    .Y(_08535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14990_ (.A(_02954_),
    .B(_10635_),
    .Y(_01643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14991_ (.A1(_02954_),
    .A2(_10635_),
    .B1(_01643_),
    .Y(_08536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14992_ (.A(_08536_),
    .Y(_08537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _14993_ (.A(_08530_),
    .B(_08532_),
    .C(_08535_),
    .D(_08537_),
    .X(_08538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14994_ (.A(_10650_),
    .X(_08539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14995_ (.A(_02996_),
    .B(_10650_),
    .Y(_02998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14996_ (.A1(_02996_),
    .A2(_08539_),
    .B1(_02998_),
    .Y(_03175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14997_ (.A(_03175_),
    .Y(_08540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14998_ (.A(_02755_),
    .X(_08541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14999_ (.A(_02979_),
    .B(_02755_),
    .Y(_02981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15000_ (.A1(_02979_),
    .A2(_08541_),
    .B1(_02981_),
    .Y(_03176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15001_ (.A(_03176_),
    .Y(_08542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15002_ (.A(_02988_),
    .B(_02761_),
    .Y(_01559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15003_ (.A(_01559_),
    .Y(_08543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15004_ (.A(_02988_),
    .B(_02761_),
    .Y(_02989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15005_ (.A(_08543_),
    .B(_02989_),
    .X(_08544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15006_ (.A(_08544_),
    .Y(_08545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15007_ (.A(_02773_),
    .X(_08546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15008_ (.A(_03005_),
    .B(_08546_),
    .Y(_01517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15009_ (.A1(_03005_),
    .A2(_08546_),
    .B1(_01517_),
    .Y(_03174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15010_ (.A(_03174_),
    .Y(_08547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _15011_ (.A(_08540_),
    .B(_08542_),
    .C(_08545_),
    .D(_08547_),
    .X(_08548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15012_ (.A(_02707_),
    .X(_08549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15013_ (.A(_02911_),
    .B(_08549_),
    .Y(_02913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15014_ (.A1(_02911_),
    .A2(_08549_),
    .B1(_02913_),
    .Y(_03184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15015_ (.A(_03184_),
    .Y(_08550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15016_ (.A(_10610_),
    .X(_08551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15017_ (.A(_02928_),
    .B(_10610_),
    .Y(_02930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15018_ (.A1(_02928_),
    .A2(_08551_),
    .B1(_02930_),
    .Y(_03182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15019_ (.A(_03182_),
    .Y(_08552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15020_ (.A(_02725_),
    .X(_08553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15021_ (.A(_02937_),
    .B(_08553_),
    .Y(_01683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15022_ (.A1(_02937_),
    .A2(_08553_),
    .B1(_01683_),
    .Y(_08554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15023_ (.A(_02920_),
    .B(_10619_),
    .Y(_01725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15024_ (.A1(_02920_),
    .A2(_10619_),
    .B1(_01725_),
    .Y(_08555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15025_ (.A(_08554_),
    .B(_08555_),
    .Y(_08556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15026_ (.A(_02885_),
    .B(_02689_),
    .Y(_02887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15027_ (.A1(_02885_),
    .A2(_02689_),
    .B1(_02887_),
    .Y(_03187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15028_ (.A(_03187_),
    .Y(_08557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15029_ (.A(_10764_),
    .B(_02876_),
    .Y(_02877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _15030_ (.A1(_10764_),
    .A2(_02876_),
    .B1(_02877_),
    .Y(_08558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15031_ (.A(_02695_),
    .X(_08559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15032_ (.A(_02894_),
    .B(_02695_),
    .Y(_02896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15033_ (.A1(_02894_),
    .A2(_08559_),
    .B1(_02896_),
    .Y(_03186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15034_ (.A(_03186_),
    .Y(_08560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15035_ (.A(_02903_),
    .B(_02701_),
    .Y(_01766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15036_ (.A1(_02903_),
    .A2(_10606_),
    .B1(_01766_),
    .Y(_03185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15037_ (.A(_03185_),
    .Y(_08561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _15038_ (.A(_08557_),
    .B(_08558_),
    .C(_08560_),
    .D(_08561_),
    .X(_08562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _15039_ (.A(_08550_),
    .B(_08552_),
    .C(_08556_),
    .D(_08562_),
    .X(_08563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _15040_ (.A(_08538_),
    .B(_08548_),
    .C(_08563_),
    .X(_08564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15041_ (.A(_03022_),
    .B(_10664_),
    .Y(_01476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15042_ (.A1(_03022_),
    .A2(_10664_),
    .B1(_01476_),
    .Y(_08565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15043_ (.A(_08565_),
    .X(_01477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15044_ (.A(_01477_),
    .Y(_08566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15045_ (.A(_02791_),
    .X(_08567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15046_ (.A(_03030_),
    .B(_08567_),
    .Y(_03032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15047_ (.A1(_03030_),
    .A2(_08567_),
    .B1(_03032_),
    .Y(_03172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15048_ (.A(_03172_),
    .Y(_08568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15049_ (.A(_03120_),
    .Y(_08569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15050_ (.A1(_03120_),
    .A2(_02634_),
    .B1(_08569_),
    .B2(_10770_),
    .X(_08570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15051_ (.A(_03013_),
    .B(_10657_),
    .Y(_03015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15052_ (.A1(_03013_),
    .A2(_10657_),
    .B1(_03015_),
    .Y(_03173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15053_ (.A(_03173_),
    .Y(_08571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15054_ (.A(_03039_),
    .B(_10672_),
    .Y(_01428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15055_ (.A1(_03039_),
    .A2(_10672_),
    .B1(_01428_),
    .Y(_08572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15056_ (.A(_08572_),
    .Y(_08573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _15057_ (.A(_08570_),
    .B(_08571_),
    .C(_08573_),
    .X(_08574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15058_ (.A(_00688_),
    .Y(_08575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15059_ (.A1(_08575_),
    .A2(_02640_),
    .B1(_00688_),
    .B2(_02637_),
    .X(_08576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15060_ (.A(_03128_),
    .B(_08576_),
    .Y(_01010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _15061_ (.A1(_03128_),
    .A2(_08576_),
    .B1(_01010_),
    .Y(_08577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15062_ (.A(_08577_),
    .X(_08578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15063_ (.A(_03087_),
    .B(_10696_),
    .Y(_01268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15064_ (.A1(_03087_),
    .A2(_10696_),
    .B1(_01268_),
    .Y(_08579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15065_ (.A(_08579_),
    .Y(_08580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15066_ (.A(_10691_),
    .B(_03094_),
    .Y(_03095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _15067_ (.A1(_10691_),
    .A2(_03094_),
    .B1(_03095_),
    .Y(_08581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15068_ (.A(_03103_),
    .B(_10693_),
    .Y(_01181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15069_ (.A1(_03103_),
    .A2(_10693_),
    .B1(_01181_),
    .Y(_08582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15070_ (.A(_08582_),
    .Y(_08583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15071_ (.A(_02827_),
    .B(_03078_),
    .Y(_03079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _15072_ (.A1(_02827_),
    .A2(_03078_),
    .B1(_03079_),
    .Y(_08584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _15073_ (.A(_08580_),
    .B(_08581_),
    .C(_08583_),
    .D(_08584_),
    .X(_08585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15074_ (.A1(_08575_),
    .A2(_02658_),
    .B1(_00688_),
    .B2(_02655_),
    .X(_08586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15075_ (.A(_03111_),
    .B(_08586_),
    .Y(_03112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _15076_ (.A1(_03111_),
    .A2(_08586_),
    .B1(_03112_),
    .Y(_08587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15077_ (.A(_10676_),
    .B(_03046_),
    .X(_08588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15078_ (.A(_10676_),
    .B(_03046_),
    .Y(_03048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15079_ (.A(_08588_),
    .B(_03048_),
    .Y(_03170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15080_ (.A(_03170_),
    .Y(_08589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15081_ (.A(_02815_),
    .X(_08590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15082_ (.A(_08590_),
    .B(_03062_),
    .Y(_03063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _15083_ (.A1(_08590_),
    .A2(_03062_),
    .B1(_03063_),
    .Y(_08591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15084_ (.A(_03071_),
    .B(_10685_),
    .Y(_01337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15085_ (.A1(_03071_),
    .A2(_10685_),
    .B1(_01337_),
    .Y(_03167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15086_ (.A(_03167_),
    .Y(_08592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15087_ (.A(_03055_),
    .B(_10682_),
    .Y(_03056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15088_ (.A(_03055_),
    .B(_10682_),
    .Y(_01383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15089_ (.A(_01383_),
    .Y(_08593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15090_ (.A(_03056_),
    .B(_08593_),
    .X(_08594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15091_ (.A(_08594_),
    .Y(_08595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _15092_ (.A(_08589_),
    .B(_08591_),
    .C(_08592_),
    .D(_08595_),
    .X(_08596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _15093_ (.A(_08578_),
    .B(_08585_),
    .C(_08587_),
    .D(_08596_),
    .X(_08597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _15094_ (.A(_08566_),
    .B(_08568_),
    .C(_08574_),
    .D(_08597_),
    .X(_08598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15095_ (.A(\design_top.core0.FCT3[2] ),
    .Y(_08599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15096_ (.A(\design_top.core0.FCT3[1] ),
    .B(\design_top.core0.FCT3[0] ),
    .X(_08600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15097_ (.A(_08600_),
    .X(_02854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _15098_ (.A1(_08564_),
    .A2(_08598_),
    .B1(_08599_),
    .C1(_02854_),
    .X(_08601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15099_ (.A1(_08528_),
    .A2(_08601_),
    .B1(\design_top.core0.XBCC ),
    .Y(_08602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _15100_ (.A1(_08486_),
    .A2(_08527_),
    .A3(_08602_),
    .B1(_10595_),
    .X(_03195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15101_ (.A(_08369_),
    .B(_03195_),
    .X(_08603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15102_ (.A(_08603_),
    .Y(_08604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15103_ (.A(_01829_),
    .Y(_08605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _15104_ (.A1(io_out[17]),
    .A2(_08604_),
    .B1(_08605_),
    .B2(_08603_),
    .C1(_08480_),
    .X(_05760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15105_ (.A(_01828_),
    .Y(_08606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _15106_ (.A1(io_out[16]),
    .A2(_08604_),
    .B1(_08606_),
    .B2(_08603_),
    .C1(_08480_),
    .X(_05759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15107_ (.A(_10926_),
    .B(_08103_),
    .X(_08607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15108_ (.A(_08607_),
    .X(_08608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _15109_ (.A1(_10987_),
    .A2(_11138_),
    .B1(_08607_),
    .X(_08609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15110_ (.A(_08609_),
    .X(_08610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _15111_ (.A1_N(_10923_),
    .A2_N(_08608_),
    .B1(\design_top.MEM[9][31] ),
    .B2(_08610_),
    .X(_05758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _15112_ (.A1_N(_10933_),
    .A2_N(_08608_),
    .B1(\design_top.MEM[9][30] ),
    .B2(_08610_),
    .X(_05757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _15113_ (.A1_N(_10936_),
    .A2_N(_08608_),
    .B1(\design_top.MEM[9][29] ),
    .B2(_08610_),
    .X(_05756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _15114_ (.A1_N(_10939_),
    .A2_N(_08608_),
    .B1(\design_top.MEM[9][28] ),
    .B2(_08610_),
    .X(_05755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _15115_ (.A1_N(_10942_),
    .A2_N(_08608_),
    .B1(\design_top.MEM[9][27] ),
    .B2(_08610_),
    .X(_05754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _15116_ (.A1_N(_10945_),
    .A2_N(_08607_),
    .B1(\design_top.MEM[9][26] ),
    .B2(_08609_),
    .X(_05753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _15117_ (.A1_N(_10948_),
    .A2_N(_08607_),
    .B1(\design_top.MEM[9][25] ),
    .B2(_08609_),
    .X(_05752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _15118_ (.A1_N(_10951_),
    .A2_N(_08607_),
    .B1(\design_top.MEM[9][24] ),
    .B2(_08609_),
    .X(_05751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _15119_ (.A(_08482_),
    .B(_00003_),
    .X(_05750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _15120_ (.A(_08482_),
    .B(_00002_),
    .X(_05749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _15121_ (.A(_08482_),
    .B(_00001_),
    .X(_05748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _15122_ (.A(_08482_),
    .B(_00000_),
    .X(_05747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _15123_ (.A(_08434_),
    .B(_00007_),
    .X(_05746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _15124_ (.A(_08434_),
    .B(_00006_),
    .X(_05745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _15125_ (.A(_08434_),
    .B(_00005_),
    .X(_05744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _15126_ (.A(_08434_),
    .B(_00004_),
    .X(_05743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _15127_ (.A(_08346_),
    .B(\design_top.DACK[0] ),
    .C(\design_top.DACK[1] ),
    .X(_05742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _15128_ (.A(_10833_),
    .B(_00012_),
    .X(_05741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15129_ (.A(\design_top.uart0.UART_XSTATE[1] ),
    .X(_08611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15130_ (.A(\design_top.uart0.UART_XSTATE[0] ),
    .Y(_08612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15131_ (.A(_08612_),
    .B(_02624_),
    .Y(_08613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _15132_ (.A(_08611_),
    .B(_08613_),
    .C(\design_top.uart0.UART_XSTATE[2] ),
    .X(_08614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15133_ (.A(\design_top.uart0.UART_XSTATE[3] ),
    .Y(_08615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15134_ (.A(_08614_),
    .Y(_08616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15135_ (.A(_08611_),
    .Y(_08617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15136_ (.A(\design_top.uart0.UART_XSTATE[2] ),
    .Y(_08618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a41o_2 _15137_ (.A1(\design_top.uart0.UART_XSTATE[0] ),
    .A2(_08617_),
    .A3(_08615_),
    .A4(_08618_),
    .B1(_08347_),
    .X(_08619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15138_ (.A(_08619_),
    .Y(_08620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _15139_ (.A1(\design_top.uart0.UART_XSTATE[3] ),
    .A2(_08614_),
    .B1(_08615_),
    .B2(_08616_),
    .C1(_08620_),
    .X(_05740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _15140_ (.A1(_08611_),
    .A2(_08613_),
    .B1(\design_top.uart0.UART_XSTATE[2] ),
    .Y(_08621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15141_ (.A1(_08614_),
    .A2(_08621_),
    .B1(_08620_),
    .Y(_05739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _15142_ (.A1_N(_08611_),
    .A2_N(_08613_),
    .B1(_08611_),
    .B2(_08613_),
    .X(_08622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15143_ (.A(_08619_),
    .B(_08622_),
    .X(_05738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211oi_2 _15144_ (.A1(_08612_),
    .A2(_02624_),
    .B1(_08613_),
    .C1(_08619_),
    .Y(_05737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15145_ (.A(\design_top.uart0.UART_RSTATE[2] ),
    .Y(_08623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15146_ (.A(_08623_),
    .X(_08624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15147_ (.A(\design_top.uart0.UART_RSTATE[0] ),
    .Y(_08625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15148_ (.A(\design_top.uart0.UART_RSTATE[1] ),
    .Y(_08626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _15149_ (.A(_08625_),
    .B(_02626_),
    .C(_08626_),
    .X(_08627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15150_ (.A(\design_top.uart0.UART_RSTATE[3] ),
    .Y(_08628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15151_ (.A(_08628_),
    .X(_08629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15152_ (.A(\design_top.uart0.UART_RSTATE[1] ),
    .X(_08630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _15153_ (.A(_08625_),
    .B(_08630_),
    .C(\design_top.uart0.UART_RSTATE[3] ),
    .D(\design_top.uart0.UART_RSTATE[2] ),
    .X(_08631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15154_ (.A(_10832_),
    .B(_08631_),
    .Y(_08632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15155_ (.A(_08632_),
    .Y(_08633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15156_ (.A1(_08624_),
    .A2(_08627_),
    .B1(_08629_),
    .Y(_08634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o311a_2 _15157_ (.A1(_08624_),
    .A2(_08627_),
    .A3(_08629_),
    .B1(_08633_),
    .C1(_08634_),
    .X(_05736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15158_ (.A(\design_top.uart0.UART_RSTATE[2] ),
    .X(_08635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15159_ (.A(_08627_),
    .Y(_08636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15160_ (.A1(_08624_),
    .A2(_08627_),
    .B1(_08635_),
    .B2(_08636_),
    .X(_08637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15161_ (.A(_08632_),
    .B(_08637_),
    .X(_05735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15162_ (.A(_08625_),
    .X(_08638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15163_ (.A(_08626_),
    .X(_08639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _15164_ (.A1(_08638_),
    .A2(_02626_),
    .B1(_08639_),
    .X(_08640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15165_ (.A1(_08636_),
    .A2(_08640_),
    .B1(_08633_),
    .Y(_05734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15166_ (.A(\design_top.uart0.UART_RSTATE[0] ),
    .X(_08641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15167_ (.A(_02626_),
    .Y(_08642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _15168_ (.A1(_08638_),
    .A2(_02626_),
    .B1(_08641_),
    .B2(_08642_),
    .C1(_08633_),
    .X(_05733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _15169_ (.A(\design_top.uart0.UART_RSTATE[0] ),
    .B(_08626_),
    .C(\design_top.uart0.UART_RSTATE[3] ),
    .D(_08623_),
    .X(_08643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15170_ (.A(_08643_),
    .Y(_02662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15171_ (.A(\design_top.uart0.UART_RBAUD[1] ),
    .B(\design_top.uart0.UART_RBAUD[0] ),
    .X(_08644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _15172_ (.A(\design_top.uart0.UART_RBAUD[2] ),
    .B(_08644_),
    .C(\design_top.uart0.UART_RBAUD[3] ),
    .X(_08645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15173_ (.A(\design_top.uart0.UART_RBAUD[4] ),
    .B(_08645_),
    .X(_08646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15174_ (.A(\design_top.uart0.UART_RBAUD[5] ),
    .B(_08646_),
    .X(_08647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15175_ (.A(\design_top.uart0.UART_RBAUD[6] ),
    .B(_08647_),
    .X(_08648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15176_ (.A(\design_top.uart0.UART_RBAUD[7] ),
    .B(_08648_),
    .X(_08649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15177_ (.A(\design_top.uart0.UART_RBAUD[8] ),
    .B(_08649_),
    .X(_08650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15178_ (.A(\design_top.uart0.UART_RBAUD[9] ),
    .B(_08650_),
    .X(_08651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15179_ (.A(_08651_),
    .Y(_08652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _15180_ (.A(\design_top.uart0.UART_RBAUD[9] ),
    .B(_08650_),
    .X(_08653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15181_ (.A(_08643_),
    .X(_08654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _15182_ (.A1(_08652_),
    .A2(_08653_),
    .B1(_08654_),
    .X(_05732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _15183_ (.A1(\design_top.uart0.UART_RBAUD[7] ),
    .A2(_08648_),
    .B1_N(_08649_),
    .Y(_08655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15184_ (.A(\design_top.uart0.UART_RBAUD[10] ),
    .B(_08651_),
    .X(_08656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15185_ (.A(\design_top.uart0.UART_RBAUD[11] ),
    .B(_08656_),
    .X(_08657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15186_ (.A(\design_top.uart0.UART_RBAUD[12] ),
    .B(_08657_),
    .X(_08658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15187_ (.A(\design_top.uart0.UART_RBAUD[13] ),
    .B(_08658_),
    .X(_08659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _15188_ (.A(\design_top.uart0.UART_RBAUD[14] ),
    .B(_08659_),
    .C(\design_top.uart0.UART_RBAUD[15] ),
    .X(_01949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15189_ (.A(_01949_),
    .Y(_08660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15190_ (.A1(_08655_),
    .A2(_08660_),
    .B1(_08654_),
    .Y(_05731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15191_ (.A(_08648_),
    .Y(_08661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _15192_ (.A(\design_top.uart0.UART_RBAUD[6] ),
    .B(_08647_),
    .X(_08662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _15193_ (.A1(_08661_),
    .A2(_08662_),
    .B1(_08654_),
    .X(_05730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _15194_ (.A1(\design_top.uart0.UART_RBAUD[4] ),
    .A2(_08645_),
    .B1_N(_08646_),
    .Y(_08663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15195_ (.A1(_08660_),
    .A2(_08663_),
    .B1(_08654_),
    .Y(_05729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _15196_ (.A1_N(\design_top.uart0.UART_RBAUD[2] ),
    .A2_N(_08644_),
    .B1(\design_top.uart0.UART_RBAUD[2] ),
    .B2(_08644_),
    .Y(_08664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15197_ (.A(_02662_),
    .B(_08664_),
    .Y(_05728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _15198_ (.A1(\design_top.uart0.UART_RBAUD[1] ),
    .A2(\design_top.uart0.UART_RBAUD[0] ),
    .B1_N(_08644_),
    .Y(_08665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15199_ (.A1(_08660_),
    .A2(_08665_),
    .B1(_08654_),
    .Y(_05727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15200_ (.A(\design_top.core0.RESMODE[2] ),
    .Y(_08666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15201_ (.A(\design_top.core0.RESMODE[0] ),
    .B(\design_top.core0.RESMODE[1] ),
    .Y(_00934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15202_ (.A(_08666_),
    .B(_00934_),
    .Y(_08667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _15203_ (.A1(\design_top.core0.RESMODE[3] ),
    .A2(_08667_),
    .B1(_08348_),
    .X(_05726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15204_ (.A1(_08666_),
    .A2(_00934_),
    .B1(_10872_),
    .Y(_08668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _15205_ (.A1(_08666_),
    .A2(_00934_),
    .A3(\design_top.core0.RESMODE[3] ),
    .B1(_08668_),
    .X(_05725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15206_ (.A(_08348_),
    .B(_00078_),
    .X(_05724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15207_ (.A(\design_top.core0.RESMODE[0] ),
    .Y(_08669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15208_ (.A(\design_top.core0.RESMODE[2] ),
    .B(\design_top.core0.RESMODE[3] ),
    .X(_08670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15209_ (.A(_08670_),
    .X(_03196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _15210_ (.A(\design_top.core0.RESMODE[0] ),
    .B(\design_top.core0.RESMODE[1] ),
    .C(_03196_),
    .X(_00046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _15211_ (.A1(_08669_),
    .A2(_00046_),
    .B1(_08348_),
    .X(_05723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15212_ (.A(_10872_),
    .X(_08671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15213_ (.A(\design_top.IRES[0] ),
    .B(\design_top.IRES[1] ),
    .X(_08672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _15214_ (.A(\design_top.IRES[2] ),
    .B(_08672_),
    .C(\design_top.IRES[3] ),
    .X(_08673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15215_ (.A(\design_top.IRES[4] ),
    .B(_08673_),
    .X(_08674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15216_ (.A(\design_top.IRES[5] ),
    .B(_08674_),
    .X(_08675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15217_ (.A(\design_top.IRES[6] ),
    .B(_08675_),
    .Y(_08676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15218_ (.A(_10795_),
    .X(_08677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15219_ (.A1(_08671_),
    .A2(_08676_),
    .B1(_08677_),
    .Y(_05722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _15220_ (.A1(\design_top.IRES[6] ),
    .A2(_08675_),
    .B1(_08676_),
    .Y(_08678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15221_ (.A1(_08671_),
    .A2(_08678_),
    .B1(_08677_),
    .Y(_05721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _15222_ (.A1(\design_top.IRES[5] ),
    .A2(_08674_),
    .B1_N(_08675_),
    .Y(_08679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15223_ (.A1(_08671_),
    .A2(_08679_),
    .B1(_08677_),
    .Y(_05720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _15224_ (.A1(\design_top.IRES[4] ),
    .A2(_08673_),
    .B1_N(_08674_),
    .Y(_08680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15225_ (.A1(_08671_),
    .A2(_08680_),
    .B1(_08677_),
    .Y(_05719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _15226_ (.A1(\design_top.IRES[2] ),
    .A2(_08672_),
    .B1(\design_top.IRES[3] ),
    .X(_08681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2b_2 _15227_ (.A_N(_08681_),
    .B(_08673_),
    .X(_08682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15228_ (.A1(_08671_),
    .A2(_08682_),
    .B1(_08677_),
    .Y(_05718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _15229_ (.A1_N(\design_top.IRES[2] ),
    .A2_N(_08672_),
    .B1(\design_top.IRES[2] ),
    .B2(_08672_),
    .Y(_08683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15230_ (.A1(_10833_),
    .A2(_08683_),
    .B1(_10795_),
    .Y(_05717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _15231_ (.A1(\design_top.IRES[0] ),
    .A2(\design_top.IRES[1] ),
    .B1_N(_08672_),
    .Y(_08684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15232_ (.A1(_10833_),
    .A2(_08684_),
    .B1(_10795_),
    .Y(_05716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15233_ (.A1(_10833_),
    .A2(\design_top.IRES[0] ),
    .B1(_10795_),
    .Y(_05715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15234_ (.A(_02662_),
    .B(_08660_),
    .X(_08685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15235_ (.A(_08685_),
    .Y(_08686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _15236_ (.A1(\design_top.uart0.UART_RBAUD[14] ),
    .A2(_08659_),
    .B1(\design_top.uart0.UART_RBAUD[15] ),
    .C1(_08686_),
    .X(_05714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15237_ (.A(_08685_),
    .X(_08687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _15238_ (.A1_N(\design_top.uart0.UART_RBAUD[14] ),
    .A2_N(_08659_),
    .B1(\design_top.uart0.UART_RBAUD[14] ),
    .B2(_08659_),
    .Y(_08688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15239_ (.A(_08687_),
    .B(_08688_),
    .Y(_05713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15240_ (.A(\design_top.uart0.UART_RBAUD[13] ),
    .B(_08658_),
    .Y(_08689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _15241_ (.A1(_08659_),
    .A2(_08689_),
    .B1(_08687_),
    .Y(_05712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15242_ (.A(\design_top.uart0.UART_RBAUD[12] ),
    .B(_08657_),
    .Y(_08690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _15243_ (.A1(_08658_),
    .A2(_08690_),
    .B1(_08687_),
    .Y(_05711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15244_ (.A(\design_top.uart0.UART_RBAUD[11] ),
    .B(_08656_),
    .Y(_08691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _15245_ (.A1(_08657_),
    .A2(_08691_),
    .B1(_08687_),
    .Y(_05710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15246_ (.A(\design_top.uart0.UART_RBAUD[10] ),
    .B(_08651_),
    .Y(_08692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _15247_ (.A1(_08656_),
    .A2(_08692_),
    .B1(_08685_),
    .Y(_05709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15248_ (.A(_08650_),
    .Y(_08693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _15249_ (.A1(\design_top.uart0.UART_RBAUD[8] ),
    .A2(_08649_),
    .B1(_08693_),
    .C1(_08685_),
    .X(_05708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15250_ (.A(_08647_),
    .Y(_08694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _15251_ (.A1(\design_top.uart0.UART_RBAUD[5] ),
    .A2(_08646_),
    .B1(_08694_),
    .C1(_08685_),
    .X(_05707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15252_ (.A(_08645_),
    .Y(_08695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _15253_ (.A1(\design_top.uart0.UART_RBAUD[2] ),
    .A2(_08644_),
    .B1(\design_top.uart0.UART_RBAUD[3] ),
    .X(_08696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _15254_ (.A1(_08695_),
    .A2(_08696_),
    .B1(_08686_),
    .X(_05706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15255_ (.A(\design_top.uart0.UART_RBAUD[0] ),
    .B(_08687_),
    .Y(_05705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _15256_ (.A(\design_top.uart0.UART_XBAUD[1] ),
    .B(\design_top.uart0.UART_XBAUD[0] ),
    .C(\design_top.uart0.UART_XBAUD[2] ),
    .D(\design_top.uart0.UART_XBAUD[3] ),
    .X(_08697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15257_ (.A(\design_top.uart0.UART_XBAUD[4] ),
    .B(_08697_),
    .X(_08698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15258_ (.A(\design_top.uart0.UART_XBAUD[5] ),
    .B(_08698_),
    .X(_08699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15259_ (.A(\design_top.uart0.UART_XBAUD[6] ),
    .B(_08699_),
    .X(_08700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15260_ (.A(\design_top.uart0.UART_XBAUD[7] ),
    .B(_08700_),
    .X(_08701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15261_ (.A(\design_top.uart0.UART_XBAUD[8] ),
    .B(_08701_),
    .X(_08702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15262_ (.A(\design_top.uart0.UART_XBAUD[9] ),
    .B(_08702_),
    .X(_08703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15263_ (.A(\design_top.uart0.UART_XBAUD[10] ),
    .B(_08703_),
    .X(_08704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15264_ (.A(\design_top.uart0.UART_XBAUD[11] ),
    .B(_08704_),
    .X(_08705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15265_ (.A(\design_top.uart0.UART_XBAUD[12] ),
    .B(_08705_),
    .X(_08706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15266_ (.A(\design_top.uart0.UART_XBAUD[13] ),
    .B(_08706_),
    .X(_08707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and4_2 _15267_ (.A(\design_top.uart0.UART_XSTATE[1] ),
    .B(_08615_),
    .C(\design_top.uart0.UART_XSTATE[2] ),
    .D(_08612_),
    .X(_02663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _15268_ (.A(\design_top.uart0.UART_XBAUD[14] ),
    .B(_08707_),
    .C(\design_top.uart0.UART_XBAUD[15] ),
    .X(_02623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2b_2 _15269_ (.A(_02663_),
    .B_N(_02623_),
    .X(_08708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15270_ (.A(_08708_),
    .Y(_08709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _15271_ (.A1(\design_top.uart0.UART_XBAUD[14] ),
    .A2(_08707_),
    .B1(\design_top.uart0.UART_XBAUD[15] ),
    .C1(_08709_),
    .X(_05704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15272_ (.A(_08708_),
    .X(_08710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15273_ (.A(_08710_),
    .X(_08711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _15274_ (.A1_N(\design_top.uart0.UART_XBAUD[14] ),
    .A2_N(_08707_),
    .B1(\design_top.uart0.UART_XBAUD[14] ),
    .B2(_08707_),
    .Y(_08712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15275_ (.A(_08711_),
    .B(_08712_),
    .Y(_05703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15276_ (.A(\design_top.uart0.UART_XBAUD[13] ),
    .B(_08706_),
    .Y(_08713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _15277_ (.A1(_08707_),
    .A2(_08713_),
    .B1(_08711_),
    .Y(_05702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15278_ (.A(\design_top.uart0.UART_XBAUD[12] ),
    .B(_08705_),
    .Y(_08714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _15279_ (.A1(_08706_),
    .A2(_08714_),
    .B1(_08711_),
    .Y(_05701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15280_ (.A(\design_top.uart0.UART_XBAUD[11] ),
    .B(_08704_),
    .Y(_08715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15281_ (.A(_08710_),
    .X(_08716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _15282_ (.A1(_08705_),
    .A2(_08715_),
    .B1(_08716_),
    .Y(_05700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15283_ (.A(\design_top.uart0.UART_XBAUD[10] ),
    .B(_08703_),
    .Y(_08717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _15284_ (.A1(_08704_),
    .A2(_08717_),
    .B1(_08716_),
    .Y(_05699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15285_ (.A(_08703_),
    .Y(_08718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _15286_ (.A1(\design_top.uart0.UART_XBAUD[9] ),
    .A2(_08702_),
    .B1(_08718_),
    .C1(_08716_),
    .X(_05698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15287_ (.A(_08702_),
    .Y(_08719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _15288_ (.A1(\design_top.uart0.UART_XBAUD[8] ),
    .A2(_08701_),
    .B1(_08719_),
    .C1(_08710_),
    .X(_05697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15289_ (.A(\design_top.uart0.UART_XBAUD[7] ),
    .B(_08700_),
    .Y(_08720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _15290_ (.A1(_08701_),
    .A2(_08720_),
    .B1(_08716_),
    .Y(_05696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15291_ (.A(_08700_),
    .Y(_08721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _15292_ (.A1(\design_top.uart0.UART_XBAUD[6] ),
    .A2(_08699_),
    .B1(_08721_),
    .C1(_08710_),
    .X(_05695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15293_ (.A(_08699_),
    .Y(_08722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _15294_ (.A1(\design_top.uart0.UART_XBAUD[5] ),
    .A2(_08698_),
    .B1(_08722_),
    .C1(_08710_),
    .X(_05694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _15295_ (.A(\design_top.uart0.UART_XBAUD[4] ),
    .B(_08697_),
    .Y(_08723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _15296_ (.A1(_08698_),
    .A2(_08723_),
    .B1(_08716_),
    .Y(_05693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15297_ (.A(_08697_),
    .Y(_08724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15298_ (.A(\design_top.uart0.UART_XBAUD[1] ),
    .X(_08725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15299_ (.A(\design_top.uart0.UART_XBAUD[0] ),
    .X(_08726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _15300_ (.A1(_08725_),
    .A2(_08726_),
    .A3(\design_top.uart0.UART_XBAUD[2] ),
    .B1(\design_top.uart0.UART_XBAUD[3] ),
    .X(_08727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _15301_ (.A1(_08724_),
    .A2(_08727_),
    .B1(_08709_),
    .X(_05692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _15302_ (.A1(_08725_),
    .A2(\design_top.uart0.UART_XBAUD[0] ),
    .B1(\design_top.uart0.UART_XBAUD[2] ),
    .Y(_08728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o311a_2 _15303_ (.A1(_08725_),
    .A2(_08726_),
    .A3(\design_top.uart0.UART_XBAUD[2] ),
    .B1(_08728_),
    .C1(_08709_),
    .X(_08729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15304_ (.A(_08729_),
    .Y(_05691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _15305_ (.A1_N(_08725_),
    .A2_N(_08726_),
    .B1(_08725_),
    .B2(_08726_),
    .Y(_08730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15306_ (.A(_08711_),
    .B(_08730_),
    .Y(_05690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15307_ (.A(_08726_),
    .B(_08711_),
    .Y(_05689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15308_ (.A(\design_top.IRES[7] ),
    .B(_10844_),
    .X(_08731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15309_ (.A(_08731_),
    .X(_08732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15310_ (.A(_08732_),
    .X(_08733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15311_ (.A(_08733_),
    .X(_08734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15312_ (.A(_08731_),
    .Y(_08735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15313_ (.A(_08735_),
    .X(_08736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15314_ (.A1(\design_top.TIMER[31] ),
    .A2(_08734_),
    .B1(_00037_),
    .B2(_08736_),
    .X(_05688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15315_ (.A1(\design_top.TIMER[30] ),
    .A2(_08734_),
    .B1(_00036_),
    .B2(_08736_),
    .X(_05687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15316_ (.A1(\design_top.TIMER[29] ),
    .A2(_08734_),
    .B1(_00034_),
    .B2(_08736_),
    .X(_05686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15317_ (.A1(\design_top.TIMER[28] ),
    .A2(_08734_),
    .B1(_00033_),
    .B2(_08736_),
    .X(_05685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15318_ (.A(_08735_),
    .X(_08737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15319_ (.A(_08737_),
    .X(_08738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15320_ (.A1(\design_top.TIMER[27] ),
    .A2(_08734_),
    .B1(_00032_),
    .B2(_08738_),
    .X(_05684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15321_ (.A(_08733_),
    .X(_08739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15322_ (.A1(\design_top.TIMER[26] ),
    .A2(_08739_),
    .B1(_00031_),
    .B2(_08738_),
    .X(_05683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15323_ (.A1(\design_top.TIMER[25] ),
    .A2(_08739_),
    .B1(_00030_),
    .B2(_08738_),
    .X(_05682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15324_ (.A1(\design_top.TIMER[24] ),
    .A2(_08739_),
    .B1(_00029_),
    .B2(_08738_),
    .X(_05681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15325_ (.A1(\design_top.TIMER[23] ),
    .A2(_08739_),
    .B1(_00028_),
    .B2(_08738_),
    .X(_05680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15326_ (.A(_08737_),
    .X(_08740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15327_ (.A1(\design_top.TIMER[22] ),
    .A2(_08739_),
    .B1(_00027_),
    .B2(_08740_),
    .X(_05679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15328_ (.A(_08732_),
    .X(_08741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15329_ (.A1(\design_top.TIMER[21] ),
    .A2(_08741_),
    .B1(_00026_),
    .B2(_08740_),
    .X(_05678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15330_ (.A1(\design_top.TIMER[20] ),
    .A2(_08741_),
    .B1(_00025_),
    .B2(_08740_),
    .X(_05677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15331_ (.A1(\design_top.TIMER[19] ),
    .A2(_08741_),
    .B1(_00023_),
    .B2(_08740_),
    .X(_05676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15332_ (.A1(\design_top.TIMER[18] ),
    .A2(_08741_),
    .B1(_00022_),
    .B2(_08740_),
    .X(_05675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15333_ (.A(_08735_),
    .X(_08742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15334_ (.A1(\design_top.TIMER[17] ),
    .A2(_08741_),
    .B1(_00021_),
    .B2(_08742_),
    .X(_05674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15335_ (.A(_08732_),
    .X(_08743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15336_ (.A1(\design_top.TIMER[16] ),
    .A2(_08743_),
    .B1(_00020_),
    .B2(_08742_),
    .X(_05673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15337_ (.A1(\design_top.TIMER[15] ),
    .A2(_08743_),
    .B1(_00019_),
    .B2(_08742_),
    .X(_05672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15338_ (.A1(\design_top.TIMER[14] ),
    .A2(_08743_),
    .B1(_00018_),
    .B2(_08742_),
    .X(_05671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15339_ (.A1(\design_top.TIMER[13] ),
    .A2(_08743_),
    .B1(_00017_),
    .B2(_08742_),
    .X(_05670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15340_ (.A(_08735_),
    .X(_08744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15341_ (.A1(\design_top.TIMER[12] ),
    .A2(_08743_),
    .B1(_00016_),
    .B2(_08744_),
    .X(_05669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15342_ (.A(_08732_),
    .X(_08745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15343_ (.A1(\design_top.TIMER[11] ),
    .A2(_08745_),
    .B1(_00015_),
    .B2(_08744_),
    .X(_05668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15344_ (.A1(\design_top.TIMER[10] ),
    .A2(_08745_),
    .B1(_00014_),
    .B2(_08744_),
    .X(_05667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15345_ (.A1(\design_top.TIMER[9] ),
    .A2(_08745_),
    .B1(_00044_),
    .B2(_08744_),
    .X(_05666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15346_ (.A1(\design_top.TIMER[8] ),
    .A2(_08745_),
    .B1(_00043_),
    .B2(_08744_),
    .X(_05665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15347_ (.A(_08735_),
    .X(_08746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15348_ (.A1(\design_top.TIMER[7] ),
    .A2(_08745_),
    .B1(_00042_),
    .B2(_08746_),
    .X(_05664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15349_ (.A(_08732_),
    .X(_08747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15350_ (.A1(\design_top.TIMER[6] ),
    .A2(_08747_),
    .B1(_00041_),
    .B2(_08746_),
    .X(_05663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15351_ (.A1(\design_top.TIMER[5] ),
    .A2(_08747_),
    .B1(_00040_),
    .B2(_08746_),
    .X(_05662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15352_ (.A1(\design_top.TIMER[4] ),
    .A2(_08747_),
    .B1(_00039_),
    .B2(_08746_),
    .X(_05661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15353_ (.A1(\design_top.TIMER[3] ),
    .A2(_08747_),
    .B1(_00038_),
    .B2(_08746_),
    .X(_05660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15354_ (.A1(\design_top.TIMER[2] ),
    .A2(_08747_),
    .B1(_00035_),
    .B2(_08737_),
    .X(_05659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15355_ (.A1(\design_top.TIMER[1] ),
    .A2(_08733_),
    .B1(_00024_),
    .B2(_08737_),
    .X(_05658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15356_ (.A1(\design_top.TIMER[0] ),
    .A2(_08733_),
    .B1(_00013_),
    .B2(_08737_),
    .X(_05657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15357_ (.A(_10868_),
    .Y(_03197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15358_ (.A(io_out[14]),
    .Y(_08748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _15359_ (.A1(_10868_),
    .A2(_08733_),
    .B1(io_out[14]),
    .X(_08749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _15360_ (.A1(_03197_),
    .A2(_08736_),
    .A3(_08748_),
    .B1(_08749_),
    .X(_05656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15361_ (.A(_03201_),
    .B(_10766_),
    .X(_08750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15362_ (.A(_08750_),
    .X(_08751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15363_ (.A1(_08137_),
    .A2(_10897_),
    .B1(_10886_),
    .B2(_08751_),
    .X(_08752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15364_ (.A(_08752_),
    .Y(_08753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15365_ (.A(_08753_),
    .X(_08754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15366_ (.A(_08752_),
    .X(_08755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15367_ (.A1(_00332_),
    .A2(_08754_),
    .B1(\design_top.MEM[27][7] ),
    .B2(_08755_),
    .X(_05655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15368_ (.A1(_00331_),
    .A2(_08754_),
    .B1(\design_top.MEM[27][6] ),
    .B2(_08755_),
    .X(_05654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15369_ (.A1(_00330_),
    .A2(_08754_),
    .B1(\design_top.MEM[27][5] ),
    .B2(_08755_),
    .X(_05653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15370_ (.A1(_00329_),
    .A2(_08754_),
    .B1(\design_top.MEM[27][4] ),
    .B2(_08755_),
    .X(_05652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15371_ (.A1(_00328_),
    .A2(_08754_),
    .B1(\design_top.MEM[27][3] ),
    .B2(_08755_),
    .X(_05651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15372_ (.A1(_00327_),
    .A2(_08753_),
    .B1(\design_top.MEM[27][2] ),
    .B2(_08752_),
    .X(_05650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15373_ (.A1(_00326_),
    .A2(_08753_),
    .B1(\design_top.MEM[27][1] ),
    .B2(_08752_),
    .X(_05649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15374_ (.A1(_00325_),
    .A2(_08753_),
    .B1(\design_top.MEM[27][0] ),
    .B2(_08752_),
    .X(_05648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15375_ (.A(_08750_),
    .X(_08756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15376_ (.A(_08756_),
    .X(_08757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15377_ (.A1(_08056_),
    .A2(_10965_),
    .B1(_10959_),
    .B2(_08757_),
    .X(_08758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15378_ (.A(_08758_),
    .Y(_08759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15379_ (.A(_08759_),
    .X(_08760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15380_ (.A(_08758_),
    .X(_08761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15381_ (.A1(_00340_),
    .A2(_08760_),
    .B1(\design_top.MEM[28][7] ),
    .B2(_08761_),
    .X(_05647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15382_ (.A1(_00339_),
    .A2(_08760_),
    .B1(\design_top.MEM[28][6] ),
    .B2(_08761_),
    .X(_05646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15383_ (.A1(_00338_),
    .A2(_08760_),
    .B1(\design_top.MEM[28][5] ),
    .B2(_08761_),
    .X(_05645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15384_ (.A1(_00337_),
    .A2(_08760_),
    .B1(\design_top.MEM[28][4] ),
    .B2(_08761_),
    .X(_05644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15385_ (.A1(_00336_),
    .A2(_08760_),
    .B1(\design_top.MEM[28][3] ),
    .B2(_08761_),
    .X(_05643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15386_ (.A1(_00335_),
    .A2(_08759_),
    .B1(\design_top.MEM[28][2] ),
    .B2(_08758_),
    .X(_05642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15387_ (.A1(_00334_),
    .A2(_08759_),
    .B1(\design_top.MEM[28][1] ),
    .B2(_08758_),
    .X(_05641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15388_ (.A1(_00333_),
    .A2(_08759_),
    .B1(\design_top.MEM[28][0] ),
    .B2(_08758_),
    .X(_05640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15389_ (.A1(_10966_),
    .A2(_11195_),
    .B1(_10981_),
    .B2(_08757_),
    .X(_08762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15390_ (.A(_08762_),
    .Y(_08763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15391_ (.A(_08763_),
    .X(_08764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15392_ (.A(_08762_),
    .X(_08765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15393_ (.A1(_00348_),
    .A2(_08764_),
    .B1(\design_top.MEM[29][7] ),
    .B2(_08765_),
    .X(_05639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15394_ (.A1(_00347_),
    .A2(_08764_),
    .B1(\design_top.MEM[29][6] ),
    .B2(_08765_),
    .X(_05638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15395_ (.A1(_00346_),
    .A2(_08764_),
    .B1(\design_top.MEM[29][5] ),
    .B2(_08765_),
    .X(_05637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15396_ (.A1(_00345_),
    .A2(_08764_),
    .B1(\design_top.MEM[29][4] ),
    .B2(_08765_),
    .X(_05636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15397_ (.A1(_00344_),
    .A2(_08764_),
    .B1(\design_top.MEM[29][3] ),
    .B2(_08765_),
    .X(_05635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15398_ (.A1(_00343_),
    .A2(_08763_),
    .B1(\design_top.MEM[29][2] ),
    .B2(_08762_),
    .X(_05634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15399_ (.A1(_00342_),
    .A2(_08763_),
    .B1(\design_top.MEM[29][1] ),
    .B2(_08762_),
    .X(_05633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15400_ (.A1(_00341_),
    .A2(_08763_),
    .B1(\design_top.MEM[29][0] ),
    .B2(_08762_),
    .X(_05632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15401_ (.A1(_10792_),
    .A2(_11134_),
    .B1(_11001_),
    .B2(_08757_),
    .X(_08766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15402_ (.A(_08766_),
    .Y(_08767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15403_ (.A(_08767_),
    .X(_08768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15404_ (.A(_08766_),
    .X(_08769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15405_ (.A1(_00356_),
    .A2(_08768_),
    .B1(\design_top.MEM[2][7] ),
    .B2(_08769_),
    .X(_05631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15406_ (.A1(_00355_),
    .A2(_08768_),
    .B1(\design_top.MEM[2][6] ),
    .B2(_08769_),
    .X(_05630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15407_ (.A1(_00354_),
    .A2(_08768_),
    .B1(\design_top.MEM[2][5] ),
    .B2(_08769_),
    .X(_05629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15408_ (.A1(_00353_),
    .A2(_08768_),
    .B1(\design_top.MEM[2][4] ),
    .B2(_08769_),
    .X(_05628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15409_ (.A1(_00352_),
    .A2(_08768_),
    .B1(\design_top.MEM[2][3] ),
    .B2(_08769_),
    .X(_05627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15410_ (.A1(_00351_),
    .A2(_08767_),
    .B1(\design_top.MEM[2][2] ),
    .B2(_08766_),
    .X(_05626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15411_ (.A1(_00350_),
    .A2(_08767_),
    .B1(\design_top.MEM[2][1] ),
    .B2(_08766_),
    .X(_05625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15412_ (.A1(_00349_),
    .A2(_08767_),
    .B1(\design_top.MEM[2][0] ),
    .B2(_08766_),
    .X(_05624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15413_ (.A1(_10965_),
    .A2(_11134_),
    .B1(_11020_),
    .B2(_08757_),
    .X(_08770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15414_ (.A(_08770_),
    .Y(_08771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15415_ (.A(_08771_),
    .X(_08772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15416_ (.A(_08770_),
    .X(_08773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15417_ (.A1(_00364_),
    .A2(_08772_),
    .B1(\design_top.MEM[30][7] ),
    .B2(_08773_),
    .X(_05623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15418_ (.A1(_00363_),
    .A2(_08772_),
    .B1(\design_top.MEM[30][6] ),
    .B2(_08773_),
    .X(_05622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15419_ (.A1(_00362_),
    .A2(_08772_),
    .B1(\design_top.MEM[30][5] ),
    .B2(_08773_),
    .X(_05621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15420_ (.A1(_00361_),
    .A2(_08772_),
    .B1(\design_top.MEM[30][4] ),
    .B2(_08773_),
    .X(_05620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15421_ (.A1(_00360_),
    .A2(_08772_),
    .B1(\design_top.MEM[30][3] ),
    .B2(_08773_),
    .X(_05619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15422_ (.A1(_00359_),
    .A2(_08771_),
    .B1(\design_top.MEM[30][2] ),
    .B2(_08770_),
    .X(_05618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15423_ (.A1(_00358_),
    .A2(_08771_),
    .B1(\design_top.MEM[30][1] ),
    .B2(_08770_),
    .X(_05617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15424_ (.A1(_00357_),
    .A2(_08771_),
    .B1(\design_top.MEM[30][0] ),
    .B2(_08770_),
    .X(_05616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15425_ (.A1(_08137_),
    .A2(_10965_),
    .B1(_11041_),
    .B2(_08757_),
    .X(_08774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15426_ (.A(_08774_),
    .Y(_08775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15427_ (.A(_08775_),
    .X(_08776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15428_ (.A(_08774_),
    .X(_08777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15429_ (.A1(_00372_),
    .A2(_08776_),
    .B1(\design_top.MEM[31][7] ),
    .B2(_08777_),
    .X(_05615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15430_ (.A1(_00371_),
    .A2(_08776_),
    .B1(\design_top.MEM[31][6] ),
    .B2(_08777_),
    .X(_05614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15431_ (.A1(_00370_),
    .A2(_08776_),
    .B1(\design_top.MEM[31][5] ),
    .B2(_08777_),
    .X(_05613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15432_ (.A1(_00369_),
    .A2(_08776_),
    .B1(\design_top.MEM[31][4] ),
    .B2(_08777_),
    .X(_05612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15433_ (.A1(_00368_),
    .A2(_08776_),
    .B1(\design_top.MEM[31][3] ),
    .B2(_08777_),
    .X(_05611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15434_ (.A1(_00367_),
    .A2(_08775_),
    .B1(\design_top.MEM[31][2] ),
    .B2(_08774_),
    .X(_05610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15435_ (.A1(_00366_),
    .A2(_08775_),
    .B1(\design_top.MEM[31][1] ),
    .B2(_08774_),
    .X(_05609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15436_ (.A1(_00365_),
    .A2(_08775_),
    .B1(\design_top.MEM[31][0] ),
    .B2(_08774_),
    .X(_05608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15437_ (.A(_00861_),
    .X(_08778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15438_ (.A(_00860_),
    .Y(_08779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15439_ (.A(_08779_),
    .X(_08780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15440_ (.A(_00863_),
    .Y(_08781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15441_ (.A(_08781_),
    .X(_08782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _15442_ (.A(_08778_),
    .B(_08780_),
    .C(_08782_),
    .D(_00862_),
    .X(_08783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _15443_ (.A(\design_top.core0.XJALR ),
    .B(\design_top.core0.XJAL ),
    .C(\design_top.core0.XRCC ),
    .D(\design_top.core0.XMCC ),
    .X(_08784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _15444_ (.A(\design_top.core0.XLCC ),
    .B(\design_top.core0.XAUIPC ),
    .C(\design_top.core0.XLUI ),
    .D(_08784_),
    .X(_08785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _15445_ (.A(_00861_),
    .B(_00860_),
    .C(_00863_),
    .D(_00862_),
    .X(_08786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15446_ (.A(_08786_),
    .Y(_08787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _15447_ (.A1(_02661_),
    .A2(_08785_),
    .B1(_08787_),
    .Y(_08788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _15448_ (.A1(_10594_),
    .A2(_08788_),
    .B1(_08432_),
    .X(_08789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15449_ (.A(_08783_),
    .B(_08789_),
    .X(_08790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15450_ (.A(_08790_),
    .X(_08791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15451_ (.A(_08791_),
    .X(_08792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15452_ (.A(_08790_),
    .Y(_08793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15453_ (.A(_08793_),
    .X(_08794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15454_ (.A(_08794_),
    .X(_08795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _15455_ (.A(\design_top.core0.XRES ),
    .B(_08787_),
    .X(_08796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15456_ (.A(_08796_),
    .X(_08797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15457_ (.A(_08797_),
    .X(_08798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15458_ (.A(_00859_),
    .B(_08798_),
    .Y(_08799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15459_ (.A(_08799_),
    .X(_08800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15460_ (.A1(\design_top.core0.REG1[9][31] ),
    .A2(_08792_),
    .B1(_08795_),
    .B2(_08800_),
    .X(_05607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15461_ (.A(_01827_),
    .B(_08798_),
    .Y(_08801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15462_ (.A(_08801_),
    .X(_08802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15463_ (.A1(\design_top.core0.REG1[9][30] ),
    .A2(_08792_),
    .B1(_08795_),
    .B2(_08802_),
    .X(_05606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15464_ (.A(_01806_),
    .B(_08798_),
    .Y(_08803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15465_ (.A(_08803_),
    .X(_08804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15466_ (.A1(\design_top.core0.REG1[9][29] ),
    .A2(_08792_),
    .B1(_08795_),
    .B2(_08804_),
    .X(_05605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15467_ (.A(_01786_),
    .B(_08798_),
    .Y(_08805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15468_ (.A(_08805_),
    .X(_08806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15469_ (.A1(\design_top.core0.REG1[9][28] ),
    .A2(_08792_),
    .B1(_08795_),
    .B2(_08806_),
    .X(_05604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15470_ (.A(_08791_),
    .X(_08807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15471_ (.A(_01764_),
    .B(_08798_),
    .Y(_08808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15472_ (.A(_08808_),
    .X(_08809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15473_ (.A1(\design_top.core0.REG1[9][27] ),
    .A2(_08807_),
    .B1(_08795_),
    .B2(_08809_),
    .X(_05603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15474_ (.A(_08794_),
    .X(_08810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15475_ (.A(_08797_),
    .X(_08811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15476_ (.A(_01745_),
    .B(_08811_),
    .Y(_08812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15477_ (.A(_08812_),
    .X(_08813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15478_ (.A1(\design_top.core0.REG1[9][26] ),
    .A2(_08807_),
    .B1(_08810_),
    .B2(_08813_),
    .X(_05602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15479_ (.A(_01723_),
    .B(_08811_),
    .Y(_08814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15480_ (.A(_08814_),
    .X(_08815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15481_ (.A1(\design_top.core0.REG1[9][25] ),
    .A2(_08807_),
    .B1(_08810_),
    .B2(_08815_),
    .X(_05601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15482_ (.A(_01703_),
    .B(_08811_),
    .Y(_08816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15483_ (.A(_08816_),
    .X(_08817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15484_ (.A1(\design_top.core0.REG1[9][24] ),
    .A2(_08807_),
    .B1(_08810_),
    .B2(_08817_),
    .X(_05600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15485_ (.A(_01681_),
    .B(_08811_),
    .Y(_08818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15486_ (.A(_08818_),
    .X(_08819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15487_ (.A1(\design_top.core0.REG1[9][23] ),
    .A2(_08807_),
    .B1(_08810_),
    .B2(_08819_),
    .X(_05599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15488_ (.A(_08791_),
    .X(_08820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15489_ (.A(_01663_),
    .B(_08811_),
    .Y(_08821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15490_ (.A(_08821_),
    .X(_08822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15491_ (.A1(\design_top.core0.REG1[9][22] ),
    .A2(_08820_),
    .B1(_08810_),
    .B2(_08822_),
    .X(_05598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15492_ (.A(_08794_),
    .X(_08823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15493_ (.A(_08797_),
    .X(_08824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15494_ (.A(_01641_),
    .B(_08824_),
    .Y(_08825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15495_ (.A(_08825_),
    .X(_08826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15496_ (.A1(\design_top.core0.REG1[9][21] ),
    .A2(_08820_),
    .B1(_08823_),
    .B2(_08826_),
    .X(_05597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15497_ (.A(_01621_),
    .B(_08824_),
    .Y(_08827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15498_ (.A(_08827_),
    .X(_08828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15499_ (.A1(\design_top.core0.REG1[9][20] ),
    .A2(_08820_),
    .B1(_08823_),
    .B2(_08828_),
    .X(_05596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15500_ (.A(_01599_),
    .B(_08824_),
    .Y(_08829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15501_ (.A(_08829_),
    .X(_08830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15502_ (.A1(\design_top.core0.REG1[9][19] ),
    .A2(_08820_),
    .B1(_08823_),
    .B2(_08830_),
    .X(_05595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15503_ (.A(_01580_),
    .B(_08824_),
    .Y(_08831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15504_ (.A(_08831_),
    .X(_08832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15505_ (.A1(\design_top.core0.REG1[9][18] ),
    .A2(_08820_),
    .B1(_08823_),
    .B2(_08832_),
    .X(_05594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15506_ (.A(_08790_),
    .X(_08833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15507_ (.A(_01557_),
    .B(_08824_),
    .Y(_08834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15508_ (.A(_08834_),
    .X(_08835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15509_ (.A1(\design_top.core0.REG1[9][17] ),
    .A2(_08833_),
    .B1(_08823_),
    .B2(_08835_),
    .X(_05593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15510_ (.A(_08793_),
    .X(_08836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15511_ (.A(_08797_),
    .X(_08837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15512_ (.A(_01537_),
    .B(_08837_),
    .Y(_08838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15513_ (.A(_08838_),
    .X(_08839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15514_ (.A1(\design_top.core0.REG1[9][16] ),
    .A2(_08833_),
    .B1(_08836_),
    .B2(_08839_),
    .X(_05592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15515_ (.A(_01515_),
    .B(_08837_),
    .Y(_08840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15516_ (.A(_08840_),
    .X(_08841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15517_ (.A1(\design_top.core0.REG1[9][15] ),
    .A2(_08833_),
    .B1(_08836_),
    .B2(_08841_),
    .X(_05591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15518_ (.A(_01499_),
    .B(_08837_),
    .Y(_08842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15519_ (.A(_08842_),
    .X(_08843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15520_ (.A1(\design_top.core0.REG1[9][14] ),
    .A2(_08833_),
    .B1(_08836_),
    .B2(_08843_),
    .X(_05590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15521_ (.A(_00045_),
    .X(_08844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15522_ (.A1(\design_top.core0.REG1[9][13] ),
    .A2(_08794_),
    .B1(_08844_),
    .B2(_08792_),
    .X(_05589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15523_ (.A(_01450_),
    .B(_08837_),
    .Y(_08845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15524_ (.A(_08845_),
    .X(_08846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15525_ (.A1(\design_top.core0.REG1[9][12] ),
    .A2(_08833_),
    .B1(_08836_),
    .B2(_08846_),
    .X(_05588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15526_ (.A(_08790_),
    .X(_08847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15527_ (.A(_01426_),
    .B(_08837_),
    .Y(_08848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15528_ (.A(_08848_),
    .X(_08849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15529_ (.A1(\design_top.core0.REG1[9][11] ),
    .A2(_08847_),
    .B1(_08836_),
    .B2(_08849_),
    .X(_05587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15530_ (.A(_08793_),
    .X(_08850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15531_ (.A(_08796_),
    .X(_08851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15532_ (.A(_01405_),
    .B(_08851_),
    .Y(_08852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15533_ (.A(_08852_),
    .X(_08853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15534_ (.A1(\design_top.core0.REG1[9][10] ),
    .A2(_08847_),
    .B1(_08850_),
    .B2(_08853_),
    .X(_05586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15535_ (.A(_01381_),
    .B(_08851_),
    .Y(_08854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15536_ (.A(_08854_),
    .X(_08855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15537_ (.A1(\design_top.core0.REG1[9][9] ),
    .A2(_08847_),
    .B1(_08850_),
    .B2(_08855_),
    .X(_05585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15538_ (.A(_01359_),
    .B(_08851_),
    .Y(_08856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15539_ (.A(_08856_),
    .X(_08857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15540_ (.A1(\design_top.core0.REG1[9][8] ),
    .A2(_08847_),
    .B1(_08850_),
    .B2(_08857_),
    .X(_05584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15541_ (.A(_01335_),
    .B(_08851_),
    .Y(_08858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15542_ (.A(_08858_),
    .X(_08859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15543_ (.A1(\design_top.core0.REG1[9][7] ),
    .A2(_08847_),
    .B1(_08850_),
    .B2(_08859_),
    .X(_05583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15544_ (.A(_08790_),
    .X(_08860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15545_ (.A(_01312_),
    .B(_08851_),
    .Y(_08861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15546_ (.A(_08861_),
    .X(_08862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15547_ (.A1(\design_top.core0.REG1[9][6] ),
    .A2(_08860_),
    .B1(_08850_),
    .B2(_08862_),
    .X(_05582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15548_ (.A(_08793_),
    .X(_08863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15549_ (.A(_08796_),
    .X(_08864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15550_ (.A(_01266_),
    .B(_08864_),
    .Y(_08865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15551_ (.A(_08865_),
    .X(_08866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15552_ (.A1(\design_top.core0.REG1[9][5] ),
    .A2(_08860_),
    .B1(_08863_),
    .B2(_08866_),
    .X(_05581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15553_ (.A(_01223_),
    .B(_08864_),
    .Y(_08867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15554_ (.A(_08867_),
    .X(_08868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15555_ (.A1(\design_top.core0.REG1[9][4] ),
    .A2(_08860_),
    .B1(_08863_),
    .B2(_08868_),
    .X(_05580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15556_ (.A(_01179_),
    .B(_08864_),
    .Y(_08869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15557_ (.A(_08869_),
    .X(_08870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15558_ (.A1(\design_top.core0.REG1[9][3] ),
    .A2(_08860_),
    .B1(_08863_),
    .B2(_08870_),
    .X(_05579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15559_ (.A(_01131_),
    .B(_08864_),
    .Y(_08871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15560_ (.A(_08871_),
    .X(_08872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15561_ (.A1(\design_top.core0.REG1[9][2] ),
    .A2(_08860_),
    .B1(_08863_),
    .B2(_08872_),
    .X(_05578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15562_ (.A(_01076_),
    .B(_08864_),
    .Y(_08873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15563_ (.A(_08873_),
    .X(_08874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15564_ (.A1(\design_top.core0.REG1[9][1] ),
    .A2(_08791_),
    .B1(_08863_),
    .B2(_08874_),
    .X(_05577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _15565_ (.A(_01008_),
    .B(_08797_),
    .Y(_08875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15566_ (.A(_08875_),
    .X(_08876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15567_ (.A1(\design_top.core0.REG1[9][0] ),
    .A2(_08791_),
    .B1(_08794_),
    .B2(_08876_),
    .X(_05576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15568_ (.A(_08756_),
    .X(_08877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15569_ (.A1(_10791_),
    .A2(_10798_),
    .B1(_10784_),
    .B2(_08877_),
    .X(_08878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15570_ (.A(_08878_),
    .Y(_08879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15571_ (.A(_08879_),
    .X(_08880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15572_ (.A(_08878_),
    .X(_08881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15573_ (.A1(_00180_),
    .A2(_08880_),
    .B1(\design_top.MEM[0][7] ),
    .B2(_08881_),
    .X(_05575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15574_ (.A1(_00179_),
    .A2(_08880_),
    .B1(\design_top.MEM[0][6] ),
    .B2(_08881_),
    .X(_05574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15575_ (.A1(_00178_),
    .A2(_08880_),
    .B1(\design_top.MEM[0][5] ),
    .B2(_08881_),
    .X(_05573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15576_ (.A1(_00177_),
    .A2(_08880_),
    .B1(\design_top.MEM[0][4] ),
    .B2(_08881_),
    .X(_05572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15577_ (.A1(_00176_),
    .A2(_08880_),
    .B1(\design_top.MEM[0][3] ),
    .B2(_08881_),
    .X(_05571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15578_ (.A1(_00175_),
    .A2(_08879_),
    .B1(\design_top.MEM[0][2] ),
    .B2(_08878_),
    .X(_05570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15579_ (.A1(_00174_),
    .A2(_08879_),
    .B1(\design_top.MEM[0][1] ),
    .B2(_08878_),
    .X(_05569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15580_ (.A1(_00173_),
    .A2(_08879_),
    .B1(\design_top.MEM[0][0] ),
    .B2(_08878_),
    .X(_05568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15581_ (.A1(_11005_),
    .A2(_11138_),
    .B1(_11131_),
    .B2(_08877_),
    .X(_08882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15582_ (.A(_08882_),
    .Y(_08883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15583_ (.A(_08883_),
    .X(_08884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15584_ (.A(_08882_),
    .X(_08885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15585_ (.A1(_00188_),
    .A2(_08884_),
    .B1(\design_top.MEM[10][7] ),
    .B2(_08885_),
    .X(_05567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15586_ (.A1(_00187_),
    .A2(_08884_),
    .B1(\design_top.MEM[10][6] ),
    .B2(_08885_),
    .X(_05566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15587_ (.A1(_00186_),
    .A2(_08884_),
    .B1(\design_top.MEM[10][5] ),
    .B2(_08885_),
    .X(_05565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15588_ (.A1(_00185_),
    .A2(_08884_),
    .B1(\design_top.MEM[10][4] ),
    .B2(_08885_),
    .X(_05564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15589_ (.A1(_00184_),
    .A2(_08884_),
    .B1(\design_top.MEM[10][3] ),
    .B2(_08885_),
    .X(_05563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15590_ (.A1(_00183_),
    .A2(_08883_),
    .B1(\design_top.MEM[10][2] ),
    .B2(_08882_),
    .X(_05562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15591_ (.A1(_00182_),
    .A2(_08883_),
    .B1(\design_top.MEM[10][1] ),
    .B2(_08882_),
    .X(_05561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15592_ (.A1(_00181_),
    .A2(_08883_),
    .B1(\design_top.MEM[10][0] ),
    .B2(_08882_),
    .X(_05560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15593_ (.A1(_08137_),
    .A2(_11137_),
    .B1(_11150_),
    .B2(_08877_),
    .X(_08886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15594_ (.A(_08886_),
    .Y(_08887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15595_ (.A(_08887_),
    .X(_08888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15596_ (.A(_08886_),
    .X(_08889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15597_ (.A1(_00196_),
    .A2(_08888_),
    .B1(\design_top.MEM[11][7] ),
    .B2(_08889_),
    .X(_05559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15598_ (.A1(_00195_),
    .A2(_08888_),
    .B1(\design_top.MEM[11][6] ),
    .B2(_08889_),
    .X(_05558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15599_ (.A1(_00194_),
    .A2(_08888_),
    .B1(\design_top.MEM[11][5] ),
    .B2(_08889_),
    .X(_05557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15600_ (.A1(_00193_),
    .A2(_08888_),
    .B1(\design_top.MEM[11][4] ),
    .B2(_08889_),
    .X(_05556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15601_ (.A1(_00192_),
    .A2(_08888_),
    .B1(\design_top.MEM[11][3] ),
    .B2(_08889_),
    .X(_05555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15602_ (.A1(_00191_),
    .A2(_08887_),
    .B1(\design_top.MEM[11][2] ),
    .B2(_08886_),
    .X(_05554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15603_ (.A1(_00190_),
    .A2(_08887_),
    .B1(\design_top.MEM[11][1] ),
    .B2(_08886_),
    .X(_05553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15604_ (.A1(_00189_),
    .A2(_08887_),
    .B1(\design_top.MEM[11][0] ),
    .B2(_08886_),
    .X(_05552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15605_ (.A1(_08056_),
    .A2(_11170_),
    .B1(_11165_),
    .B2(_08877_),
    .X(_08890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15606_ (.A(_08890_),
    .Y(_08891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15607_ (.A(_08891_),
    .X(_08892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15608_ (.A(_08890_),
    .X(_08893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15609_ (.A1(_00204_),
    .A2(_08892_),
    .B1(\design_top.MEM[12][7] ),
    .B2(_08893_),
    .X(_05551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15610_ (.A1(_00203_),
    .A2(_08892_),
    .B1(\design_top.MEM[12][6] ),
    .B2(_08893_),
    .X(_05550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15611_ (.A1(_00202_),
    .A2(_08892_),
    .B1(\design_top.MEM[12][5] ),
    .B2(_08893_),
    .X(_05549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15612_ (.A1(_00201_),
    .A2(_08892_),
    .B1(\design_top.MEM[12][4] ),
    .B2(_08893_),
    .X(_05548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15613_ (.A1(_00200_),
    .A2(_08892_),
    .B1(\design_top.MEM[12][3] ),
    .B2(_08893_),
    .X(_05547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15614_ (.A1(_00199_),
    .A2(_08891_),
    .B1(\design_top.MEM[12][2] ),
    .B2(_08890_),
    .X(_05546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15615_ (.A1(_00198_),
    .A2(_08891_),
    .B1(\design_top.MEM[12][1] ),
    .B2(_08890_),
    .X(_05545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15616_ (.A1(_00197_),
    .A2(_08891_),
    .B1(\design_top.MEM[12][0] ),
    .B2(_08890_),
    .X(_05544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15617_ (.A1(_10986_),
    .A2(_11169_),
    .B1(_11192_),
    .B2(_08877_),
    .X(_08894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15618_ (.A(_08894_),
    .Y(_08895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15619_ (.A(_08895_),
    .X(_08896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15620_ (.A(_08894_),
    .X(_08897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15621_ (.A1(_00212_),
    .A2(_08896_),
    .B1(\design_top.MEM[13][7] ),
    .B2(_08897_),
    .X(_05543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15622_ (.A1(_00211_),
    .A2(_08896_),
    .B1(\design_top.MEM[13][6] ),
    .B2(_08897_),
    .X(_05542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15623_ (.A1(_00210_),
    .A2(_08896_),
    .B1(\design_top.MEM[13][5] ),
    .B2(_08897_),
    .X(_05541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15624_ (.A1(_00209_),
    .A2(_08896_),
    .B1(\design_top.MEM[13][4] ),
    .B2(_08897_),
    .X(_05540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15625_ (.A1(_00208_),
    .A2(_08896_),
    .B1(\design_top.MEM[13][3] ),
    .B2(_08897_),
    .X(_05539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15626_ (.A1(_00207_),
    .A2(_08895_),
    .B1(\design_top.MEM[13][2] ),
    .B2(_08894_),
    .X(_05538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15627_ (.A1(_00206_),
    .A2(_08895_),
    .B1(\design_top.MEM[13][1] ),
    .B2(_08894_),
    .X(_05537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15628_ (.A1(_00205_),
    .A2(_08895_),
    .B1(\design_top.MEM[13][0] ),
    .B2(_08894_),
    .X(_05536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15629_ (.A(_08750_),
    .X(_08898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15630_ (.A(_08898_),
    .X(_08899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15631_ (.A1(_11005_),
    .A2(_11169_),
    .B1(_11226_),
    .B2(_08899_),
    .X(_08900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15632_ (.A(_08900_),
    .Y(_08901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15633_ (.A(_08901_),
    .X(_08902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15634_ (.A(_08900_),
    .X(_08903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15635_ (.A1(_00220_),
    .A2(_08902_),
    .B1(\design_top.MEM[14][7] ),
    .B2(_08903_),
    .X(_05535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15636_ (.A1(_00219_),
    .A2(_08902_),
    .B1(\design_top.MEM[14][6] ),
    .B2(_08903_),
    .X(_05534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15637_ (.A1(_00218_),
    .A2(_08902_),
    .B1(\design_top.MEM[14][5] ),
    .B2(_08903_),
    .X(_05533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15638_ (.A1(_00217_),
    .A2(_08902_),
    .B1(\design_top.MEM[14][4] ),
    .B2(_08903_),
    .X(_05532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15639_ (.A1(_00216_),
    .A2(_08902_),
    .B1(\design_top.MEM[14][3] ),
    .B2(_08903_),
    .X(_05531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15640_ (.A1(_00215_),
    .A2(_08901_),
    .B1(\design_top.MEM[14][2] ),
    .B2(_08900_),
    .X(_05530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15641_ (.A1(_00214_),
    .A2(_08901_),
    .B1(\design_top.MEM[14][1] ),
    .B2(_08900_),
    .X(_05529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15642_ (.A1(_00213_),
    .A2(_08901_),
    .B1(\design_top.MEM[14][0] ),
    .B2(_08900_),
    .X(_05528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15643_ (.A(_10889_),
    .X(_08904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15644_ (.A1(_08904_),
    .A2(_11169_),
    .B1(_11240_),
    .B2(_08899_),
    .X(_08905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15645_ (.A(_08905_),
    .Y(_08906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15646_ (.A(_08906_),
    .X(_08907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15647_ (.A(_08905_),
    .X(_08908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15648_ (.A1(_00228_),
    .A2(_08907_),
    .B1(\design_top.MEM[15][7] ),
    .B2(_08908_),
    .X(_05527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15649_ (.A1(_00227_),
    .A2(_08907_),
    .B1(\design_top.MEM[15][6] ),
    .B2(_08908_),
    .X(_05526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15650_ (.A1(_00226_),
    .A2(_08907_),
    .B1(\design_top.MEM[15][5] ),
    .B2(_08908_),
    .X(_05525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15651_ (.A1(_00225_),
    .A2(_08907_),
    .B1(\design_top.MEM[15][4] ),
    .B2(_08908_),
    .X(_05524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15652_ (.A1(_00224_),
    .A2(_08907_),
    .B1(\design_top.MEM[15][3] ),
    .B2(_08908_),
    .X(_05523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15653_ (.A1(_00223_),
    .A2(_08906_),
    .B1(\design_top.MEM[15][2] ),
    .B2(_08905_),
    .X(_05522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15654_ (.A1(_00222_),
    .A2(_08906_),
    .B1(\design_top.MEM[15][1] ),
    .B2(_08905_),
    .X(_05521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15655_ (.A1(_00221_),
    .A2(_08906_),
    .B1(\design_top.MEM[15][0] ),
    .B2(_08905_),
    .X(_05520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15656_ (.A1(_08056_),
    .A2(_11261_),
    .B1(_11257_),
    .B2(_08899_),
    .X(_08909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15657_ (.A(_08909_),
    .Y(_08910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15658_ (.A(_08910_),
    .X(_08911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15659_ (.A(_08909_),
    .X(_08912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15660_ (.A1(_00236_),
    .A2(_08911_),
    .B1(\design_top.MEM[16][7] ),
    .B2(_08912_),
    .X(_05519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15661_ (.A1(_00235_),
    .A2(_08911_),
    .B1(\design_top.MEM[16][6] ),
    .B2(_08912_),
    .X(_05518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15662_ (.A1(_00234_),
    .A2(_08911_),
    .B1(\design_top.MEM[16][5] ),
    .B2(_08912_),
    .X(_05517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15663_ (.A1(_00233_),
    .A2(_08911_),
    .B1(\design_top.MEM[16][4] ),
    .B2(_08912_),
    .X(_05516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15664_ (.A1(_00232_),
    .A2(_08911_),
    .B1(\design_top.MEM[16][3] ),
    .B2(_08912_),
    .X(_05515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15665_ (.A1(_00231_),
    .A2(_08910_),
    .B1(\design_top.MEM[16][2] ),
    .B2(_08909_),
    .X(_05514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15666_ (.A1(_00230_),
    .A2(_08910_),
    .B1(\design_top.MEM[16][1] ),
    .B2(_08909_),
    .X(_05513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15667_ (.A1(_00229_),
    .A2(_08910_),
    .B1(\design_top.MEM[16][0] ),
    .B2(_08909_),
    .X(_05512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15668_ (.A1(_10986_),
    .A2(_11260_),
    .B1(_11277_),
    .B2(_08899_),
    .X(_08913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15669_ (.A(_08913_),
    .Y(_08914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15670_ (.A(_08914_),
    .X(_08915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15671_ (.A(_08913_),
    .X(_08916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15672_ (.A1(_00244_),
    .A2(_08915_),
    .B1(\design_top.MEM[17][7] ),
    .B2(_08916_),
    .X(_05511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15673_ (.A1(_00243_),
    .A2(_08915_),
    .B1(\design_top.MEM[17][6] ),
    .B2(_08916_),
    .X(_05510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15674_ (.A1(_00242_),
    .A2(_08915_),
    .B1(\design_top.MEM[17][5] ),
    .B2(_08916_),
    .X(_05509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15675_ (.A1(_00241_),
    .A2(_08915_),
    .B1(\design_top.MEM[17][4] ),
    .B2(_08916_),
    .X(_05508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15676_ (.A1(_00240_),
    .A2(_08915_),
    .B1(\design_top.MEM[17][3] ),
    .B2(_08916_),
    .X(_05507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15677_ (.A1(_00239_),
    .A2(_08914_),
    .B1(\design_top.MEM[17][2] ),
    .B2(_08913_),
    .X(_05506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15678_ (.A1(_00238_),
    .A2(_08914_),
    .B1(\design_top.MEM[17][1] ),
    .B2(_08913_),
    .X(_05505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15679_ (.A1(_00237_),
    .A2(_08914_),
    .B1(\design_top.MEM[17][0] ),
    .B2(_08913_),
    .X(_05504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15680_ (.A(_10797_),
    .X(_08917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15681_ (.A1(_08917_),
    .A2(_11112_),
    .B1(_11106_),
    .B2(_08899_),
    .X(_08918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15682_ (.A(_08918_),
    .Y(_08919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15683_ (.A(_08919_),
    .X(_08920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15684_ (.A(_08918_),
    .X(_08921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15685_ (.A1(_00380_),
    .A2(_08920_),
    .B1(\design_top.MEM[32][7] ),
    .B2(_08921_),
    .X(_05503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15686_ (.A1(_00379_),
    .A2(_08920_),
    .B1(\design_top.MEM[32][6] ),
    .B2(_08921_),
    .X(_05502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15687_ (.A1(_00378_),
    .A2(_08920_),
    .B1(\design_top.MEM[32][5] ),
    .B2(_08921_),
    .X(_05501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15688_ (.A1(_00377_),
    .A2(_08920_),
    .B1(\design_top.MEM[32][4] ),
    .B2(_08921_),
    .X(_05500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15689_ (.A1(_00376_),
    .A2(_08920_),
    .B1(\design_top.MEM[32][3] ),
    .B2(_08921_),
    .X(_05499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15690_ (.A1(_00375_),
    .A2(_08919_),
    .B1(\design_top.MEM[32][2] ),
    .B2(_08918_),
    .X(_05498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15691_ (.A1(_00374_),
    .A2(_08919_),
    .B1(\design_top.MEM[32][1] ),
    .B2(_08918_),
    .X(_05497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15692_ (.A1(_00373_),
    .A2(_08919_),
    .B1(\design_top.MEM[32][0] ),
    .B2(_08918_),
    .X(_05496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15693_ (.A(_08898_),
    .X(_08922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15694_ (.A1(_10986_),
    .A2(_11111_),
    .B1(_11287_),
    .B2(_08922_),
    .X(_08923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15695_ (.A(_08923_),
    .Y(_08924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15696_ (.A(_08924_),
    .X(_08925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15697_ (.A(_08923_),
    .X(_08926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15698_ (.A1(_00388_),
    .A2(_08925_),
    .B1(\design_top.MEM[33][7] ),
    .B2(_08926_),
    .X(_05495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15699_ (.A1(_00387_),
    .A2(_08925_),
    .B1(\design_top.MEM[33][6] ),
    .B2(_08926_),
    .X(_05494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15700_ (.A1(_00386_),
    .A2(_08925_),
    .B1(\design_top.MEM[33][5] ),
    .B2(_08926_),
    .X(_05493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15701_ (.A1(_00385_),
    .A2(_08925_),
    .B1(\design_top.MEM[33][4] ),
    .B2(_08926_),
    .X(_05492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15702_ (.A1(_00384_),
    .A2(_08925_),
    .B1(\design_top.MEM[33][3] ),
    .B2(_08926_),
    .X(_05491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15703_ (.A1(_00383_),
    .A2(_08924_),
    .B1(\design_top.MEM[33][2] ),
    .B2(_08923_),
    .X(_05490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15704_ (.A1(_00382_),
    .A2(_08924_),
    .B1(\design_top.MEM[33][1] ),
    .B2(_08923_),
    .X(_05489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15705_ (.A1(_00381_),
    .A2(_08924_),
    .B1(\design_top.MEM[33][0] ),
    .B2(_08923_),
    .X(_05488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15706_ (.A1(_11005_),
    .A2(_11260_),
    .B1(_11342_),
    .B2(_08922_),
    .X(_08927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15707_ (.A(_08927_),
    .Y(_08928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15708_ (.A(_08928_),
    .X(_08929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15709_ (.A(_08927_),
    .X(_08930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15710_ (.A1(_00252_),
    .A2(_08929_),
    .B1(\design_top.MEM[18][7] ),
    .B2(_08930_),
    .X(_05487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15711_ (.A1(_00251_),
    .A2(_08929_),
    .B1(\design_top.MEM[18][6] ),
    .B2(_08930_),
    .X(_05486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15712_ (.A1(_00250_),
    .A2(_08929_),
    .B1(\design_top.MEM[18][5] ),
    .B2(_08930_),
    .X(_05485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15713_ (.A1(_00249_),
    .A2(_08929_),
    .B1(\design_top.MEM[18][4] ),
    .B2(_08930_),
    .X(_05484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15714_ (.A1(_00248_),
    .A2(_08929_),
    .B1(\design_top.MEM[18][3] ),
    .B2(_08930_),
    .X(_05483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15715_ (.A1(_00247_),
    .A2(_08928_),
    .B1(\design_top.MEM[18][2] ),
    .B2(_08927_),
    .X(_05482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15716_ (.A1(_00246_),
    .A2(_08928_),
    .B1(\design_top.MEM[18][1] ),
    .B2(_08927_),
    .X(_05481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15717_ (.A1(_00245_),
    .A2(_08928_),
    .B1(\design_top.MEM[18][0] ),
    .B2(_08927_),
    .X(_05480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15718_ (.A1(_08904_),
    .A2(_11260_),
    .B1(_11355_),
    .B2(_08922_),
    .X(_08931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15719_ (.A(_08931_),
    .Y(_08932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15720_ (.A(_08932_),
    .X(_08933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15721_ (.A(_08931_),
    .X(_08934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15722_ (.A1(_00260_),
    .A2(_08933_),
    .B1(\design_top.MEM[19][7] ),
    .B2(_08934_),
    .X(_05479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15723_ (.A1(_00259_),
    .A2(_08933_),
    .B1(\design_top.MEM[19][6] ),
    .B2(_08934_),
    .X(_05478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15724_ (.A1(_00258_),
    .A2(_08933_),
    .B1(\design_top.MEM[19][5] ),
    .B2(_08934_),
    .X(_05477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15725_ (.A1(_00257_),
    .A2(_08933_),
    .B1(\design_top.MEM[19][4] ),
    .B2(_08934_),
    .X(_05476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15726_ (.A1(_00256_),
    .A2(_08933_),
    .B1(\design_top.MEM[19][3] ),
    .B2(_08934_),
    .X(_05475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15727_ (.A1(_00255_),
    .A2(_08932_),
    .B1(\design_top.MEM[19][2] ),
    .B2(_08931_),
    .X(_05474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15728_ (.A1(_00254_),
    .A2(_08932_),
    .B1(\design_top.MEM[19][1] ),
    .B2(_08931_),
    .X(_05473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15729_ (.A1(_00253_),
    .A2(_08932_),
    .B1(\design_top.MEM[19][0] ),
    .B2(_08931_),
    .X(_05472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15730_ (.A(_11004_),
    .X(_08935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15731_ (.A1(_08935_),
    .A2(_11111_),
    .B1(_11327_),
    .B2(_08922_),
    .X(_08936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15732_ (.A(_08936_),
    .Y(_08937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15733_ (.A(_08937_),
    .X(_08938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15734_ (.A(_08936_),
    .X(_08939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15735_ (.A1(_00396_),
    .A2(_08938_),
    .B1(\design_top.MEM[34][7] ),
    .B2(_08939_),
    .X(_05471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15736_ (.A1(_00395_),
    .A2(_08938_),
    .B1(\design_top.MEM[34][6] ),
    .B2(_08939_),
    .X(_05470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15737_ (.A1(_00394_),
    .A2(_08938_),
    .B1(\design_top.MEM[34][5] ),
    .B2(_08939_),
    .X(_05469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15738_ (.A1(_00393_),
    .A2(_08938_),
    .B1(\design_top.MEM[34][4] ),
    .B2(_08939_),
    .X(_05468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15739_ (.A1(_00392_),
    .A2(_08938_),
    .B1(\design_top.MEM[34][3] ),
    .B2(_08939_),
    .X(_05467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15740_ (.A1(_00391_),
    .A2(_08937_),
    .B1(\design_top.MEM[34][2] ),
    .B2(_08936_),
    .X(_05466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15741_ (.A1(_00390_),
    .A2(_08937_),
    .B1(\design_top.MEM[34][1] ),
    .B2(_08936_),
    .X(_05465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15742_ (.A1(_00389_),
    .A2(_08937_),
    .B1(\design_top.MEM[34][0] ),
    .B2(_08936_),
    .X(_05464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15743_ (.A(_10985_),
    .X(_08940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15744_ (.A1(_08940_),
    .A2(_07572_),
    .B1(_07643_),
    .B2(_08922_),
    .X(_08941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15745_ (.A(_08941_),
    .Y(_08942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15746_ (.A(_08942_),
    .X(_08943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15747_ (.A(_08941_),
    .X(_08944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15748_ (.A1(_00564_),
    .A2(_08943_),
    .B1(\design_top.MEM[53][7] ),
    .B2(_08944_),
    .X(_05463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15749_ (.A1(_00563_),
    .A2(_08943_),
    .B1(\design_top.MEM[53][6] ),
    .B2(_08944_),
    .X(_05462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15750_ (.A1(_00562_),
    .A2(_08943_),
    .B1(\design_top.MEM[53][5] ),
    .B2(_08944_),
    .X(_05461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15751_ (.A1(_00561_),
    .A2(_08943_),
    .B1(\design_top.MEM[53][4] ),
    .B2(_08944_),
    .X(_05460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15752_ (.A1(_00560_),
    .A2(_08943_),
    .B1(\design_top.MEM[53][3] ),
    .B2(_08944_),
    .X(_05459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15753_ (.A1(_00559_),
    .A2(_08942_),
    .B1(\design_top.MEM[53][2] ),
    .B2(_08941_),
    .X(_05458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15754_ (.A1(_00558_),
    .A2(_08942_),
    .B1(\design_top.MEM[53][1] ),
    .B2(_08941_),
    .X(_05457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15755_ (.A1(_00557_),
    .A2(_08942_),
    .B1(\design_top.MEM[53][0] ),
    .B2(_08941_),
    .X(_05456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15756_ (.A(_08898_),
    .X(_08945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15757_ (.A1(_08904_),
    .A2(_11111_),
    .B1(_07442_),
    .B2(_08945_),
    .X(_08946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15758_ (.A(_08946_),
    .Y(_08947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15759_ (.A(_08947_),
    .X(_08948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15760_ (.A(_08946_),
    .X(_08949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15761_ (.A1(_00404_),
    .A2(_08948_),
    .B1(\design_top.MEM[35][7] ),
    .B2(_08949_),
    .X(_05455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15762_ (.A1(_00403_),
    .A2(_08948_),
    .B1(\design_top.MEM[35][6] ),
    .B2(_08949_),
    .X(_05454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15763_ (.A1(_00402_),
    .A2(_08948_),
    .B1(\design_top.MEM[35][5] ),
    .B2(_08949_),
    .X(_05453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15764_ (.A1(_00401_),
    .A2(_08948_),
    .B1(\design_top.MEM[35][4] ),
    .B2(_08949_),
    .X(_05452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15765_ (.A1(_00400_),
    .A2(_08948_),
    .B1(\design_top.MEM[35][3] ),
    .B2(_08949_),
    .X(_05451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15766_ (.A1(_00399_),
    .A2(_08947_),
    .B1(\design_top.MEM[35][2] ),
    .B2(_08946_),
    .X(_05450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15767_ (.A1(_00398_),
    .A2(_08947_),
    .B1(\design_top.MEM[35][1] ),
    .B2(_08946_),
    .X(_05449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15768_ (.A1(_00397_),
    .A2(_08947_),
    .B1(\design_top.MEM[35][0] ),
    .B2(_08946_),
    .X(_05448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15769_ (.A1(_10791_),
    .A2(_11195_),
    .B1(_07956_),
    .B2(_08945_),
    .X(_08950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15770_ (.A(_08950_),
    .Y(_08951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15771_ (.A(_08951_),
    .X(_08952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15772_ (.A(_08950_),
    .X(_08953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15773_ (.A1(_00268_),
    .A2(_08952_),
    .B1(\design_top.MEM[1][7] ),
    .B2(_08953_),
    .X(_05447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15774_ (.A1(_00267_),
    .A2(_08952_),
    .B1(\design_top.MEM[1][6] ),
    .B2(_08953_),
    .X(_05446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15775_ (.A1(_00266_),
    .A2(_08952_),
    .B1(\design_top.MEM[1][5] ),
    .B2(_08953_),
    .X(_05445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15776_ (.A1(_00265_),
    .A2(_08952_),
    .B1(\design_top.MEM[1][4] ),
    .B2(_08953_),
    .X(_05444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15777_ (.A1(_00264_),
    .A2(_08952_),
    .B1(\design_top.MEM[1][3] ),
    .B2(_08953_),
    .X(_05443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15778_ (.A1(_00263_),
    .A2(_08951_),
    .B1(\design_top.MEM[1][2] ),
    .B2(_08950_),
    .X(_05442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15779_ (.A1(_00262_),
    .A2(_08951_),
    .B1(\design_top.MEM[1][1] ),
    .B2(_08950_),
    .X(_05441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15780_ (.A1(_00261_),
    .A2(_08951_),
    .B1(\design_top.MEM[1][0] ),
    .B2(_08950_),
    .X(_05440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15781_ (.A1(_08917_),
    .A2(_07476_),
    .B1(_07472_),
    .B2(_08945_),
    .X(_08954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15782_ (.A(_08954_),
    .Y(_08955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15783_ (.A(_08955_),
    .X(_08956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15784_ (.A(_08954_),
    .X(_08957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15785_ (.A1(_00276_),
    .A2(_08956_),
    .B1(\design_top.MEM[20][7] ),
    .B2(_08957_),
    .X(_05439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15786_ (.A1(_00275_),
    .A2(_08956_),
    .B1(\design_top.MEM[20][6] ),
    .B2(_08957_),
    .X(_05438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15787_ (.A1(_00274_),
    .A2(_08956_),
    .B1(\design_top.MEM[20][5] ),
    .B2(_08957_),
    .X(_05437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15788_ (.A1(_00273_),
    .A2(_08956_),
    .B1(\design_top.MEM[20][4] ),
    .B2(_08957_),
    .X(_05436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15789_ (.A1(_00272_),
    .A2(_08956_),
    .B1(\design_top.MEM[20][3] ),
    .B2(_08957_),
    .X(_05435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15790_ (.A1(_00271_),
    .A2(_08955_),
    .B1(\design_top.MEM[20][2] ),
    .B2(_08954_),
    .X(_05434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15791_ (.A1(_00270_),
    .A2(_08955_),
    .B1(\design_top.MEM[20][1] ),
    .B2(_08954_),
    .X(_05433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15792_ (.A1(_00269_),
    .A2(_08955_),
    .B1(\design_top.MEM[20][0] ),
    .B2(_08954_),
    .X(_05432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15793_ (.A1(_08940_),
    .A2(_07475_),
    .B1(_07505_),
    .B2(_08945_),
    .X(_08958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15794_ (.A(_08958_),
    .Y(_08959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15795_ (.A(_08959_),
    .X(_08960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15796_ (.A(_08958_),
    .X(_08961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15797_ (.A1(_00284_),
    .A2(_08960_),
    .B1(\design_top.MEM[21][7] ),
    .B2(_08961_),
    .X(_05431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15798_ (.A1(_00283_),
    .A2(_08960_),
    .B1(\design_top.MEM[21][6] ),
    .B2(_08961_),
    .X(_05430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15799_ (.A1(_00282_),
    .A2(_08960_),
    .B1(\design_top.MEM[21][5] ),
    .B2(_08961_),
    .X(_05429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15800_ (.A1(_00281_),
    .A2(_08960_),
    .B1(\design_top.MEM[21][4] ),
    .B2(_08961_),
    .X(_05428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15801_ (.A1(_00280_),
    .A2(_08960_),
    .B1(\design_top.MEM[21][3] ),
    .B2(_08961_),
    .X(_05427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15802_ (.A1(_00279_),
    .A2(_08959_),
    .B1(\design_top.MEM[21][2] ),
    .B2(_08958_),
    .X(_05426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15803_ (.A1(_00278_),
    .A2(_08959_),
    .B1(\design_top.MEM[21][1] ),
    .B2(_08958_),
    .X(_05425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15804_ (.A1(_00277_),
    .A2(_08959_),
    .B1(\design_top.MEM[21][0] ),
    .B2(_08958_),
    .X(_05424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15805_ (.A1(_08917_),
    .A2(_07520_),
    .B1(_07516_),
    .B2(_08945_),
    .X(_08962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15806_ (.A(_08962_),
    .Y(_08963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15807_ (.A(_08963_),
    .X(_08964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15808_ (.A(_08962_),
    .X(_08965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15809_ (.A1(_00412_),
    .A2(_08964_),
    .B1(\design_top.MEM[36][7] ),
    .B2(_08965_),
    .X(_05423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15810_ (.A1(_00411_),
    .A2(_08964_),
    .B1(\design_top.MEM[36][6] ),
    .B2(_08965_),
    .X(_05422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15811_ (.A1(_00410_),
    .A2(_08964_),
    .B1(\design_top.MEM[36][5] ),
    .B2(_08965_),
    .X(_05421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15812_ (.A1(_00409_),
    .A2(_08964_),
    .B1(\design_top.MEM[36][4] ),
    .B2(_08965_),
    .X(_05420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15813_ (.A1(_00408_),
    .A2(_08964_),
    .B1(\design_top.MEM[36][3] ),
    .B2(_08965_),
    .X(_05419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15814_ (.A1(_00407_),
    .A2(_08963_),
    .B1(\design_top.MEM[36][2] ),
    .B2(_08962_),
    .X(_05418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15815_ (.A1(_00406_),
    .A2(_08963_),
    .B1(\design_top.MEM[36][1] ),
    .B2(_08962_),
    .X(_05417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15816_ (.A1(_00405_),
    .A2(_08963_),
    .B1(\design_top.MEM[36][0] ),
    .B2(_08962_),
    .X(_05416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15817_ (.A(_08898_),
    .X(_08966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15818_ (.A1(_08935_),
    .A2(_07475_),
    .B1(_07528_),
    .B2(_08966_),
    .X(_08967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15819_ (.A(_08967_),
    .Y(_08968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15820_ (.A(_08968_),
    .X(_08969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15821_ (.A(_08967_),
    .X(_08970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15822_ (.A1(_00292_),
    .A2(_08969_),
    .B1(\design_top.MEM[22][7] ),
    .B2(_08970_),
    .X(_05415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15823_ (.A1(_00291_),
    .A2(_08969_),
    .B1(\design_top.MEM[22][6] ),
    .B2(_08970_),
    .X(_05414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15824_ (.A1(_00290_),
    .A2(_08969_),
    .B1(\design_top.MEM[22][5] ),
    .B2(_08970_),
    .X(_05413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15825_ (.A1(_00289_),
    .A2(_08969_),
    .B1(\design_top.MEM[22][4] ),
    .B2(_08970_),
    .X(_05412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15826_ (.A1(_00288_),
    .A2(_08969_),
    .B1(\design_top.MEM[22][3] ),
    .B2(_08970_),
    .X(_05411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15827_ (.A1(_00287_),
    .A2(_08968_),
    .B1(\design_top.MEM[22][2] ),
    .B2(_08967_),
    .X(_05410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15828_ (.A1(_00286_),
    .A2(_08968_),
    .B1(\design_top.MEM[22][1] ),
    .B2(_08967_),
    .X(_05409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15829_ (.A1(_00285_),
    .A2(_08968_),
    .B1(\design_top.MEM[22][0] ),
    .B2(_08967_),
    .X(_05408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15830_ (.A1(_08904_),
    .A2(_07563_),
    .B1(_07577_),
    .B2(_08966_),
    .X(_08971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15831_ (.A(_08971_),
    .Y(_08972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15832_ (.A(_08972_),
    .X(_08973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15833_ (.A(_08971_),
    .X(_08974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15834_ (.A1(_00548_),
    .A2(_08973_),
    .B1(\design_top.MEM[51][7] ),
    .B2(_08974_),
    .X(_05407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15835_ (.A1(_00547_),
    .A2(_08973_),
    .B1(\design_top.MEM[51][6] ),
    .B2(_08974_),
    .X(_05406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15836_ (.A1(_00546_),
    .A2(_08973_),
    .B1(\design_top.MEM[51][5] ),
    .B2(_08974_),
    .X(_05405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15837_ (.A1(_00545_),
    .A2(_08973_),
    .B1(\design_top.MEM[51][4] ),
    .B2(_08974_),
    .X(_05404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15838_ (.A1(_00544_),
    .A2(_08973_),
    .B1(\design_top.MEM[51][3] ),
    .B2(_08974_),
    .X(_05403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15839_ (.A1(_00543_),
    .A2(_08972_),
    .B1(\design_top.MEM[51][2] ),
    .B2(_08971_),
    .X(_05402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15840_ (.A1(_00542_),
    .A2(_08972_),
    .B1(\design_top.MEM[51][1] ),
    .B2(_08971_),
    .X(_05401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15841_ (.A1(_00541_),
    .A2(_08972_),
    .B1(\design_top.MEM[51][0] ),
    .B2(_08971_),
    .X(_05400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15842_ (.A1(_08935_),
    .A2(_07571_),
    .B1(_07567_),
    .B2(_08966_),
    .X(_08975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15843_ (.A(_08975_),
    .Y(_08976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15844_ (.A(_08976_),
    .X(_08977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15845_ (.A(_08975_),
    .X(_08978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15846_ (.A1(_00572_),
    .A2(_08977_),
    .B1(\design_top.MEM[54][7] ),
    .B2(_08978_),
    .X(_05399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15847_ (.A1(_00571_),
    .A2(_08977_),
    .B1(\design_top.MEM[54][6] ),
    .B2(_08978_),
    .X(_05398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15848_ (.A1(_00570_),
    .A2(_08977_),
    .B1(\design_top.MEM[54][5] ),
    .B2(_08978_),
    .X(_05397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15849_ (.A1(_00569_),
    .A2(_08977_),
    .B1(\design_top.MEM[54][4] ),
    .B2(_08978_),
    .X(_05396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15850_ (.A1(_00568_),
    .A2(_08977_),
    .B1(\design_top.MEM[54][3] ),
    .B2(_08978_),
    .X(_05395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15851_ (.A1(_00567_),
    .A2(_08976_),
    .B1(\design_top.MEM[54][2] ),
    .B2(_08975_),
    .X(_05394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15852_ (.A1(_00566_),
    .A2(_08976_),
    .B1(\design_top.MEM[54][1] ),
    .B2(_08975_),
    .X(_05393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15853_ (.A1(_00565_),
    .A2(_08976_),
    .B1(\design_top.MEM[54][0] ),
    .B2(_08975_),
    .X(_05392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15854_ (.A1(_08917_),
    .A2(_07571_),
    .B1(_07602_),
    .B2(_08966_),
    .X(_08979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15855_ (.A(_08979_),
    .Y(_08980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15856_ (.A(_08980_),
    .X(_08981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15857_ (.A(_08979_),
    .X(_08982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15858_ (.A1(_00556_),
    .A2(_08981_),
    .B1(\design_top.MEM[52][7] ),
    .B2(_08982_),
    .X(_05391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15859_ (.A1(_00555_),
    .A2(_08981_),
    .B1(\design_top.MEM[52][6] ),
    .B2(_08982_),
    .X(_05390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15860_ (.A1(_00554_),
    .A2(_08981_),
    .B1(\design_top.MEM[52][5] ),
    .B2(_08982_),
    .X(_05389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15861_ (.A1(_00553_),
    .A2(_08981_),
    .B1(\design_top.MEM[52][4] ),
    .B2(_08982_),
    .X(_05388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15862_ (.A1(_00552_),
    .A2(_08981_),
    .B1(\design_top.MEM[52][3] ),
    .B2(_08982_),
    .X(_05387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15863_ (.A1(_00551_),
    .A2(_08980_),
    .B1(\design_top.MEM[52][2] ),
    .B2(_08979_),
    .X(_05386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15864_ (.A1(_00550_),
    .A2(_08980_),
    .B1(\design_top.MEM[52][1] ),
    .B2(_08979_),
    .X(_05385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15865_ (.A1(_00549_),
    .A2(_08980_),
    .B1(\design_top.MEM[52][0] ),
    .B2(_08979_),
    .X(_05384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15866_ (.A1(_08904_),
    .A2(_07519_),
    .B1(_07698_),
    .B2(_08966_),
    .X(_08983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15867_ (.A(_08983_),
    .Y(_08984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15868_ (.A(_08984_),
    .X(_08985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15869_ (.A(_08983_),
    .X(_08986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15870_ (.A1(_00436_),
    .A2(_08985_),
    .B1(\design_top.MEM[39][7] ),
    .B2(_08986_),
    .X(_05383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15871_ (.A1(_00435_),
    .A2(_08985_),
    .B1(\design_top.MEM[39][6] ),
    .B2(_08986_),
    .X(_05382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15872_ (.A1(_00434_),
    .A2(_08985_),
    .B1(\design_top.MEM[39][5] ),
    .B2(_08986_),
    .X(_05381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15873_ (.A1(_00433_),
    .A2(_08985_),
    .B1(\design_top.MEM[39][4] ),
    .B2(_08986_),
    .X(_05380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15874_ (.A1(_00432_),
    .A2(_08985_),
    .B1(\design_top.MEM[39][3] ),
    .B2(_08986_),
    .X(_05379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15875_ (.A1(_00431_),
    .A2(_08984_),
    .B1(\design_top.MEM[39][2] ),
    .B2(_08983_),
    .X(_05378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15876_ (.A1(_00430_),
    .A2(_08984_),
    .B1(\design_top.MEM[39][1] ),
    .B2(_08983_),
    .X(_05377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15877_ (.A1(_00429_),
    .A2(_08984_),
    .B1(\design_top.MEM[39][0] ),
    .B2(_08983_),
    .X(_05376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15878_ (.A(_08898_),
    .X(_08987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15879_ (.A1(_08935_),
    .A2(_07455_),
    .B1(_07703_),
    .B2(_08987_),
    .X(_08988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15880_ (.A(_08988_),
    .Y(_08989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15881_ (.A(_08989_),
    .X(_08990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15882_ (.A(_08988_),
    .X(_08991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15883_ (.A1(_00500_),
    .A2(_08990_),
    .B1(\design_top.MEM[46][7] ),
    .B2(_08991_),
    .X(_05375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15884_ (.A1(_00499_),
    .A2(_08990_),
    .B1(\design_top.MEM[46][6] ),
    .B2(_08991_),
    .X(_05374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15885_ (.A1(_00498_),
    .A2(_08990_),
    .B1(\design_top.MEM[46][5] ),
    .B2(_08991_),
    .X(_05373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15886_ (.A1(_00497_),
    .A2(_08990_),
    .B1(\design_top.MEM[46][4] ),
    .B2(_08991_),
    .X(_05372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15887_ (.A1(_00496_),
    .A2(_08990_),
    .B1(\design_top.MEM[46][3] ),
    .B2(_08991_),
    .X(_05371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15888_ (.A1(_00495_),
    .A2(_08989_),
    .B1(\design_top.MEM[46][2] ),
    .B2(_08988_),
    .X(_05370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15889_ (.A1(_00494_),
    .A2(_08989_),
    .B1(\design_top.MEM[46][1] ),
    .B2(_08988_),
    .X(_05369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15890_ (.A1(_00493_),
    .A2(_08989_),
    .B1(\design_top.MEM[46][0] ),
    .B2(_08988_),
    .X(_05368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15891_ (.A(_10889_),
    .X(_08992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15892_ (.A1(_08992_),
    .A2(_07454_),
    .B1(_07728_),
    .B2(_08987_),
    .X(_08993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15893_ (.A(_08993_),
    .Y(_08994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15894_ (.A(_08994_),
    .X(_08995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15895_ (.A(_08993_),
    .X(_08996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15896_ (.A1(_00508_),
    .A2(_08995_),
    .B1(\design_top.MEM[47][7] ),
    .B2(_08996_),
    .X(_05367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15897_ (.A1(_00507_),
    .A2(_08995_),
    .B1(\design_top.MEM[47][6] ),
    .B2(_08996_),
    .X(_05366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15898_ (.A1(_00506_),
    .A2(_08995_),
    .B1(\design_top.MEM[47][5] ),
    .B2(_08996_),
    .X(_05365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15899_ (.A1(_00505_),
    .A2(_08995_),
    .B1(\design_top.MEM[47][4] ),
    .B2(_08996_),
    .X(_05364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15900_ (.A1(_00504_),
    .A2(_08995_),
    .B1(\design_top.MEM[47][3] ),
    .B2(_08996_),
    .X(_05363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15901_ (.A1(_00503_),
    .A2(_08994_),
    .B1(\design_top.MEM[47][2] ),
    .B2(_08993_),
    .X(_05362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15902_ (.A1(_00502_),
    .A2(_08994_),
    .B1(\design_top.MEM[47][1] ),
    .B2(_08993_),
    .X(_05361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15903_ (.A1(_00501_),
    .A2(_08994_),
    .B1(\design_top.MEM[47][0] ),
    .B2(_08993_),
    .X(_05360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15904_ (.A1(_10791_),
    .A2(_10890_),
    .B1(_07751_),
    .B2(_08987_),
    .X(_08997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15905_ (.A(_08997_),
    .Y(_08998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15906_ (.A(_08998_),
    .X(_08999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15907_ (.A(_08997_),
    .X(_09000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15908_ (.A1(_00444_),
    .A2(_08999_),
    .B1(\design_top.MEM[3][7] ),
    .B2(_09000_),
    .X(_05359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15909_ (.A1(_00443_),
    .A2(_08999_),
    .B1(\design_top.MEM[3][6] ),
    .B2(_09000_),
    .X(_05358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15910_ (.A1(_00442_),
    .A2(_08999_),
    .B1(\design_top.MEM[3][5] ),
    .B2(_09000_),
    .X(_05357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15911_ (.A1(_00441_),
    .A2(_08999_),
    .B1(\design_top.MEM[3][4] ),
    .B2(_09000_),
    .X(_05356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15912_ (.A1(_00440_),
    .A2(_08999_),
    .B1(\design_top.MEM[3][3] ),
    .B2(_09000_),
    .X(_05355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15913_ (.A1(_00439_),
    .A2(_08998_),
    .B1(\design_top.MEM[3][2] ),
    .B2(_08997_),
    .X(_05354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15914_ (.A1(_00438_),
    .A2(_08998_),
    .B1(\design_top.MEM[3][1] ),
    .B2(_08997_),
    .X(_05353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15915_ (.A1(_00437_),
    .A2(_08998_),
    .B1(\design_top.MEM[3][0] ),
    .B2(_08997_),
    .X(_05352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15916_ (.A1(_08917_),
    .A2(_07777_),
    .B1(_07772_),
    .B2(_08987_),
    .X(_09001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15917_ (.A(_09001_),
    .Y(_09002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15918_ (.A(_09002_),
    .X(_09003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15919_ (.A(_09001_),
    .X(_09004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15920_ (.A1(_00452_),
    .A2(_09003_),
    .B1(\design_top.MEM[40][7] ),
    .B2(_09004_),
    .X(_05351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15921_ (.A1(_00451_),
    .A2(_09003_),
    .B1(\design_top.MEM[40][6] ),
    .B2(_09004_),
    .X(_05350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15922_ (.A1(_00450_),
    .A2(_09003_),
    .B1(\design_top.MEM[40][5] ),
    .B2(_09004_),
    .X(_05349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15923_ (.A1(_00449_),
    .A2(_09003_),
    .B1(\design_top.MEM[40][4] ),
    .B2(_09004_),
    .X(_05348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15924_ (.A1(_00448_),
    .A2(_09003_),
    .B1(\design_top.MEM[40][3] ),
    .B2(_09004_),
    .X(_05347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15925_ (.A1(_00447_),
    .A2(_09002_),
    .B1(\design_top.MEM[40][2] ),
    .B2(_09001_),
    .X(_05346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15926_ (.A1(_00446_),
    .A2(_09002_),
    .B1(\design_top.MEM[40][1] ),
    .B2(_09001_),
    .X(_05345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15927_ (.A1(_00445_),
    .A2(_09002_),
    .B1(\design_top.MEM[40][0] ),
    .B2(_09001_),
    .X(_05344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15928_ (.A(_10797_),
    .X(_09005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15929_ (.A1(_09005_),
    .A2(_07562_),
    .B1(_07781_),
    .B2(_08987_),
    .X(_09006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15930_ (.A(_09006_),
    .Y(_09007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15931_ (.A(_09007_),
    .X(_09008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15932_ (.A(_09006_),
    .X(_09009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15933_ (.A1(_00516_),
    .A2(_09008_),
    .B1(\design_top.MEM[48][7] ),
    .B2(_09009_),
    .X(_05343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15934_ (.A1(_00515_),
    .A2(_09008_),
    .B1(\design_top.MEM[48][6] ),
    .B2(_09009_),
    .X(_05342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15935_ (.A1(_00514_),
    .A2(_09008_),
    .B1(\design_top.MEM[48][5] ),
    .B2(_09009_),
    .X(_05341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15936_ (.A1(_00513_),
    .A2(_09008_),
    .B1(\design_top.MEM[48][4] ),
    .B2(_09009_),
    .X(_05340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15937_ (.A1(_00512_),
    .A2(_09008_),
    .B1(\design_top.MEM[48][3] ),
    .B2(_09009_),
    .X(_05339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15938_ (.A1(_00511_),
    .A2(_09007_),
    .B1(\design_top.MEM[48][2] ),
    .B2(_09006_),
    .X(_05338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15939_ (.A1(_00510_),
    .A2(_09007_),
    .B1(\design_top.MEM[48][1] ),
    .B2(_09006_),
    .X(_05337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15940_ (.A1(_00509_),
    .A2(_09007_),
    .B1(\design_top.MEM[48][0] ),
    .B2(_09006_),
    .X(_05336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15941_ (.A(_08750_),
    .X(_09010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15942_ (.A(_09010_),
    .X(_09011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15943_ (.A1(_08940_),
    .A2(_07776_),
    .B1(_07822_),
    .B2(_09011_),
    .X(_09012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15944_ (.A(_09012_),
    .Y(_09013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15945_ (.A(_09013_),
    .X(_09014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15946_ (.A(_09012_),
    .X(_09015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15947_ (.A1(_00460_),
    .A2(_09014_),
    .B1(\design_top.MEM[41][7] ),
    .B2(_09015_),
    .X(_05335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15948_ (.A1(_00459_),
    .A2(_09014_),
    .B1(\design_top.MEM[41][6] ),
    .B2(_09015_),
    .X(_05334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15949_ (.A1(_00458_),
    .A2(_09014_),
    .B1(\design_top.MEM[41][5] ),
    .B2(_09015_),
    .X(_05333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15950_ (.A1(_00457_),
    .A2(_09014_),
    .B1(\design_top.MEM[41][4] ),
    .B2(_09015_),
    .X(_05332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15951_ (.A1(_00456_),
    .A2(_09014_),
    .B1(\design_top.MEM[41][3] ),
    .B2(_09015_),
    .X(_05331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15952_ (.A1(_00455_),
    .A2(_09013_),
    .B1(\design_top.MEM[41][2] ),
    .B2(_09012_),
    .X(_05330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15953_ (.A1(_00454_),
    .A2(_09013_),
    .B1(\design_top.MEM[41][1] ),
    .B2(_09012_),
    .X(_05329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15954_ (.A1(_00453_),
    .A2(_09013_),
    .B1(\design_top.MEM[41][0] ),
    .B2(_09012_),
    .X(_05328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15955_ (.A1(_08940_),
    .A2(_07562_),
    .B1(_07828_),
    .B2(_09011_),
    .X(_09016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15956_ (.A(_09016_),
    .Y(_09017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15957_ (.A(_09017_),
    .X(_09018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15958_ (.A(_09016_),
    .X(_09019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15959_ (.A1(_00524_),
    .A2(_09018_),
    .B1(\design_top.MEM[49][7] ),
    .B2(_09019_),
    .X(_05327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15960_ (.A1(_00523_),
    .A2(_09018_),
    .B1(\design_top.MEM[49][6] ),
    .B2(_09019_),
    .X(_05326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15961_ (.A1(_00522_),
    .A2(_09018_),
    .B1(\design_top.MEM[49][5] ),
    .B2(_09019_),
    .X(_05325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15962_ (.A1(_00521_),
    .A2(_09018_),
    .B1(\design_top.MEM[49][4] ),
    .B2(_09019_),
    .X(_05324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15963_ (.A1(_00520_),
    .A2(_09018_),
    .B1(\design_top.MEM[49][3] ),
    .B2(_09019_),
    .X(_05323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15964_ (.A1(_00519_),
    .A2(_09017_),
    .B1(\design_top.MEM[49][2] ),
    .B2(_09016_),
    .X(_05322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15965_ (.A1(_00518_),
    .A2(_09017_),
    .B1(\design_top.MEM[49][1] ),
    .B2(_09016_),
    .X(_05321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15966_ (.A1(_00517_),
    .A2(_09017_),
    .B1(\design_top.MEM[49][0] ),
    .B2(_09016_),
    .X(_05320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15967_ (.A1(_08935_),
    .A2(_07776_),
    .B1(_07851_),
    .B2(_09011_),
    .X(_09020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15968_ (.A(_09020_),
    .Y(_09021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15969_ (.A(_09021_),
    .X(_09022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15970_ (.A(_09020_),
    .X(_09023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15971_ (.A1(_00468_),
    .A2(_09022_),
    .B1(\design_top.MEM[42][7] ),
    .B2(_09023_),
    .X(_05319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15972_ (.A1(_00467_),
    .A2(_09022_),
    .B1(\design_top.MEM[42][6] ),
    .B2(_09023_),
    .X(_05318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15973_ (.A1(_00466_),
    .A2(_09022_),
    .B1(\design_top.MEM[42][5] ),
    .B2(_09023_),
    .X(_05317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15974_ (.A1(_00465_),
    .A2(_09022_),
    .B1(\design_top.MEM[42][4] ),
    .B2(_09023_),
    .X(_05316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15975_ (.A1(_00464_),
    .A2(_09022_),
    .B1(\design_top.MEM[42][3] ),
    .B2(_09023_),
    .X(_05315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15976_ (.A1(_00463_),
    .A2(_09021_),
    .B1(\design_top.MEM[42][2] ),
    .B2(_09020_),
    .X(_05314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15977_ (.A1(_00462_),
    .A2(_09021_),
    .B1(\design_top.MEM[42][1] ),
    .B2(_09020_),
    .X(_05313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15978_ (.A1(_00461_),
    .A2(_09021_),
    .B1(\design_top.MEM[42][0] ),
    .B2(_09020_),
    .X(_05312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15979_ (.A1(_09005_),
    .A2(_07868_),
    .B1(_07864_),
    .B2(_09011_),
    .X(_09024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15980_ (.A(_09024_),
    .Y(_09025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15981_ (.A(_09025_),
    .X(_09026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15982_ (.A(_09024_),
    .X(_09027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15983_ (.A1(_00532_),
    .A2(_09026_),
    .B1(\design_top.MEM[4][7] ),
    .B2(_09027_),
    .X(_05311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15984_ (.A1(_00531_),
    .A2(_09026_),
    .B1(\design_top.MEM[4][6] ),
    .B2(_09027_),
    .X(_05310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15985_ (.A1(_00530_),
    .A2(_09026_),
    .B1(\design_top.MEM[4][5] ),
    .B2(_09027_),
    .X(_05309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15986_ (.A1(_00529_),
    .A2(_09026_),
    .B1(\design_top.MEM[4][4] ),
    .B2(_09027_),
    .X(_05308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15987_ (.A1(_00528_),
    .A2(_09026_),
    .B1(\design_top.MEM[4][3] ),
    .B2(_09027_),
    .X(_05307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15988_ (.A1(_00527_),
    .A2(_09025_),
    .B1(\design_top.MEM[4][2] ),
    .B2(_09024_),
    .X(_05306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15989_ (.A1(_00526_),
    .A2(_09025_),
    .B1(\design_top.MEM[4][1] ),
    .B2(_09024_),
    .X(_05305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15990_ (.A1(_00525_),
    .A2(_09025_),
    .B1(\design_top.MEM[4][0] ),
    .B2(_09024_),
    .X(_05304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _15991_ (.A1(_08992_),
    .A2(_07776_),
    .B1(_07906_),
    .B2(_09011_),
    .X(_09028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _15992_ (.A(_09028_),
    .Y(_09029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15993_ (.A(_09029_),
    .X(_09030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _15994_ (.A(_09028_),
    .X(_09031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15995_ (.A1(_00476_),
    .A2(_09030_),
    .B1(\design_top.MEM[43][7] ),
    .B2(_09031_),
    .X(_05303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15996_ (.A1(_00475_),
    .A2(_09030_),
    .B1(\design_top.MEM[43][6] ),
    .B2(_09031_),
    .X(_05302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15997_ (.A1(_00474_),
    .A2(_09030_),
    .B1(\design_top.MEM[43][5] ),
    .B2(_09031_),
    .X(_05301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15998_ (.A1(_00473_),
    .A2(_09030_),
    .B1(\design_top.MEM[43][4] ),
    .B2(_09031_),
    .X(_05300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _15999_ (.A1(_00472_),
    .A2(_09030_),
    .B1(\design_top.MEM[43][3] ),
    .B2(_09031_),
    .X(_05299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16000_ (.A1(_00471_),
    .A2(_09029_),
    .B1(\design_top.MEM[43][2] ),
    .B2(_09028_),
    .X(_05298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16001_ (.A1(_00470_),
    .A2(_09029_),
    .B1(\design_top.MEM[43][1] ),
    .B2(_09028_),
    .X(_05297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16002_ (.A1(_00469_),
    .A2(_09029_),
    .B1(\design_top.MEM[43][0] ),
    .B2(_09028_),
    .X(_05296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16003_ (.A(_11004_),
    .X(_09032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16004_ (.A(_09010_),
    .X(_09033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16005_ (.A1(_09032_),
    .A2(_07562_),
    .B1(_07559_),
    .B2(_09033_),
    .X(_09034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16006_ (.A(_09034_),
    .Y(_09035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16007_ (.A(_09035_),
    .X(_09036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16008_ (.A(_09034_),
    .X(_09037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16009_ (.A1(_00540_),
    .A2(_09036_),
    .B1(\design_top.MEM[50][7] ),
    .B2(_09037_),
    .X(_05295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16010_ (.A1(_00539_),
    .A2(_09036_),
    .B1(\design_top.MEM[50][6] ),
    .B2(_09037_),
    .X(_05294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16011_ (.A1(_00538_),
    .A2(_09036_),
    .B1(\design_top.MEM[50][5] ),
    .B2(_09037_),
    .X(_05293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16012_ (.A1(_00537_),
    .A2(_09036_),
    .B1(\design_top.MEM[50][4] ),
    .B2(_09037_),
    .X(_05292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16013_ (.A1(_00536_),
    .A2(_09036_),
    .B1(\design_top.MEM[50][3] ),
    .B2(_09037_),
    .X(_05291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16014_ (.A1(_00535_),
    .A2(_09035_),
    .B1(\design_top.MEM[50][2] ),
    .B2(_09034_),
    .X(_05290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16015_ (.A1(_00534_),
    .A2(_09035_),
    .B1(\design_top.MEM[50][1] ),
    .B2(_09034_),
    .X(_05289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16016_ (.A1(_00533_),
    .A2(_09035_),
    .B1(\design_top.MEM[50][0] ),
    .B2(_09034_),
    .X(_05288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16017_ (.A1(_09005_),
    .A2(_07454_),
    .B1(_07930_),
    .B2(_09033_),
    .X(_09038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16018_ (.A(_09038_),
    .Y(_09039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16019_ (.A(_09039_),
    .X(_09040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16020_ (.A(_09038_),
    .X(_09041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16021_ (.A1(_00484_),
    .A2(_09040_),
    .B1(\design_top.MEM[44][7] ),
    .B2(_09041_),
    .X(_05287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16022_ (.A1(_00483_),
    .A2(_09040_),
    .B1(\design_top.MEM[44][6] ),
    .B2(_09041_),
    .X(_05286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16023_ (.A1(_00482_),
    .A2(_09040_),
    .B1(\design_top.MEM[44][5] ),
    .B2(_09041_),
    .X(_05285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16024_ (.A1(_00481_),
    .A2(_09040_),
    .B1(\design_top.MEM[44][4] ),
    .B2(_09041_),
    .X(_05284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16025_ (.A1(_00480_),
    .A2(_09040_),
    .B1(\design_top.MEM[44][3] ),
    .B2(_09041_),
    .X(_05283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16026_ (.A1(_00479_),
    .A2(_09039_),
    .B1(\design_top.MEM[44][2] ),
    .B2(_09038_),
    .X(_05282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16027_ (.A1(_00478_),
    .A2(_09039_),
    .B1(\design_top.MEM[44][1] ),
    .B2(_09038_),
    .X(_05281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16028_ (.A1(_00477_),
    .A2(_09039_),
    .B1(\design_top.MEM[44][0] ),
    .B2(_09038_),
    .X(_05280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16029_ (.A1(_08940_),
    .A2(_07454_),
    .B1(_07451_),
    .B2(_09033_),
    .X(_09042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16030_ (.A(_09042_),
    .Y(_09043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16031_ (.A(_09043_),
    .X(_09044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16032_ (.A(_09042_),
    .X(_09045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16033_ (.A1(_00492_),
    .A2(_09044_),
    .B1(\design_top.MEM[45][7] ),
    .B2(_09045_),
    .X(_05279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16034_ (.A1(_00491_),
    .A2(_09044_),
    .B1(\design_top.MEM[45][6] ),
    .B2(_09045_),
    .X(_05278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16035_ (.A1(_00490_),
    .A2(_09044_),
    .B1(\design_top.MEM[45][5] ),
    .B2(_09045_),
    .X(_05277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16036_ (.A1(_00489_),
    .A2(_09044_),
    .B1(\design_top.MEM[45][4] ),
    .B2(_09045_),
    .X(_05276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16037_ (.A1(_00488_),
    .A2(_09044_),
    .B1(\design_top.MEM[45][3] ),
    .B2(_09045_),
    .X(_05275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16038_ (.A1(_00487_),
    .A2(_09043_),
    .B1(\design_top.MEM[45][2] ),
    .B2(_09042_),
    .X(_05274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16039_ (.A1(_00486_),
    .A2(_09043_),
    .B1(\design_top.MEM[45][1] ),
    .B2(_09042_),
    .X(_05273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16040_ (.A1(_00485_),
    .A2(_09043_),
    .B1(\design_top.MEM[45][0] ),
    .B2(_09042_),
    .X(_05272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16041_ (.A1(_08992_),
    .A2(_07475_),
    .B1(_07973_),
    .B2(_09033_),
    .X(_09046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16042_ (.A(_09046_),
    .Y(_09047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16043_ (.A(_09047_),
    .X(_09048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16044_ (.A(_09046_),
    .X(_09049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16045_ (.A1(_00300_),
    .A2(_09048_),
    .B1(\design_top.MEM[23][7] ),
    .B2(_09049_),
    .X(_05271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16046_ (.A1(_00299_),
    .A2(_09048_),
    .B1(\design_top.MEM[23][6] ),
    .B2(_09049_),
    .X(_05270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16047_ (.A1(_00298_),
    .A2(_09048_),
    .B1(\design_top.MEM[23][5] ),
    .B2(_09049_),
    .X(_05269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16048_ (.A1(_00297_),
    .A2(_09048_),
    .B1(\design_top.MEM[23][4] ),
    .B2(_09049_),
    .X(_05268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16049_ (.A1(_00296_),
    .A2(_09048_),
    .B1(\design_top.MEM[23][3] ),
    .B2(_09049_),
    .X(_05267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16050_ (.A1(_00295_),
    .A2(_09047_),
    .B1(\design_top.MEM[23][2] ),
    .B2(_09046_),
    .X(_05266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16051_ (.A1(_00294_),
    .A2(_09047_),
    .B1(\design_top.MEM[23][1] ),
    .B2(_09046_),
    .X(_05265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16052_ (.A1(_00293_),
    .A2(_09047_),
    .B1(\design_top.MEM[23][0] ),
    .B2(_09046_),
    .X(_05264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16053_ (.A(_10985_),
    .X(_09050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16054_ (.A1(_09050_),
    .A2(_07519_),
    .B1(_07978_),
    .B2(_09033_),
    .X(_09051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16055_ (.A(_09051_),
    .Y(_09052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16056_ (.A(_09052_),
    .X(_09053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16057_ (.A(_09051_),
    .X(_09054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16058_ (.A1(_00420_),
    .A2(_09053_),
    .B1(\design_top.MEM[37][7] ),
    .B2(_09054_),
    .X(_05263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16059_ (.A1(_00419_),
    .A2(_09053_),
    .B1(\design_top.MEM[37][6] ),
    .B2(_09054_),
    .X(_05262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16060_ (.A1(_00418_),
    .A2(_09053_),
    .B1(\design_top.MEM[37][5] ),
    .B2(_09054_),
    .X(_05261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16061_ (.A1(_00417_),
    .A2(_09053_),
    .B1(\design_top.MEM[37][4] ),
    .B2(_09054_),
    .X(_05260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16062_ (.A1(_00416_),
    .A2(_09053_),
    .B1(\design_top.MEM[37][3] ),
    .B2(_09054_),
    .X(_05259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16063_ (.A1(_00415_),
    .A2(_09052_),
    .B1(\design_top.MEM[37][2] ),
    .B2(_09051_),
    .X(_05258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16064_ (.A1(_00414_),
    .A2(_09052_),
    .B1(\design_top.MEM[37][1] ),
    .B2(_09051_),
    .X(_05257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16065_ (.A1(_00413_),
    .A2(_09052_),
    .B1(\design_top.MEM[37][0] ),
    .B2(_09051_),
    .X(_05256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16066_ (.A(_09010_),
    .X(_09055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16067_ (.A1(_09005_),
    .A2(_10897_),
    .B1(_08019_),
    .B2(_09055_),
    .X(_09056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16068_ (.A(_09056_),
    .Y(_09057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16069_ (.A(_09057_),
    .X(_09058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16070_ (.A(_09056_),
    .X(_09059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16071_ (.A1(_00308_),
    .A2(_09058_),
    .B1(\design_top.MEM[24][7] ),
    .B2(_09059_),
    .X(_05255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16072_ (.A1(_00307_),
    .A2(_09058_),
    .B1(\design_top.MEM[24][6] ),
    .B2(_09059_),
    .X(_05254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16073_ (.A1(_00306_),
    .A2(_09058_),
    .B1(\design_top.MEM[24][5] ),
    .B2(_09059_),
    .X(_05253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16074_ (.A1(_00305_),
    .A2(_09058_),
    .B1(\design_top.MEM[24][4] ),
    .B2(_09059_),
    .X(_05252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16075_ (.A1(_00304_),
    .A2(_09058_),
    .B1(\design_top.MEM[24][3] ),
    .B2(_09059_),
    .X(_05251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16076_ (.A1(_00303_),
    .A2(_09057_),
    .B1(\design_top.MEM[24][2] ),
    .B2(_09056_),
    .X(_05250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16077_ (.A1(_00302_),
    .A2(_09057_),
    .B1(\design_top.MEM[24][1] ),
    .B2(_09056_),
    .X(_05249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16078_ (.A1(_00301_),
    .A2(_09057_),
    .B1(\design_top.MEM[24][0] ),
    .B2(_09056_),
    .X(_05248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16079_ (.A1(_09032_),
    .A2(_07519_),
    .B1(_07671_),
    .B2(_09055_),
    .X(_09060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16080_ (.A(_09060_),
    .Y(_09061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16081_ (.A(_09061_),
    .X(_09062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16082_ (.A(_09060_),
    .X(_09063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16083_ (.A1(_00428_),
    .A2(_09062_),
    .B1(\design_top.MEM[38][7] ),
    .B2(_09063_),
    .X(_05247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16084_ (.A1(_00427_),
    .A2(_09062_),
    .B1(\design_top.MEM[38][6] ),
    .B2(_09063_),
    .X(_05246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16085_ (.A1(_00426_),
    .A2(_09062_),
    .B1(\design_top.MEM[38][5] ),
    .B2(_09063_),
    .X(_05245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16086_ (.A1(_00425_),
    .A2(_09062_),
    .B1(\design_top.MEM[38][4] ),
    .B2(_09063_),
    .X(_05244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16087_ (.A1(_00424_),
    .A2(_09062_),
    .B1(\design_top.MEM[38][3] ),
    .B2(_09063_),
    .X(_05243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16088_ (.A1(_00423_),
    .A2(_09061_),
    .B1(\design_top.MEM[38][2] ),
    .B2(_09060_),
    .X(_05242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16089_ (.A1(_00422_),
    .A2(_09061_),
    .B1(\design_top.MEM[38][1] ),
    .B2(_09060_),
    .X(_05241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16090_ (.A1(_00421_),
    .A2(_09061_),
    .B1(\design_top.MEM[38][0] ),
    .B2(_09060_),
    .X(_05240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16091_ (.A1(_10898_),
    .A2(_11195_),
    .B1(_08044_),
    .B2(_09055_),
    .X(_09064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16092_ (.A(_09064_),
    .Y(_09065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16093_ (.A(_09065_),
    .X(_09066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16094_ (.A(_09064_),
    .X(_09067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16095_ (.A1(_00316_),
    .A2(_09066_),
    .B1(\design_top.MEM[25][7] ),
    .B2(_09067_),
    .X(_05239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16096_ (.A1(_00315_),
    .A2(_09066_),
    .B1(\design_top.MEM[25][6] ),
    .B2(_09067_),
    .X(_05238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16097_ (.A1(_00314_),
    .A2(_09066_),
    .B1(\design_top.MEM[25][5] ),
    .B2(_09067_),
    .X(_05237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16098_ (.A1(_00313_),
    .A2(_09066_),
    .B1(\design_top.MEM[25][4] ),
    .B2(_09067_),
    .X(_05236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16099_ (.A1(_00312_),
    .A2(_09066_),
    .B1(\design_top.MEM[25][3] ),
    .B2(_09067_),
    .X(_05235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16100_ (.A1(_00311_),
    .A2(_09065_),
    .B1(\design_top.MEM[25][2] ),
    .B2(_09064_),
    .X(_05234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16101_ (.A1(_00310_),
    .A2(_09065_),
    .B1(\design_top.MEM[25][1] ),
    .B2(_09064_),
    .X(_05233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16102_ (.A1(_00309_),
    .A2(_09065_),
    .B1(\design_top.MEM[25][0] ),
    .B2(_09064_),
    .X(_05232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16103_ (.A1(_10897_),
    .A2(_11134_),
    .B1(_08068_),
    .B2(_09055_),
    .X(_09068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16104_ (.A(_09068_),
    .Y(_09069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16105_ (.A(_09069_),
    .X(_09070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16106_ (.A(_09068_),
    .X(_09071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16107_ (.A1(_00324_),
    .A2(_09070_),
    .B1(\design_top.MEM[26][7] ),
    .B2(_09071_),
    .X(_05231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16108_ (.A1(_00323_),
    .A2(_09070_),
    .B1(\design_top.MEM[26][6] ),
    .B2(_09071_),
    .X(_05230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16109_ (.A1(_00322_),
    .A2(_09070_),
    .B1(\design_top.MEM[26][5] ),
    .B2(_09071_),
    .X(_05229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16110_ (.A1(_00321_),
    .A2(_09070_),
    .B1(\design_top.MEM[26][4] ),
    .B2(_09071_),
    .X(_05228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16111_ (.A1(_00320_),
    .A2(_09070_),
    .B1(\design_top.MEM[26][3] ),
    .B2(_09071_),
    .X(_05227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16112_ (.A1(_00319_),
    .A2(_09069_),
    .B1(\design_top.MEM[26][2] ),
    .B2(_09068_),
    .X(_05226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16113_ (.A1(_00318_),
    .A2(_09069_),
    .B1(\design_top.MEM[26][1] ),
    .B2(_09068_),
    .X(_05225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16114_ (.A1(_00317_),
    .A2(_09069_),
    .B1(\design_top.MEM[26][0] ),
    .B2(_09068_),
    .X(_05224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16115_ (.A1(_09050_),
    .A2(_11137_),
    .B1(_08103_),
    .B2(_09055_),
    .X(_09072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16116_ (.A(_09072_),
    .Y(_09073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16117_ (.A(_09073_),
    .X(_09074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16118_ (.A(_09072_),
    .X(_09075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16119_ (.A1(_00684_),
    .A2(_09074_),
    .B1(\design_top.MEM[9][7] ),
    .B2(_09075_),
    .X(_05223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16120_ (.A1(_00683_),
    .A2(_09074_),
    .B1(\design_top.MEM[9][6] ),
    .B2(_09075_),
    .X(_05222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16121_ (.A1(_00682_),
    .A2(_09074_),
    .B1(\design_top.MEM[9][5] ),
    .B2(_09075_),
    .X(_05221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16122_ (.A1(_00681_),
    .A2(_09074_),
    .B1(\design_top.MEM[9][4] ),
    .B2(_09075_),
    .X(_05220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16123_ (.A1(_00680_),
    .A2(_09074_),
    .B1(\design_top.MEM[9][3] ),
    .B2(_09075_),
    .X(_05219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16124_ (.A1(_00679_),
    .A2(_09073_),
    .B1(\design_top.MEM[9][2] ),
    .B2(_09072_),
    .X(_05218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16125_ (.A1(_00678_),
    .A2(_09073_),
    .B1(\design_top.MEM[9][1] ),
    .B2(_09072_),
    .X(_05217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16126_ (.A1(_00677_),
    .A2(_09073_),
    .B1(\design_top.MEM[9][0] ),
    .B2(_09072_),
    .X(_05216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16127_ (.A(_09010_),
    .X(_09076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16128_ (.A1(_09005_),
    .A2(_11137_),
    .B1(_08120_),
    .B2(_09076_),
    .X(_09077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16129_ (.A(_09077_),
    .Y(_09078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16130_ (.A(_09078_),
    .X(_09079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16131_ (.A(_09077_),
    .X(_09080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16132_ (.A1(_00676_),
    .A2(_09079_),
    .B1(\design_top.MEM[8][7] ),
    .B2(_09080_),
    .X(_05215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16133_ (.A1(_00675_),
    .A2(_09079_),
    .B1(\design_top.MEM[8][6] ),
    .B2(_09080_),
    .X(_05214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16134_ (.A1(_00674_),
    .A2(_09079_),
    .B1(\design_top.MEM[8][5] ),
    .B2(_09080_),
    .X(_05213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16135_ (.A1(_00673_),
    .A2(_09079_),
    .B1(\design_top.MEM[8][4] ),
    .B2(_09080_),
    .X(_05212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16136_ (.A1(_00672_),
    .A2(_09079_),
    .B1(\design_top.MEM[8][3] ),
    .B2(_09080_),
    .X(_05211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16137_ (.A1(_00671_),
    .A2(_09078_),
    .B1(\design_top.MEM[8][2] ),
    .B2(_09077_),
    .X(_05210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16138_ (.A1(_00670_),
    .A2(_09078_),
    .B1(\design_top.MEM[8][1] ),
    .B2(_09077_),
    .X(_05209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16139_ (.A1(_00669_),
    .A2(_09078_),
    .B1(\design_top.MEM[8][0] ),
    .B2(_09077_),
    .X(_05208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16140_ (.A(_08799_),
    .X(_09081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16141_ (.A(_09081_),
    .X(_09082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16142_ (.A(_00861_),
    .Y(_09083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16143_ (.A(_09083_),
    .X(_09084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16144_ (.A(_00860_),
    .X(_09085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16145_ (.A(_00862_),
    .Y(_09086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16146_ (.A(_09086_),
    .X(_09087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _16147_ (.A(_09084_),
    .B(_09085_),
    .C(_08781_),
    .D(_09087_),
    .X(_09088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16148_ (.A(_09088_),
    .X(_09089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16149_ (.A(_09089_),
    .X(_09090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16150_ (.A(_09090_),
    .X(_09091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16151_ (.A(_09089_),
    .Y(_09092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16152_ (.A(_09092_),
    .X(_09093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16153_ (.A(_09093_),
    .X(_09094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16154_ (.A1(_09082_),
    .A2(_09091_),
    .B1(\design_top.core0.REG2[14][31] ),
    .B2(_09094_),
    .X(_05207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16155_ (.A(_08801_),
    .X(_09095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16156_ (.A(_09095_),
    .X(_09096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16157_ (.A1(_09096_),
    .A2(_09091_),
    .B1(\design_top.core0.REG2[14][30] ),
    .B2(_09094_),
    .X(_05206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16158_ (.A(_08803_),
    .X(_09097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16159_ (.A(_09097_),
    .X(_09098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16160_ (.A1(_09098_),
    .A2(_09091_),
    .B1(\design_top.core0.REG2[14][29] ),
    .B2(_09094_),
    .X(_05205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16161_ (.A(_08805_),
    .X(_09099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16162_ (.A(_09099_),
    .X(_09100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16163_ (.A1(_09100_),
    .A2(_09091_),
    .B1(\design_top.core0.REG2[14][28] ),
    .B2(_09094_),
    .X(_05204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16164_ (.A(_08808_),
    .X(_09101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16165_ (.A(_09101_),
    .X(_09102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16166_ (.A1(_09102_),
    .A2(_09091_),
    .B1(\design_top.core0.REG2[14][27] ),
    .B2(_09094_),
    .X(_05203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16167_ (.A(_08812_),
    .X(_09103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16168_ (.A(_09103_),
    .X(_09104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16169_ (.A(_09090_),
    .X(_09105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16170_ (.A(_09093_),
    .X(_09106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16171_ (.A1(_09104_),
    .A2(_09105_),
    .B1(\design_top.core0.REG2[14][26] ),
    .B2(_09106_),
    .X(_05202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16172_ (.A(_08814_),
    .X(_09107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16173_ (.A(_09107_),
    .X(_09108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16174_ (.A1(_09108_),
    .A2(_09105_),
    .B1(\design_top.core0.REG2[14][25] ),
    .B2(_09106_),
    .X(_05201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16175_ (.A(_08816_),
    .X(_09109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16176_ (.A(_09109_),
    .X(_09110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16177_ (.A1(_09110_),
    .A2(_09105_),
    .B1(\design_top.core0.REG2[14][24] ),
    .B2(_09106_),
    .X(_05200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16178_ (.A(_08818_),
    .X(_09111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16179_ (.A(_09111_),
    .X(_09112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16180_ (.A1(_09112_),
    .A2(_09105_),
    .B1(\design_top.core0.REG2[14][23] ),
    .B2(_09106_),
    .X(_05199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16181_ (.A(_08821_),
    .X(_09113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16182_ (.A(_09113_),
    .X(_09114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16183_ (.A1(_09114_),
    .A2(_09105_),
    .B1(\design_top.core0.REG2[14][22] ),
    .B2(_09106_),
    .X(_05198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16184_ (.A(_08825_),
    .X(_09115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16185_ (.A(_09115_),
    .X(_09116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16186_ (.A(_09090_),
    .X(_09117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16187_ (.A(_09093_),
    .X(_09118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16188_ (.A1(_09116_),
    .A2(_09117_),
    .B1(\design_top.core0.REG2[14][21] ),
    .B2(_09118_),
    .X(_05197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16189_ (.A(_08827_),
    .X(_09119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16190_ (.A(_09119_),
    .X(_09120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16191_ (.A1(_09120_),
    .A2(_09117_),
    .B1(\design_top.core0.REG2[14][20] ),
    .B2(_09118_),
    .X(_05196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16192_ (.A(_08829_),
    .X(_09121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16193_ (.A(_09121_),
    .X(_09122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16194_ (.A1(_09122_),
    .A2(_09117_),
    .B1(\design_top.core0.REG2[14][19] ),
    .B2(_09118_),
    .X(_05195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16195_ (.A(_08831_),
    .X(_09123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16196_ (.A(_09123_),
    .X(_09124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16197_ (.A1(_09124_),
    .A2(_09117_),
    .B1(\design_top.core0.REG2[14][18] ),
    .B2(_09118_),
    .X(_05194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16198_ (.A(_08834_),
    .X(_09125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16199_ (.A(_09125_),
    .X(_09126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16200_ (.A1(_09126_),
    .A2(_09117_),
    .B1(\design_top.core0.REG2[14][17] ),
    .B2(_09118_),
    .X(_05193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16201_ (.A(_08838_),
    .X(_09127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16202_ (.A(_09127_),
    .X(_09128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16203_ (.A(_09089_),
    .X(_09129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16204_ (.A(_09092_),
    .X(_09130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16205_ (.A1(_09128_),
    .A2(_09129_),
    .B1(\design_top.core0.REG2[14][16] ),
    .B2(_09130_),
    .X(_05192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16206_ (.A(_08840_),
    .X(_09131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16207_ (.A(_09131_),
    .X(_09132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16208_ (.A1(_09132_),
    .A2(_09129_),
    .B1(\design_top.core0.REG2[14][15] ),
    .B2(_09130_),
    .X(_05191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16209_ (.A(_08842_),
    .X(_09133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16210_ (.A(_09133_),
    .X(_09134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16211_ (.A1(_09134_),
    .A2(_09129_),
    .B1(\design_top.core0.REG2[14][14] ),
    .B2(_09130_),
    .X(_05190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16212_ (.A(_08844_),
    .X(_09135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16213_ (.A1(\design_top.core0.REG2[14][13] ),
    .A2(_09090_),
    .B1(_09135_),
    .B2(_09093_),
    .X(_05189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16214_ (.A(_08845_),
    .X(_09136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16215_ (.A(_09136_),
    .X(_09137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16216_ (.A1(_09137_),
    .A2(_09129_),
    .B1(\design_top.core0.REG2[14][12] ),
    .B2(_09130_),
    .X(_05188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16217_ (.A(_08848_),
    .X(_09138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16218_ (.A(_09138_),
    .X(_09139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16219_ (.A1(_09139_),
    .A2(_09129_),
    .B1(\design_top.core0.REG2[14][11] ),
    .B2(_09130_),
    .X(_05187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16220_ (.A(_08852_),
    .X(_09140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16221_ (.A(_09140_),
    .X(_09141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16222_ (.A(_09089_),
    .X(_09142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16223_ (.A(_09092_),
    .X(_09143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16224_ (.A1(_09141_),
    .A2(_09142_),
    .B1(\design_top.core0.REG2[14][10] ),
    .B2(_09143_),
    .X(_05186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16225_ (.A(_08854_),
    .X(_09144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16226_ (.A(_09144_),
    .X(_09145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16227_ (.A1(_09145_),
    .A2(_09142_),
    .B1(\design_top.core0.REG2[14][9] ),
    .B2(_09143_),
    .X(_05185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16228_ (.A(_08856_),
    .X(_09146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16229_ (.A(_09146_),
    .X(_09147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16230_ (.A1(_09147_),
    .A2(_09142_),
    .B1(\design_top.core0.REG2[14][8] ),
    .B2(_09143_),
    .X(_05184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16231_ (.A(_08858_),
    .X(_09148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16232_ (.A(_09148_),
    .X(_09149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16233_ (.A1(_09149_),
    .A2(_09142_),
    .B1(\design_top.core0.REG2[14][7] ),
    .B2(_09143_),
    .X(_05183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16234_ (.A(_08861_),
    .X(_09150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16235_ (.A(_09150_),
    .X(_09151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16236_ (.A1(_09151_),
    .A2(_09142_),
    .B1(\design_top.core0.REG2[14][6] ),
    .B2(_09143_),
    .X(_05182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16237_ (.A(_08865_),
    .X(_09152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16238_ (.A(_09152_),
    .X(_09153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16239_ (.A(_09089_),
    .X(_09154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16240_ (.A(_09092_),
    .X(_09155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16241_ (.A1(_09153_),
    .A2(_09154_),
    .B1(\design_top.core0.REG2[14][5] ),
    .B2(_09155_),
    .X(_05181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16242_ (.A(_08867_),
    .X(_09156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16243_ (.A(_09156_),
    .X(_09157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16244_ (.A1(_09157_),
    .A2(_09154_),
    .B1(\design_top.core0.REG2[14][4] ),
    .B2(_09155_),
    .X(_05180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16245_ (.A(_08869_),
    .X(_09158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16246_ (.A(_09158_),
    .X(_09159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16247_ (.A1(_09159_),
    .A2(_09154_),
    .B1(\design_top.core0.REG2[14][3] ),
    .B2(_09155_),
    .X(_05179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16248_ (.A(_08871_),
    .X(_09160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16249_ (.A(_09160_),
    .X(_09161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16250_ (.A1(_09161_),
    .A2(_09154_),
    .B1(\design_top.core0.REG2[14][2] ),
    .B2(_09155_),
    .X(_05178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16251_ (.A(_08873_),
    .X(_09162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16252_ (.A(_09162_),
    .X(_09163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16253_ (.A1(_09163_),
    .A2(_09154_),
    .B1(\design_top.core0.REG2[14][1] ),
    .B2(_09155_),
    .X(_05177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16254_ (.A(_08875_),
    .X(_09164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16255_ (.A(_09164_),
    .X(_09165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16256_ (.A1(_09165_),
    .A2(_09090_),
    .B1(\design_top.core0.REG2[14][0] ),
    .B2(_09093_),
    .X(_05176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _16257_ (.A(_08778_),
    .B(_08780_),
    .C(_08781_),
    .D(_09087_),
    .X(_09166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16258_ (.A(_09166_),
    .X(_09167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16259_ (.A(_09167_),
    .X(_09168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16260_ (.A(_09168_),
    .X(_09169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16261_ (.A(_09167_),
    .Y(_09170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16262_ (.A(_09170_),
    .X(_09171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16263_ (.A(_09171_),
    .X(_09172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16264_ (.A1(_09082_),
    .A2(_09169_),
    .B1(\design_top.core0.REG2[13][31] ),
    .B2(_09172_),
    .X(_05175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16265_ (.A1(_09096_),
    .A2(_09169_),
    .B1(\design_top.core0.REG2[13][30] ),
    .B2(_09172_),
    .X(_05174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16266_ (.A1(_09098_),
    .A2(_09169_),
    .B1(\design_top.core0.REG2[13][29] ),
    .B2(_09172_),
    .X(_05173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16267_ (.A1(_09100_),
    .A2(_09169_),
    .B1(\design_top.core0.REG2[13][28] ),
    .B2(_09172_),
    .X(_05172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16268_ (.A1(_09102_),
    .A2(_09169_),
    .B1(\design_top.core0.REG2[13][27] ),
    .B2(_09172_),
    .X(_05171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16269_ (.A(_09168_),
    .X(_09173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16270_ (.A(_09171_),
    .X(_09174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16271_ (.A1(_09104_),
    .A2(_09173_),
    .B1(\design_top.core0.REG2[13][26] ),
    .B2(_09174_),
    .X(_05170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16272_ (.A1(_09108_),
    .A2(_09173_),
    .B1(\design_top.core0.REG2[13][25] ),
    .B2(_09174_),
    .X(_05169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16273_ (.A1(_09110_),
    .A2(_09173_),
    .B1(\design_top.core0.REG2[13][24] ),
    .B2(_09174_),
    .X(_05168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16274_ (.A1(_09112_),
    .A2(_09173_),
    .B1(\design_top.core0.REG2[13][23] ),
    .B2(_09174_),
    .X(_05167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16275_ (.A1(_09114_),
    .A2(_09173_),
    .B1(\design_top.core0.REG2[13][22] ),
    .B2(_09174_),
    .X(_05166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16276_ (.A(_09168_),
    .X(_09175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16277_ (.A(_09171_),
    .X(_09176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16278_ (.A1(_09116_),
    .A2(_09175_),
    .B1(\design_top.core0.REG2[13][21] ),
    .B2(_09176_),
    .X(_05165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16279_ (.A1(_09120_),
    .A2(_09175_),
    .B1(\design_top.core0.REG2[13][20] ),
    .B2(_09176_),
    .X(_05164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16280_ (.A1(_09122_),
    .A2(_09175_),
    .B1(\design_top.core0.REG2[13][19] ),
    .B2(_09176_),
    .X(_05163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16281_ (.A1(_09124_),
    .A2(_09175_),
    .B1(\design_top.core0.REG2[13][18] ),
    .B2(_09176_),
    .X(_05162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16282_ (.A1(_09126_),
    .A2(_09175_),
    .B1(\design_top.core0.REG2[13][17] ),
    .B2(_09176_),
    .X(_05161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16283_ (.A(_09167_),
    .X(_09177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16284_ (.A(_09170_),
    .X(_09178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16285_ (.A1(_09128_),
    .A2(_09177_),
    .B1(\design_top.core0.REG2[13][16] ),
    .B2(_09178_),
    .X(_05160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16286_ (.A1(_09132_),
    .A2(_09177_),
    .B1(\design_top.core0.REG2[13][15] ),
    .B2(_09178_),
    .X(_05159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16287_ (.A1(_09134_),
    .A2(_09177_),
    .B1(\design_top.core0.REG2[13][14] ),
    .B2(_09178_),
    .X(_05158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16288_ (.A1(\design_top.core0.REG2[13][13] ),
    .A2(_09168_),
    .B1(_09135_),
    .B2(_09171_),
    .X(_05157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16289_ (.A1(_09137_),
    .A2(_09177_),
    .B1(\design_top.core0.REG2[13][12] ),
    .B2(_09178_),
    .X(_05156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16290_ (.A1(_09139_),
    .A2(_09177_),
    .B1(\design_top.core0.REG2[13][11] ),
    .B2(_09178_),
    .X(_05155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16291_ (.A(_09167_),
    .X(_09179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16292_ (.A(_09170_),
    .X(_09180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16293_ (.A1(_09141_),
    .A2(_09179_),
    .B1(\design_top.core0.REG2[13][10] ),
    .B2(_09180_),
    .X(_05154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16294_ (.A1(_09145_),
    .A2(_09179_),
    .B1(\design_top.core0.REG2[13][9] ),
    .B2(_09180_),
    .X(_05153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16295_ (.A1(_09147_),
    .A2(_09179_),
    .B1(\design_top.core0.REG2[13][8] ),
    .B2(_09180_),
    .X(_05152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16296_ (.A1(_09149_),
    .A2(_09179_),
    .B1(\design_top.core0.REG2[13][7] ),
    .B2(_09180_),
    .X(_05151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16297_ (.A1(_09151_),
    .A2(_09179_),
    .B1(\design_top.core0.REG2[13][6] ),
    .B2(_09180_),
    .X(_05150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16298_ (.A(_09167_),
    .X(_09181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16299_ (.A(_09170_),
    .X(_09182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16300_ (.A1(_09153_),
    .A2(_09181_),
    .B1(\design_top.core0.REG2[13][5] ),
    .B2(_09182_),
    .X(_05149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16301_ (.A1(_09157_),
    .A2(_09181_),
    .B1(\design_top.core0.REG2[13][4] ),
    .B2(_09182_),
    .X(_05148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16302_ (.A1(_09159_),
    .A2(_09181_),
    .B1(\design_top.core0.REG2[13][3] ),
    .B2(_09182_),
    .X(_05147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16303_ (.A1(_09161_),
    .A2(_09181_),
    .B1(\design_top.core0.REG2[13][2] ),
    .B2(_09182_),
    .X(_05146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16304_ (.A1(_09163_),
    .A2(_09181_),
    .B1(\design_top.core0.REG2[13][1] ),
    .B2(_09182_),
    .X(_05145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16305_ (.A1(_09165_),
    .A2(_09168_),
    .B1(\design_top.core0.REG2[13][0] ),
    .B2(_09171_),
    .X(_05144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _16306_ (.A(_08778_),
    .B(_09085_),
    .C(_08781_),
    .D(_09087_),
    .X(_09183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16307_ (.A(_09183_),
    .X(_09184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16308_ (.A(_09184_),
    .X(_09185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16309_ (.A(_09185_),
    .X(_09186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16310_ (.A(_09184_),
    .Y(_09187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16311_ (.A(_09187_),
    .X(_09188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16312_ (.A(_09188_),
    .X(_09189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16313_ (.A1(_09082_),
    .A2(_09186_),
    .B1(\design_top.core0.REG2[12][31] ),
    .B2(_09189_),
    .X(_05143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16314_ (.A1(_09096_),
    .A2(_09186_),
    .B1(\design_top.core0.REG2[12][30] ),
    .B2(_09189_),
    .X(_05142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16315_ (.A1(_09098_),
    .A2(_09186_),
    .B1(\design_top.core0.REG2[12][29] ),
    .B2(_09189_),
    .X(_05141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16316_ (.A1(_09100_),
    .A2(_09186_),
    .B1(\design_top.core0.REG2[12][28] ),
    .B2(_09189_),
    .X(_05140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16317_ (.A1(_09102_),
    .A2(_09186_),
    .B1(\design_top.core0.REG2[12][27] ),
    .B2(_09189_),
    .X(_05139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16318_ (.A(_09185_),
    .X(_09190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16319_ (.A(_09188_),
    .X(_09191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16320_ (.A1(_09104_),
    .A2(_09190_),
    .B1(\design_top.core0.REG2[12][26] ),
    .B2(_09191_),
    .X(_05138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16321_ (.A1(_09108_),
    .A2(_09190_),
    .B1(\design_top.core0.REG2[12][25] ),
    .B2(_09191_),
    .X(_05137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16322_ (.A1(_09110_),
    .A2(_09190_),
    .B1(\design_top.core0.REG2[12][24] ),
    .B2(_09191_),
    .X(_05136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16323_ (.A1(_09112_),
    .A2(_09190_),
    .B1(\design_top.core0.REG2[12][23] ),
    .B2(_09191_),
    .X(_05135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16324_ (.A1(_09114_),
    .A2(_09190_),
    .B1(\design_top.core0.REG2[12][22] ),
    .B2(_09191_),
    .X(_05134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16325_ (.A(_09185_),
    .X(_09192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16326_ (.A(_09188_),
    .X(_09193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16327_ (.A1(_09116_),
    .A2(_09192_),
    .B1(\design_top.core0.REG2[12][21] ),
    .B2(_09193_),
    .X(_05133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16328_ (.A1(_09120_),
    .A2(_09192_),
    .B1(\design_top.core0.REG2[12][20] ),
    .B2(_09193_),
    .X(_05132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16329_ (.A1(_09122_),
    .A2(_09192_),
    .B1(\design_top.core0.REG2[12][19] ),
    .B2(_09193_),
    .X(_05131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16330_ (.A1(_09124_),
    .A2(_09192_),
    .B1(\design_top.core0.REG2[12][18] ),
    .B2(_09193_),
    .X(_05130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16331_ (.A1(_09126_),
    .A2(_09192_),
    .B1(\design_top.core0.REG2[12][17] ),
    .B2(_09193_),
    .X(_05129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16332_ (.A(_09184_),
    .X(_09194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16333_ (.A(_09187_),
    .X(_09195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16334_ (.A1(_09128_),
    .A2(_09194_),
    .B1(\design_top.core0.REG2[12][16] ),
    .B2(_09195_),
    .X(_05128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16335_ (.A1(_09132_),
    .A2(_09194_),
    .B1(\design_top.core0.REG2[12][15] ),
    .B2(_09195_),
    .X(_05127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16336_ (.A1(_09134_),
    .A2(_09194_),
    .B1(\design_top.core0.REG2[12][14] ),
    .B2(_09195_),
    .X(_05126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16337_ (.A1(\design_top.core0.REG2[12][13] ),
    .A2(_09185_),
    .B1(_09135_),
    .B2(_09188_),
    .X(_05125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16338_ (.A1(_09137_),
    .A2(_09194_),
    .B1(\design_top.core0.REG2[12][12] ),
    .B2(_09195_),
    .X(_05124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16339_ (.A1(_09139_),
    .A2(_09194_),
    .B1(\design_top.core0.REG2[12][11] ),
    .B2(_09195_),
    .X(_05123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16340_ (.A(_09184_),
    .X(_09196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16341_ (.A(_09187_),
    .X(_09197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16342_ (.A1(_09141_),
    .A2(_09196_),
    .B1(\design_top.core0.REG2[12][10] ),
    .B2(_09197_),
    .X(_05122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16343_ (.A1(_09145_),
    .A2(_09196_),
    .B1(\design_top.core0.REG2[12][9] ),
    .B2(_09197_),
    .X(_05121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16344_ (.A1(_09147_),
    .A2(_09196_),
    .B1(\design_top.core0.REG2[12][8] ),
    .B2(_09197_),
    .X(_05120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16345_ (.A1(_09149_),
    .A2(_09196_),
    .B1(\design_top.core0.REG2[12][7] ),
    .B2(_09197_),
    .X(_05119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16346_ (.A1(_09151_),
    .A2(_09196_),
    .B1(\design_top.core0.REG2[12][6] ),
    .B2(_09197_),
    .X(_05118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16347_ (.A(_09184_),
    .X(_09198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16348_ (.A(_09187_),
    .X(_09199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16349_ (.A1(_09153_),
    .A2(_09198_),
    .B1(\design_top.core0.REG2[12][5] ),
    .B2(_09199_),
    .X(_05117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16350_ (.A1(_09157_),
    .A2(_09198_),
    .B1(\design_top.core0.REG2[12][4] ),
    .B2(_09199_),
    .X(_05116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16351_ (.A1(_09159_),
    .A2(_09198_),
    .B1(\design_top.core0.REG2[12][3] ),
    .B2(_09199_),
    .X(_05115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16352_ (.A1(_09161_),
    .A2(_09198_),
    .B1(\design_top.core0.REG2[12][2] ),
    .B2(_09199_),
    .X(_05114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16353_ (.A1(_09163_),
    .A2(_09198_),
    .B1(\design_top.core0.REG2[12][1] ),
    .B2(_09199_),
    .X(_05113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16354_ (.A1(_09165_),
    .A2(_09185_),
    .B1(\design_top.core0.REG2[12][0] ),
    .B2(_09188_),
    .X(_05112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16355_ (.A(_00862_),
    .X(_09200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _16356_ (.A(_08782_),
    .B(_09200_),
    .C(_09084_),
    .D(_08779_),
    .X(_09201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16357_ (.A(_09201_),
    .X(_09202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16358_ (.A(_09202_),
    .X(_09203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16359_ (.A(_09203_),
    .X(_09204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16360_ (.A(_09202_),
    .Y(_09205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16361_ (.A(_09205_),
    .X(_09206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16362_ (.A(_09206_),
    .X(_09207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16363_ (.A1(_09082_),
    .A2(_09204_),
    .B1(\design_top.core0.REG2[11][31] ),
    .B2(_09207_),
    .X(_05111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16364_ (.A1(_09096_),
    .A2(_09204_),
    .B1(\design_top.core0.REG2[11][30] ),
    .B2(_09207_),
    .X(_05110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16365_ (.A1(_09098_),
    .A2(_09204_),
    .B1(\design_top.core0.REG2[11][29] ),
    .B2(_09207_),
    .X(_05109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16366_ (.A1(_09100_),
    .A2(_09204_),
    .B1(\design_top.core0.REG2[11][28] ),
    .B2(_09207_),
    .X(_05108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16367_ (.A1(_09102_),
    .A2(_09204_),
    .B1(\design_top.core0.REG2[11][27] ),
    .B2(_09207_),
    .X(_05107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16368_ (.A(_09203_),
    .X(_09208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16369_ (.A(_09206_),
    .X(_09209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16370_ (.A1(_09104_),
    .A2(_09208_),
    .B1(\design_top.core0.REG2[11][26] ),
    .B2(_09209_),
    .X(_05106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16371_ (.A1(_09108_),
    .A2(_09208_),
    .B1(\design_top.core0.REG2[11][25] ),
    .B2(_09209_),
    .X(_05105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16372_ (.A1(_09110_),
    .A2(_09208_),
    .B1(\design_top.core0.REG2[11][24] ),
    .B2(_09209_),
    .X(_05104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16373_ (.A1(_09112_),
    .A2(_09208_),
    .B1(\design_top.core0.REG2[11][23] ),
    .B2(_09209_),
    .X(_05103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16374_ (.A1(_09114_),
    .A2(_09208_),
    .B1(\design_top.core0.REG2[11][22] ),
    .B2(_09209_),
    .X(_05102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16375_ (.A(_09203_),
    .X(_09210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16376_ (.A(_09206_),
    .X(_09211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16377_ (.A1(_09116_),
    .A2(_09210_),
    .B1(\design_top.core0.REG2[11][21] ),
    .B2(_09211_),
    .X(_05101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16378_ (.A1(_09120_),
    .A2(_09210_),
    .B1(\design_top.core0.REG2[11][20] ),
    .B2(_09211_),
    .X(_05100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16379_ (.A1(_09122_),
    .A2(_09210_),
    .B1(\design_top.core0.REG2[11][19] ),
    .B2(_09211_),
    .X(_05099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16380_ (.A1(_09124_),
    .A2(_09210_),
    .B1(\design_top.core0.REG2[11][18] ),
    .B2(_09211_),
    .X(_05098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16381_ (.A1(_09126_),
    .A2(_09210_),
    .B1(\design_top.core0.REG2[11][17] ),
    .B2(_09211_),
    .X(_05097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16382_ (.A(_09202_),
    .X(_09212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16383_ (.A(_09205_),
    .X(_09213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16384_ (.A1(_09128_),
    .A2(_09212_),
    .B1(\design_top.core0.REG2[11][16] ),
    .B2(_09213_),
    .X(_05096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16385_ (.A1(_09132_),
    .A2(_09212_),
    .B1(\design_top.core0.REG2[11][15] ),
    .B2(_09213_),
    .X(_05095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16386_ (.A1(_09134_),
    .A2(_09212_),
    .B1(\design_top.core0.REG2[11][14] ),
    .B2(_09213_),
    .X(_05094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16387_ (.A1(\design_top.core0.REG2[11][13] ),
    .A2(_09203_),
    .B1(_09135_),
    .B2(_09206_),
    .X(_05093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16388_ (.A1(_09137_),
    .A2(_09212_),
    .B1(\design_top.core0.REG2[11][12] ),
    .B2(_09213_),
    .X(_05092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16389_ (.A1(_09139_),
    .A2(_09212_),
    .B1(\design_top.core0.REG2[11][11] ),
    .B2(_09213_),
    .X(_05091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16390_ (.A(_09202_),
    .X(_09214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16391_ (.A(_09205_),
    .X(_09215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16392_ (.A1(_09141_),
    .A2(_09214_),
    .B1(\design_top.core0.REG2[11][10] ),
    .B2(_09215_),
    .X(_05090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16393_ (.A1(_09145_),
    .A2(_09214_),
    .B1(\design_top.core0.REG2[11][9] ),
    .B2(_09215_),
    .X(_05089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16394_ (.A1(_09147_),
    .A2(_09214_),
    .B1(\design_top.core0.REG2[11][8] ),
    .B2(_09215_),
    .X(_05088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16395_ (.A1(_09149_),
    .A2(_09214_),
    .B1(\design_top.core0.REG2[11][7] ),
    .B2(_09215_),
    .X(_05087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16396_ (.A1(_09151_),
    .A2(_09214_),
    .B1(\design_top.core0.REG2[11][6] ),
    .B2(_09215_),
    .X(_05086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16397_ (.A(_09202_),
    .X(_09216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16398_ (.A(_09205_),
    .X(_09217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16399_ (.A1(_09153_),
    .A2(_09216_),
    .B1(\design_top.core0.REG2[11][5] ),
    .B2(_09217_),
    .X(_05085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16400_ (.A1(_09157_),
    .A2(_09216_),
    .B1(\design_top.core0.REG2[11][4] ),
    .B2(_09217_),
    .X(_05084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16401_ (.A1(_09159_),
    .A2(_09216_),
    .B1(\design_top.core0.REG2[11][3] ),
    .B2(_09217_),
    .X(_05083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16402_ (.A1(_09161_),
    .A2(_09216_),
    .B1(\design_top.core0.REG2[11][2] ),
    .B2(_09217_),
    .X(_05082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16403_ (.A1(_09163_),
    .A2(_09216_),
    .B1(\design_top.core0.REG2[11][1] ),
    .B2(_09217_),
    .X(_05081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16404_ (.A1(_09165_),
    .A2(_09203_),
    .B1(\design_top.core0.REG2[11][0] ),
    .B2(_09206_),
    .X(_05080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _16405_ (.A(_08782_),
    .B(_09200_),
    .C(_09084_),
    .D(_09085_),
    .X(_09218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16406_ (.A(_09218_),
    .X(_09219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16407_ (.A(_09219_),
    .X(_09220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16408_ (.A(_09220_),
    .X(_09221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16409_ (.A(_09219_),
    .Y(_09222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16410_ (.A(_09222_),
    .X(_09223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16411_ (.A(_09223_),
    .X(_09224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16412_ (.A1(_09082_),
    .A2(_09221_),
    .B1(\design_top.core0.REG2[10][31] ),
    .B2(_09224_),
    .X(_05079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16413_ (.A1(_09096_),
    .A2(_09221_),
    .B1(\design_top.core0.REG2[10][30] ),
    .B2(_09224_),
    .X(_05078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16414_ (.A1(_09098_),
    .A2(_09221_),
    .B1(\design_top.core0.REG2[10][29] ),
    .B2(_09224_),
    .X(_05077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16415_ (.A1(_09100_),
    .A2(_09221_),
    .B1(\design_top.core0.REG2[10][28] ),
    .B2(_09224_),
    .X(_05076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16416_ (.A1(_09102_),
    .A2(_09221_),
    .B1(\design_top.core0.REG2[10][27] ),
    .B2(_09224_),
    .X(_05075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16417_ (.A(_09220_),
    .X(_09225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16418_ (.A(_09223_),
    .X(_09226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16419_ (.A1(_09104_),
    .A2(_09225_),
    .B1(\design_top.core0.REG2[10][26] ),
    .B2(_09226_),
    .X(_05074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16420_ (.A1(_09108_),
    .A2(_09225_),
    .B1(\design_top.core0.REG2[10][25] ),
    .B2(_09226_),
    .X(_05073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16421_ (.A1(_09110_),
    .A2(_09225_),
    .B1(\design_top.core0.REG2[10][24] ),
    .B2(_09226_),
    .X(_05072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16422_ (.A1(_09112_),
    .A2(_09225_),
    .B1(\design_top.core0.REG2[10][23] ),
    .B2(_09226_),
    .X(_05071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16423_ (.A1(_09114_),
    .A2(_09225_),
    .B1(\design_top.core0.REG2[10][22] ),
    .B2(_09226_),
    .X(_05070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16424_ (.A(_09220_),
    .X(_09227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16425_ (.A(_09223_),
    .X(_09228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16426_ (.A1(_09116_),
    .A2(_09227_),
    .B1(\design_top.core0.REG2[10][21] ),
    .B2(_09228_),
    .X(_05069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16427_ (.A1(_09120_),
    .A2(_09227_),
    .B1(\design_top.core0.REG2[10][20] ),
    .B2(_09228_),
    .X(_05068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16428_ (.A1(_09122_),
    .A2(_09227_),
    .B1(\design_top.core0.REG2[10][19] ),
    .B2(_09228_),
    .X(_05067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16429_ (.A1(_09124_),
    .A2(_09227_),
    .B1(\design_top.core0.REG2[10][18] ),
    .B2(_09228_),
    .X(_05066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16430_ (.A1(_09126_),
    .A2(_09227_),
    .B1(\design_top.core0.REG2[10][17] ),
    .B2(_09228_),
    .X(_05065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16431_ (.A(_09219_),
    .X(_09229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16432_ (.A(_09222_),
    .X(_09230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16433_ (.A1(_09128_),
    .A2(_09229_),
    .B1(\design_top.core0.REG2[10][16] ),
    .B2(_09230_),
    .X(_05064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16434_ (.A1(_09132_),
    .A2(_09229_),
    .B1(\design_top.core0.REG2[10][15] ),
    .B2(_09230_),
    .X(_05063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16435_ (.A1(_09134_),
    .A2(_09229_),
    .B1(\design_top.core0.REG2[10][14] ),
    .B2(_09230_),
    .X(_05062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16436_ (.A1(\design_top.core0.REG2[10][13] ),
    .A2(_09220_),
    .B1(_09135_),
    .B2(_09223_),
    .X(_05061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16437_ (.A1(_09137_),
    .A2(_09229_),
    .B1(\design_top.core0.REG2[10][12] ),
    .B2(_09230_),
    .X(_05060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16438_ (.A1(_09139_),
    .A2(_09229_),
    .B1(\design_top.core0.REG2[10][11] ),
    .B2(_09230_),
    .X(_05059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16439_ (.A(_09219_),
    .X(_09231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16440_ (.A(_09222_),
    .X(_09232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16441_ (.A1(_09141_),
    .A2(_09231_),
    .B1(\design_top.core0.REG2[10][10] ),
    .B2(_09232_),
    .X(_05058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16442_ (.A1(_09145_),
    .A2(_09231_),
    .B1(\design_top.core0.REG2[10][9] ),
    .B2(_09232_),
    .X(_05057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16443_ (.A1(_09147_),
    .A2(_09231_),
    .B1(\design_top.core0.REG2[10][8] ),
    .B2(_09232_),
    .X(_05056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16444_ (.A1(_09149_),
    .A2(_09231_),
    .B1(\design_top.core0.REG2[10][7] ),
    .B2(_09232_),
    .X(_05055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16445_ (.A1(_09151_),
    .A2(_09231_),
    .B1(\design_top.core0.REG2[10][6] ),
    .B2(_09232_),
    .X(_05054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16446_ (.A(_09219_),
    .X(_09233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16447_ (.A(_09222_),
    .X(_09234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16448_ (.A1(_09153_),
    .A2(_09233_),
    .B1(\design_top.core0.REG2[10][5] ),
    .B2(_09234_),
    .X(_05053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16449_ (.A1(_09157_),
    .A2(_09233_),
    .B1(\design_top.core0.REG2[10][4] ),
    .B2(_09234_),
    .X(_05052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16450_ (.A1(_09159_),
    .A2(_09233_),
    .B1(\design_top.core0.REG2[10][3] ),
    .B2(_09234_),
    .X(_05051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16451_ (.A1(_09161_),
    .A2(_09233_),
    .B1(\design_top.core0.REG2[10][2] ),
    .B2(_09234_),
    .X(_05050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16452_ (.A1(_09163_),
    .A2(_09233_),
    .B1(\design_top.core0.REG2[10][1] ),
    .B2(_09234_),
    .X(_05049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16453_ (.A1(_09165_),
    .A2(_09220_),
    .B1(\design_top.core0.REG2[10][0] ),
    .B2(_09223_),
    .X(_05048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16454_ (.A(_08786_),
    .X(_09235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16455_ (.A(_09235_),
    .X(_09236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16456_ (.A(_09236_),
    .X(_09237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16457_ (.A(\design_top.core0.REG2[0][31] ),
    .B(_09237_),
    .X(_05047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16458_ (.A(\design_top.core0.REG2[0][30] ),
    .B(_09237_),
    .X(_05046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16459_ (.A(\design_top.core0.REG2[0][29] ),
    .B(_09237_),
    .X(_05045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16460_ (.A(\design_top.core0.REG2[0][28] ),
    .B(_09237_),
    .X(_05044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16461_ (.A(\design_top.core0.REG2[0][27] ),
    .B(_09237_),
    .X(_05043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16462_ (.A(_09236_),
    .X(_09238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16463_ (.A(\design_top.core0.REG2[0][26] ),
    .B(_09238_),
    .X(_05042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16464_ (.A(\design_top.core0.REG2[0][25] ),
    .B(_09238_),
    .X(_05041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16465_ (.A(\design_top.core0.REG2[0][24] ),
    .B(_09238_),
    .X(_05040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16466_ (.A(\design_top.core0.REG2[0][23] ),
    .B(_09238_),
    .X(_05039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16467_ (.A(\design_top.core0.REG2[0][22] ),
    .B(_09238_),
    .X(_05038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16468_ (.A(_09236_),
    .X(_09239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16469_ (.A(\design_top.core0.REG2[0][21] ),
    .B(_09239_),
    .X(_05037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16470_ (.A(\design_top.core0.REG2[0][20] ),
    .B(_09239_),
    .X(_05036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16471_ (.A(\design_top.core0.REG2[0][19] ),
    .B(_09239_),
    .X(_05035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16472_ (.A(\design_top.core0.REG2[0][18] ),
    .B(_09239_),
    .X(_05034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16473_ (.A(\design_top.core0.REG2[0][17] ),
    .B(_09239_),
    .X(_05033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16474_ (.A(_09235_),
    .X(_09240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16475_ (.A(\design_top.core0.REG2[0][16] ),
    .B(_09240_),
    .X(_05032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16476_ (.A(\design_top.core0.REG2[0][15] ),
    .B(_09240_),
    .X(_05031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16477_ (.A(\design_top.core0.REG2[0][14] ),
    .B(_09240_),
    .X(_05030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16478_ (.A(_08844_),
    .X(_09241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16479_ (.A1(\design_top.core0.REG2[0][13] ),
    .A2(_09236_),
    .B1(_09241_),
    .B2(_08787_),
    .X(_05029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16480_ (.A(\design_top.core0.REG2[0][12] ),
    .B(_09240_),
    .X(_05028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16481_ (.A(\design_top.core0.REG2[0][11] ),
    .B(_09240_),
    .X(_05027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16482_ (.A(_09235_),
    .X(_09242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16483_ (.A(\design_top.core0.REG2[0][10] ),
    .B(_09242_),
    .X(_05026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16484_ (.A(\design_top.core0.REG2[0][9] ),
    .B(_09242_),
    .X(_05025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16485_ (.A(\design_top.core0.REG2[0][8] ),
    .B(_09242_),
    .X(_05024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16486_ (.A(\design_top.core0.REG2[0][7] ),
    .B(_09242_),
    .X(_05023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16487_ (.A(\design_top.core0.REG2[0][6] ),
    .B(_09242_),
    .X(_05022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16488_ (.A(_09235_),
    .X(_09243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16489_ (.A(\design_top.core0.REG2[0][5] ),
    .B(_09243_),
    .X(_05021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16490_ (.A(\design_top.core0.REG2[0][4] ),
    .B(_09243_),
    .X(_05020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16491_ (.A(\design_top.core0.REG2[0][3] ),
    .B(_09243_),
    .X(_05019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16492_ (.A(\design_top.core0.REG2[0][2] ),
    .B(_09243_),
    .X(_05018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16493_ (.A(\design_top.core0.REG2[0][1] ),
    .B(_09243_),
    .X(_05017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _16494_ (.A(\design_top.core0.REG2[0][0] ),
    .B(_09236_),
    .X(_05016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16495_ (.A(_09081_),
    .X(_09244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _16496_ (.A(_08782_),
    .B(_09200_),
    .C(_00861_),
    .D(_00860_),
    .X(_09245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16497_ (.A(_09245_),
    .X(_09246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16498_ (.A(_09246_),
    .X(_09247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16499_ (.A(_09247_),
    .X(_09248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16500_ (.A(_09246_),
    .Y(_09249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16501_ (.A(_09249_),
    .X(_09250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16502_ (.A(_09250_),
    .X(_09251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16503_ (.A1(_09244_),
    .A2(_09248_),
    .B1(\design_top.core0.REG2[8][31] ),
    .B2(_09251_),
    .X(_05015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16504_ (.A(_09095_),
    .X(_09252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16505_ (.A1(_09252_),
    .A2(_09248_),
    .B1(\design_top.core0.REG2[8][30] ),
    .B2(_09251_),
    .X(_05014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16506_ (.A(_09097_),
    .X(_09253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16507_ (.A1(_09253_),
    .A2(_09248_),
    .B1(\design_top.core0.REG2[8][29] ),
    .B2(_09251_),
    .X(_05013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16508_ (.A(_09099_),
    .X(_09254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16509_ (.A1(_09254_),
    .A2(_09248_),
    .B1(\design_top.core0.REG2[8][28] ),
    .B2(_09251_),
    .X(_05012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16510_ (.A(_09101_),
    .X(_09255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16511_ (.A1(_09255_),
    .A2(_09248_),
    .B1(\design_top.core0.REG2[8][27] ),
    .B2(_09251_),
    .X(_05011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16512_ (.A(_09103_),
    .X(_09256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16513_ (.A(_09247_),
    .X(_09257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16514_ (.A(_09250_),
    .X(_09258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16515_ (.A1(_09256_),
    .A2(_09257_),
    .B1(\design_top.core0.REG2[8][26] ),
    .B2(_09258_),
    .X(_05010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16516_ (.A(_09107_),
    .X(_09259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16517_ (.A1(_09259_),
    .A2(_09257_),
    .B1(\design_top.core0.REG2[8][25] ),
    .B2(_09258_),
    .X(_05009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16518_ (.A(_09109_),
    .X(_09260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16519_ (.A1(_09260_),
    .A2(_09257_),
    .B1(\design_top.core0.REG2[8][24] ),
    .B2(_09258_),
    .X(_05008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16520_ (.A(_09111_),
    .X(_09261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16521_ (.A1(_09261_),
    .A2(_09257_),
    .B1(\design_top.core0.REG2[8][23] ),
    .B2(_09258_),
    .X(_05007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16522_ (.A(_09113_),
    .X(_09262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16523_ (.A1(_09262_),
    .A2(_09257_),
    .B1(\design_top.core0.REG2[8][22] ),
    .B2(_09258_),
    .X(_05006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16524_ (.A(_09115_),
    .X(_09263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16525_ (.A(_09247_),
    .X(_09264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16526_ (.A(_09250_),
    .X(_09265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16527_ (.A1(_09263_),
    .A2(_09264_),
    .B1(\design_top.core0.REG2[8][21] ),
    .B2(_09265_),
    .X(_05005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16528_ (.A(_09119_),
    .X(_09266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16529_ (.A1(_09266_),
    .A2(_09264_),
    .B1(\design_top.core0.REG2[8][20] ),
    .B2(_09265_),
    .X(_05004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16530_ (.A(_09121_),
    .X(_09267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16531_ (.A1(_09267_),
    .A2(_09264_),
    .B1(\design_top.core0.REG2[8][19] ),
    .B2(_09265_),
    .X(_05003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16532_ (.A(_09123_),
    .X(_09268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16533_ (.A1(_09268_),
    .A2(_09264_),
    .B1(\design_top.core0.REG2[8][18] ),
    .B2(_09265_),
    .X(_05002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16534_ (.A(_09125_),
    .X(_09269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16535_ (.A1(_09269_),
    .A2(_09264_),
    .B1(\design_top.core0.REG2[8][17] ),
    .B2(_09265_),
    .X(_05001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16536_ (.A(_09127_),
    .X(_09270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16537_ (.A(_09246_),
    .X(_09271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16538_ (.A(_09249_),
    .X(_09272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16539_ (.A1(_09270_),
    .A2(_09271_),
    .B1(\design_top.core0.REG2[8][16] ),
    .B2(_09272_),
    .X(_05000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16540_ (.A(_09131_),
    .X(_09273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16541_ (.A1(_09273_),
    .A2(_09271_),
    .B1(\design_top.core0.REG2[8][15] ),
    .B2(_09272_),
    .X(_04999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16542_ (.A(_09133_),
    .X(_09274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16543_ (.A1(_09274_),
    .A2(_09271_),
    .B1(\design_top.core0.REG2[8][14] ),
    .B2(_09272_),
    .X(_04998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16544_ (.A1(\design_top.core0.REG2[8][13] ),
    .A2(_09247_),
    .B1(_09241_),
    .B2(_09250_),
    .X(_04997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16545_ (.A(_09136_),
    .X(_09275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16546_ (.A1(_09275_),
    .A2(_09271_),
    .B1(\design_top.core0.REG2[8][12] ),
    .B2(_09272_),
    .X(_04996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16547_ (.A(_09138_),
    .X(_09276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16548_ (.A1(_09276_),
    .A2(_09271_),
    .B1(\design_top.core0.REG2[8][11] ),
    .B2(_09272_),
    .X(_04995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16549_ (.A(_09140_),
    .X(_09277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16550_ (.A(_09246_),
    .X(_09278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16551_ (.A(_09249_),
    .X(_09279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16552_ (.A1(_09277_),
    .A2(_09278_),
    .B1(\design_top.core0.REG2[8][10] ),
    .B2(_09279_),
    .X(_04994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16553_ (.A(_09144_),
    .X(_09280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16554_ (.A1(_09280_),
    .A2(_09278_),
    .B1(\design_top.core0.REG2[8][9] ),
    .B2(_09279_),
    .X(_04993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16555_ (.A(_09146_),
    .X(_09281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16556_ (.A1(_09281_),
    .A2(_09278_),
    .B1(\design_top.core0.REG2[8][8] ),
    .B2(_09279_),
    .X(_04992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16557_ (.A(_09148_),
    .X(_09282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16558_ (.A1(_09282_),
    .A2(_09278_),
    .B1(\design_top.core0.REG2[8][7] ),
    .B2(_09279_),
    .X(_04991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16559_ (.A(_09150_),
    .X(_09283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16560_ (.A1(_09283_),
    .A2(_09278_),
    .B1(\design_top.core0.REG2[8][6] ),
    .B2(_09279_),
    .X(_04990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16561_ (.A(_09152_),
    .X(_09284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16562_ (.A(_09246_),
    .X(_09285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16563_ (.A(_09249_),
    .X(_09286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16564_ (.A1(_09284_),
    .A2(_09285_),
    .B1(\design_top.core0.REG2[8][5] ),
    .B2(_09286_),
    .X(_04989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16565_ (.A(_09156_),
    .X(_09287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16566_ (.A1(_09287_),
    .A2(_09285_),
    .B1(\design_top.core0.REG2[8][4] ),
    .B2(_09286_),
    .X(_04988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16567_ (.A(_09158_),
    .X(_09288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16568_ (.A1(_09288_),
    .A2(_09285_),
    .B1(\design_top.core0.REG2[8][3] ),
    .B2(_09286_),
    .X(_04987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16569_ (.A(_09160_),
    .X(_09289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16570_ (.A1(_09289_),
    .A2(_09285_),
    .B1(\design_top.core0.REG2[8][2] ),
    .B2(_09286_),
    .X(_04986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16571_ (.A(_09162_),
    .X(_09290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16572_ (.A1(_09290_),
    .A2(_09285_),
    .B1(\design_top.core0.REG2[8][1] ),
    .B2(_09286_),
    .X(_04985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16573_ (.A(_09164_),
    .X(_09291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16574_ (.A1(_09291_),
    .A2(_09247_),
    .B1(\design_top.core0.REG2[8][0] ),
    .B2(_09250_),
    .X(_04984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16575_ (.A(_00863_),
    .X(_09292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _16576_ (.A(_09084_),
    .B(_08780_),
    .C(_09292_),
    .D(_09087_),
    .X(_09293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16577_ (.A(_09293_),
    .X(_09294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16578_ (.A(_09294_),
    .X(_09295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16579_ (.A(_09295_),
    .X(_09296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16580_ (.A(_09294_),
    .Y(_09297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16581_ (.A(_09297_),
    .X(_09298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16582_ (.A(_09298_),
    .X(_09299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16583_ (.A1(_09244_),
    .A2(_09296_),
    .B1(\design_top.core0.REG2[7][31] ),
    .B2(_09299_),
    .X(_04983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16584_ (.A1(_09252_),
    .A2(_09296_),
    .B1(\design_top.core0.REG2[7][30] ),
    .B2(_09299_),
    .X(_04982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16585_ (.A1(_09253_),
    .A2(_09296_),
    .B1(\design_top.core0.REG2[7][29] ),
    .B2(_09299_),
    .X(_04981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16586_ (.A1(_09254_),
    .A2(_09296_),
    .B1(\design_top.core0.REG2[7][28] ),
    .B2(_09299_),
    .X(_04980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16587_ (.A1(_09255_),
    .A2(_09296_),
    .B1(\design_top.core0.REG2[7][27] ),
    .B2(_09299_),
    .X(_04979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16588_ (.A(_09295_),
    .X(_09300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16589_ (.A(_09298_),
    .X(_09301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16590_ (.A1(_09256_),
    .A2(_09300_),
    .B1(\design_top.core0.REG2[7][26] ),
    .B2(_09301_),
    .X(_04978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16591_ (.A1(_09259_),
    .A2(_09300_),
    .B1(\design_top.core0.REG2[7][25] ),
    .B2(_09301_),
    .X(_04977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16592_ (.A1(_09260_),
    .A2(_09300_),
    .B1(\design_top.core0.REG2[7][24] ),
    .B2(_09301_),
    .X(_04976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16593_ (.A1(_09261_),
    .A2(_09300_),
    .B1(\design_top.core0.REG2[7][23] ),
    .B2(_09301_),
    .X(_04975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16594_ (.A1(_09262_),
    .A2(_09300_),
    .B1(\design_top.core0.REG2[7][22] ),
    .B2(_09301_),
    .X(_04974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16595_ (.A(_09295_),
    .X(_09302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16596_ (.A(_09298_),
    .X(_09303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16597_ (.A1(_09263_),
    .A2(_09302_),
    .B1(\design_top.core0.REG2[7][21] ),
    .B2(_09303_),
    .X(_04973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16598_ (.A1(_09266_),
    .A2(_09302_),
    .B1(\design_top.core0.REG2[7][20] ),
    .B2(_09303_),
    .X(_04972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16599_ (.A1(_09267_),
    .A2(_09302_),
    .B1(\design_top.core0.REG2[7][19] ),
    .B2(_09303_),
    .X(_04971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16600_ (.A1(_09268_),
    .A2(_09302_),
    .B1(\design_top.core0.REG2[7][18] ),
    .B2(_09303_),
    .X(_04970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16601_ (.A1(_09269_),
    .A2(_09302_),
    .B1(\design_top.core0.REG2[7][17] ),
    .B2(_09303_),
    .X(_04969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16602_ (.A(_09294_),
    .X(_09304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16603_ (.A(_09297_),
    .X(_09305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16604_ (.A1(_09270_),
    .A2(_09304_),
    .B1(\design_top.core0.REG2[7][16] ),
    .B2(_09305_),
    .X(_04968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16605_ (.A1(_09273_),
    .A2(_09304_),
    .B1(\design_top.core0.REG2[7][15] ),
    .B2(_09305_),
    .X(_04967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16606_ (.A1(_09274_),
    .A2(_09304_),
    .B1(\design_top.core0.REG2[7][14] ),
    .B2(_09305_),
    .X(_04966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16607_ (.A1(\design_top.core0.REG2[7][13] ),
    .A2(_09295_),
    .B1(_09241_),
    .B2(_09298_),
    .X(_04965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16608_ (.A1(_09275_),
    .A2(_09304_),
    .B1(\design_top.core0.REG2[7][12] ),
    .B2(_09305_),
    .X(_04964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16609_ (.A1(_09276_),
    .A2(_09304_),
    .B1(\design_top.core0.REG2[7][11] ),
    .B2(_09305_),
    .X(_04963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16610_ (.A(_09294_),
    .X(_09306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16611_ (.A(_09297_),
    .X(_09307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16612_ (.A1(_09277_),
    .A2(_09306_),
    .B1(\design_top.core0.REG2[7][10] ),
    .B2(_09307_),
    .X(_04962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16613_ (.A1(_09280_),
    .A2(_09306_),
    .B1(\design_top.core0.REG2[7][9] ),
    .B2(_09307_),
    .X(_04961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16614_ (.A1(_09281_),
    .A2(_09306_),
    .B1(\design_top.core0.REG2[7][8] ),
    .B2(_09307_),
    .X(_04960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16615_ (.A1(_09282_),
    .A2(_09306_),
    .B1(\design_top.core0.REG2[7][7] ),
    .B2(_09307_),
    .X(_04959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16616_ (.A1(_09283_),
    .A2(_09306_),
    .B1(\design_top.core0.REG2[7][6] ),
    .B2(_09307_),
    .X(_04958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16617_ (.A(_09294_),
    .X(_09308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16618_ (.A(_09297_),
    .X(_09309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16619_ (.A1(_09284_),
    .A2(_09308_),
    .B1(\design_top.core0.REG2[7][5] ),
    .B2(_09309_),
    .X(_04957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16620_ (.A1(_09287_),
    .A2(_09308_),
    .B1(\design_top.core0.REG2[7][4] ),
    .B2(_09309_),
    .X(_04956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16621_ (.A1(_09288_),
    .A2(_09308_),
    .B1(\design_top.core0.REG2[7][3] ),
    .B2(_09309_),
    .X(_04955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16622_ (.A1(_09289_),
    .A2(_09308_),
    .B1(\design_top.core0.REG2[7][2] ),
    .B2(_09309_),
    .X(_04954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16623_ (.A1(_09290_),
    .A2(_09308_),
    .B1(\design_top.core0.REG2[7][1] ),
    .B2(_09309_),
    .X(_04953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16624_ (.A1(_09291_),
    .A2(_09295_),
    .B1(\design_top.core0.REG2[7][0] ),
    .B2(_09298_),
    .X(_04952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _16625_ (.A(_09084_),
    .B(_09085_),
    .C(_09292_),
    .D(_09086_),
    .X(_09310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16626_ (.A(_09310_),
    .X(_09311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16627_ (.A(_09311_),
    .X(_09312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16628_ (.A(_09312_),
    .X(_09313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16629_ (.A(_09311_),
    .Y(_09314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16630_ (.A(_09314_),
    .X(_09315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16631_ (.A(_09315_),
    .X(_09316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16632_ (.A1(_09244_),
    .A2(_09313_),
    .B1(\design_top.core0.REG2[6][31] ),
    .B2(_09316_),
    .X(_04951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16633_ (.A1(_09252_),
    .A2(_09313_),
    .B1(\design_top.core0.REG2[6][30] ),
    .B2(_09316_),
    .X(_04950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16634_ (.A1(_09253_),
    .A2(_09313_),
    .B1(\design_top.core0.REG2[6][29] ),
    .B2(_09316_),
    .X(_04949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16635_ (.A1(_09254_),
    .A2(_09313_),
    .B1(\design_top.core0.REG2[6][28] ),
    .B2(_09316_),
    .X(_04948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16636_ (.A1(_09255_),
    .A2(_09313_),
    .B1(\design_top.core0.REG2[6][27] ),
    .B2(_09316_),
    .X(_04947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16637_ (.A(_09312_),
    .X(_09317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16638_ (.A(_09315_),
    .X(_09318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16639_ (.A1(_09256_),
    .A2(_09317_),
    .B1(\design_top.core0.REG2[6][26] ),
    .B2(_09318_),
    .X(_04946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16640_ (.A1(_09259_),
    .A2(_09317_),
    .B1(\design_top.core0.REG2[6][25] ),
    .B2(_09318_),
    .X(_04945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16641_ (.A1(_09260_),
    .A2(_09317_),
    .B1(\design_top.core0.REG2[6][24] ),
    .B2(_09318_),
    .X(_04944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16642_ (.A1(_09261_),
    .A2(_09317_),
    .B1(\design_top.core0.REG2[6][23] ),
    .B2(_09318_),
    .X(_04943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16643_ (.A1(_09262_),
    .A2(_09317_),
    .B1(\design_top.core0.REG2[6][22] ),
    .B2(_09318_),
    .X(_04942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16644_ (.A(_09312_),
    .X(_09319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16645_ (.A(_09315_),
    .X(_09320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16646_ (.A1(_09263_),
    .A2(_09319_),
    .B1(\design_top.core0.REG2[6][21] ),
    .B2(_09320_),
    .X(_04941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16647_ (.A1(_09266_),
    .A2(_09319_),
    .B1(\design_top.core0.REG2[6][20] ),
    .B2(_09320_),
    .X(_04940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16648_ (.A1(_09267_),
    .A2(_09319_),
    .B1(\design_top.core0.REG2[6][19] ),
    .B2(_09320_),
    .X(_04939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16649_ (.A1(_09268_),
    .A2(_09319_),
    .B1(\design_top.core0.REG2[6][18] ),
    .B2(_09320_),
    .X(_04938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16650_ (.A1(_09269_),
    .A2(_09319_),
    .B1(\design_top.core0.REG2[6][17] ),
    .B2(_09320_),
    .X(_04937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16651_ (.A(_09311_),
    .X(_09321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16652_ (.A(_09314_),
    .X(_09322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16653_ (.A1(_09270_),
    .A2(_09321_),
    .B1(\design_top.core0.REG2[6][16] ),
    .B2(_09322_),
    .X(_04936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16654_ (.A1(_09273_),
    .A2(_09321_),
    .B1(\design_top.core0.REG2[6][15] ),
    .B2(_09322_),
    .X(_04935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16655_ (.A1(_09274_),
    .A2(_09321_),
    .B1(\design_top.core0.REG2[6][14] ),
    .B2(_09322_),
    .X(_04934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16656_ (.A1(\design_top.core0.REG2[6][13] ),
    .A2(_09312_),
    .B1(_09241_),
    .B2(_09315_),
    .X(_04933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16657_ (.A1(_09275_),
    .A2(_09321_),
    .B1(\design_top.core0.REG2[6][12] ),
    .B2(_09322_),
    .X(_04932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16658_ (.A1(_09276_),
    .A2(_09321_),
    .B1(\design_top.core0.REG2[6][11] ),
    .B2(_09322_),
    .X(_04931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16659_ (.A(_09311_),
    .X(_09323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16660_ (.A(_09314_),
    .X(_09324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16661_ (.A1(_09277_),
    .A2(_09323_),
    .B1(\design_top.core0.REG2[6][10] ),
    .B2(_09324_),
    .X(_04930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16662_ (.A1(_09280_),
    .A2(_09323_),
    .B1(\design_top.core0.REG2[6][9] ),
    .B2(_09324_),
    .X(_04929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16663_ (.A1(_09281_),
    .A2(_09323_),
    .B1(\design_top.core0.REG2[6][8] ),
    .B2(_09324_),
    .X(_04928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16664_ (.A1(_09282_),
    .A2(_09323_),
    .B1(\design_top.core0.REG2[6][7] ),
    .B2(_09324_),
    .X(_04927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16665_ (.A1(_09283_),
    .A2(_09323_),
    .B1(\design_top.core0.REG2[6][6] ),
    .B2(_09324_),
    .X(_04926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16666_ (.A(_09311_),
    .X(_09325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16667_ (.A(_09314_),
    .X(_09326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16668_ (.A1(_09284_),
    .A2(_09325_),
    .B1(\design_top.core0.REG2[6][5] ),
    .B2(_09326_),
    .X(_04925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16669_ (.A1(_09287_),
    .A2(_09325_),
    .B1(\design_top.core0.REG2[6][4] ),
    .B2(_09326_),
    .X(_04924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16670_ (.A1(_09288_),
    .A2(_09325_),
    .B1(\design_top.core0.REG2[6][3] ),
    .B2(_09326_),
    .X(_04923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16671_ (.A1(_09289_),
    .A2(_09325_),
    .B1(\design_top.core0.REG2[6][2] ),
    .B2(_09326_),
    .X(_04922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16672_ (.A1(_09290_),
    .A2(_09325_),
    .B1(\design_top.core0.REG2[6][1] ),
    .B2(_09326_),
    .X(_04921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16673_ (.A1(_09291_),
    .A2(_09312_),
    .B1(\design_top.core0.REG2[6][0] ),
    .B2(_09315_),
    .X(_04920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _16674_ (.A(_08778_),
    .B(_08780_),
    .C(_09292_),
    .D(_09086_),
    .X(_09327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16675_ (.A(_09327_),
    .X(_09328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16676_ (.A(_09328_),
    .X(_09329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16677_ (.A(_09329_),
    .X(_09330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16678_ (.A(_09328_),
    .Y(_09331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16679_ (.A(_09331_),
    .X(_09332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16680_ (.A(_09332_),
    .X(_09333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16681_ (.A1(_09244_),
    .A2(_09330_),
    .B1(\design_top.core0.REG2[5][31] ),
    .B2(_09333_),
    .X(_04919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16682_ (.A1(_09252_),
    .A2(_09330_),
    .B1(\design_top.core0.REG2[5][30] ),
    .B2(_09333_),
    .X(_04918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16683_ (.A1(_09253_),
    .A2(_09330_),
    .B1(\design_top.core0.REG2[5][29] ),
    .B2(_09333_),
    .X(_04917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16684_ (.A1(_09254_),
    .A2(_09330_),
    .B1(\design_top.core0.REG2[5][28] ),
    .B2(_09333_),
    .X(_04916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16685_ (.A1(_09255_),
    .A2(_09330_),
    .B1(\design_top.core0.REG2[5][27] ),
    .B2(_09333_),
    .X(_04915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16686_ (.A(_09329_),
    .X(_09334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16687_ (.A(_09332_),
    .X(_09335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16688_ (.A1(_09256_),
    .A2(_09334_),
    .B1(\design_top.core0.REG2[5][26] ),
    .B2(_09335_),
    .X(_04914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16689_ (.A1(_09259_),
    .A2(_09334_),
    .B1(\design_top.core0.REG2[5][25] ),
    .B2(_09335_),
    .X(_04913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16690_ (.A1(_09260_),
    .A2(_09334_),
    .B1(\design_top.core0.REG2[5][24] ),
    .B2(_09335_),
    .X(_04912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16691_ (.A1(_09261_),
    .A2(_09334_),
    .B1(\design_top.core0.REG2[5][23] ),
    .B2(_09335_),
    .X(_04911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16692_ (.A1(_09262_),
    .A2(_09334_),
    .B1(\design_top.core0.REG2[5][22] ),
    .B2(_09335_),
    .X(_04910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16693_ (.A(_09329_),
    .X(_09336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16694_ (.A(_09332_),
    .X(_09337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16695_ (.A1(_09263_),
    .A2(_09336_),
    .B1(\design_top.core0.REG2[5][21] ),
    .B2(_09337_),
    .X(_04909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16696_ (.A1(_09266_),
    .A2(_09336_),
    .B1(\design_top.core0.REG2[5][20] ),
    .B2(_09337_),
    .X(_04908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16697_ (.A1(_09267_),
    .A2(_09336_),
    .B1(\design_top.core0.REG2[5][19] ),
    .B2(_09337_),
    .X(_04907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16698_ (.A1(_09268_),
    .A2(_09336_),
    .B1(\design_top.core0.REG2[5][18] ),
    .B2(_09337_),
    .X(_04906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16699_ (.A1(_09269_),
    .A2(_09336_),
    .B1(\design_top.core0.REG2[5][17] ),
    .B2(_09337_),
    .X(_04905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16700_ (.A(_09328_),
    .X(_09338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16701_ (.A(_09331_),
    .X(_09339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16702_ (.A1(_09270_),
    .A2(_09338_),
    .B1(\design_top.core0.REG2[5][16] ),
    .B2(_09339_),
    .X(_04904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16703_ (.A1(_09273_),
    .A2(_09338_),
    .B1(\design_top.core0.REG2[5][15] ),
    .B2(_09339_),
    .X(_04903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16704_ (.A1(_09274_),
    .A2(_09338_),
    .B1(\design_top.core0.REG2[5][14] ),
    .B2(_09339_),
    .X(_04902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16705_ (.A1(\design_top.core0.REG2[5][13] ),
    .A2(_09329_),
    .B1(_09241_),
    .B2(_09332_),
    .X(_04901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16706_ (.A1(_09275_),
    .A2(_09338_),
    .B1(\design_top.core0.REG2[5][12] ),
    .B2(_09339_),
    .X(_04900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16707_ (.A1(_09276_),
    .A2(_09338_),
    .B1(\design_top.core0.REG2[5][11] ),
    .B2(_09339_),
    .X(_04899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16708_ (.A(_09328_),
    .X(_09340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16709_ (.A(_09331_),
    .X(_09341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16710_ (.A1(_09277_),
    .A2(_09340_),
    .B1(\design_top.core0.REG2[5][10] ),
    .B2(_09341_),
    .X(_04898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16711_ (.A1(_09280_),
    .A2(_09340_),
    .B1(\design_top.core0.REG2[5][9] ),
    .B2(_09341_),
    .X(_04897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16712_ (.A1(_09281_),
    .A2(_09340_),
    .B1(\design_top.core0.REG2[5][8] ),
    .B2(_09341_),
    .X(_04896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16713_ (.A1(_09282_),
    .A2(_09340_),
    .B1(\design_top.core0.REG2[5][7] ),
    .B2(_09341_),
    .X(_04895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16714_ (.A1(_09283_),
    .A2(_09340_),
    .B1(\design_top.core0.REG2[5][6] ),
    .B2(_09341_),
    .X(_04894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16715_ (.A(_09328_),
    .X(_09342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16716_ (.A(_09331_),
    .X(_09343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16717_ (.A1(_09284_),
    .A2(_09342_),
    .B1(\design_top.core0.REG2[5][5] ),
    .B2(_09343_),
    .X(_04893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16718_ (.A1(_09287_),
    .A2(_09342_),
    .B1(\design_top.core0.REG2[5][4] ),
    .B2(_09343_),
    .X(_04892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16719_ (.A1(_09288_),
    .A2(_09342_),
    .B1(\design_top.core0.REG2[5][3] ),
    .B2(_09343_),
    .X(_04891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16720_ (.A1(_09289_),
    .A2(_09342_),
    .B1(\design_top.core0.REG2[5][2] ),
    .B2(_09343_),
    .X(_04890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16721_ (.A1(_09290_),
    .A2(_09342_),
    .B1(\design_top.core0.REG2[5][1] ),
    .B2(_09343_),
    .X(_04889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16722_ (.A1(_09291_),
    .A2(_09329_),
    .B1(\design_top.core0.REG2[5][0] ),
    .B2(_09332_),
    .X(_04888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16723_ (.A1(_08992_),
    .A2(_07867_),
    .B1(_08134_),
    .B2(_09076_),
    .X(_09344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16724_ (.A(_09344_),
    .Y(_09345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16725_ (.A(_09345_),
    .X(_09346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16726_ (.A(_09344_),
    .X(_09347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16727_ (.A1(_00668_),
    .A2(_09346_),
    .B1(\design_top.MEM[7][7] ),
    .B2(_09347_),
    .X(_04887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16728_ (.A1(_00667_),
    .A2(_09346_),
    .B1(\design_top.MEM[7][6] ),
    .B2(_09347_),
    .X(_04886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16729_ (.A1(_00666_),
    .A2(_09346_),
    .B1(\design_top.MEM[7][5] ),
    .B2(_09347_),
    .X(_04885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16730_ (.A1(_00665_),
    .A2(_09346_),
    .B1(\design_top.MEM[7][4] ),
    .B2(_09347_),
    .X(_04884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16731_ (.A1(_00664_),
    .A2(_09346_),
    .B1(\design_top.MEM[7][3] ),
    .B2(_09347_),
    .X(_04883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16732_ (.A1(_00663_),
    .A2(_09345_),
    .B1(\design_top.MEM[7][2] ),
    .B2(_09344_),
    .X(_04882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16733_ (.A1(_00662_),
    .A2(_09345_),
    .B1(\design_top.MEM[7][1] ),
    .B2(_09344_),
    .X(_04881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16734_ (.A1(_00661_),
    .A2(_09345_),
    .B1(\design_top.MEM[7][0] ),
    .B2(_09344_),
    .X(_04880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _16735_ (.A(_08778_),
    .B(_09085_),
    .C(_00863_),
    .D(_09086_),
    .X(_09348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16736_ (.A(_09348_),
    .X(_09349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16737_ (.A(_09349_),
    .X(_09350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16738_ (.A(_09350_),
    .X(_09351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16739_ (.A(_09349_),
    .Y(_09352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16740_ (.A(_09352_),
    .X(_09353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16741_ (.A(_09353_),
    .X(_09354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16742_ (.A1(_09244_),
    .A2(_09351_),
    .B1(\design_top.core0.REG2[4][31] ),
    .B2(_09354_),
    .X(_04879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16743_ (.A1(_09252_),
    .A2(_09351_),
    .B1(\design_top.core0.REG2[4][30] ),
    .B2(_09354_),
    .X(_04878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16744_ (.A1(_09253_),
    .A2(_09351_),
    .B1(\design_top.core0.REG2[4][29] ),
    .B2(_09354_),
    .X(_04877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16745_ (.A1(_09254_),
    .A2(_09351_),
    .B1(\design_top.core0.REG2[4][28] ),
    .B2(_09354_),
    .X(_04876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16746_ (.A1(_09255_),
    .A2(_09351_),
    .B1(\design_top.core0.REG2[4][27] ),
    .B2(_09354_),
    .X(_04875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16747_ (.A(_09350_),
    .X(_09355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16748_ (.A(_09353_),
    .X(_09356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16749_ (.A1(_09256_),
    .A2(_09355_),
    .B1(\design_top.core0.REG2[4][26] ),
    .B2(_09356_),
    .X(_04874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16750_ (.A1(_09259_),
    .A2(_09355_),
    .B1(\design_top.core0.REG2[4][25] ),
    .B2(_09356_),
    .X(_04873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16751_ (.A1(_09260_),
    .A2(_09355_),
    .B1(\design_top.core0.REG2[4][24] ),
    .B2(_09356_),
    .X(_04872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16752_ (.A1(_09261_),
    .A2(_09355_),
    .B1(\design_top.core0.REG2[4][23] ),
    .B2(_09356_),
    .X(_04871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16753_ (.A1(_09262_),
    .A2(_09355_),
    .B1(\design_top.core0.REG2[4][22] ),
    .B2(_09356_),
    .X(_04870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16754_ (.A(_09350_),
    .X(_09357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16755_ (.A(_09353_),
    .X(_09358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16756_ (.A1(_09263_),
    .A2(_09357_),
    .B1(\design_top.core0.REG2[4][21] ),
    .B2(_09358_),
    .X(_04869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16757_ (.A1(_09266_),
    .A2(_09357_),
    .B1(\design_top.core0.REG2[4][20] ),
    .B2(_09358_),
    .X(_04868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16758_ (.A1(_09267_),
    .A2(_09357_),
    .B1(\design_top.core0.REG2[4][19] ),
    .B2(_09358_),
    .X(_04867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16759_ (.A1(_09268_),
    .A2(_09357_),
    .B1(\design_top.core0.REG2[4][18] ),
    .B2(_09358_),
    .X(_04866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16760_ (.A1(_09269_),
    .A2(_09357_),
    .B1(\design_top.core0.REG2[4][17] ),
    .B2(_09358_),
    .X(_04865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16761_ (.A(_09349_),
    .X(_09359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16762_ (.A(_09352_),
    .X(_09360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16763_ (.A1(_09270_),
    .A2(_09359_),
    .B1(\design_top.core0.REG2[4][16] ),
    .B2(_09360_),
    .X(_04864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16764_ (.A1(_09273_),
    .A2(_09359_),
    .B1(\design_top.core0.REG2[4][15] ),
    .B2(_09360_),
    .X(_04863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16765_ (.A1(_09274_),
    .A2(_09359_),
    .B1(\design_top.core0.REG2[4][14] ),
    .B2(_09360_),
    .X(_04862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16766_ (.A(_08844_),
    .X(_09361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16767_ (.A1(\design_top.core0.REG2[4][13] ),
    .A2(_09350_),
    .B1(_09361_),
    .B2(_09353_),
    .X(_04861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16768_ (.A1(_09275_),
    .A2(_09359_),
    .B1(\design_top.core0.REG2[4][12] ),
    .B2(_09360_),
    .X(_04860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16769_ (.A1(_09276_),
    .A2(_09359_),
    .B1(\design_top.core0.REG2[4][11] ),
    .B2(_09360_),
    .X(_04859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16770_ (.A(_09349_),
    .X(_09362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16771_ (.A(_09352_),
    .X(_09363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16772_ (.A1(_09277_),
    .A2(_09362_),
    .B1(\design_top.core0.REG2[4][10] ),
    .B2(_09363_),
    .X(_04858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16773_ (.A1(_09280_),
    .A2(_09362_),
    .B1(\design_top.core0.REG2[4][9] ),
    .B2(_09363_),
    .X(_04857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16774_ (.A1(_09281_),
    .A2(_09362_),
    .B1(\design_top.core0.REG2[4][8] ),
    .B2(_09363_),
    .X(_04856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16775_ (.A1(_09282_),
    .A2(_09362_),
    .B1(\design_top.core0.REG2[4][7] ),
    .B2(_09363_),
    .X(_04855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16776_ (.A1(_09283_),
    .A2(_09362_),
    .B1(\design_top.core0.REG2[4][6] ),
    .B2(_09363_),
    .X(_04854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16777_ (.A(_09349_),
    .X(_09364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16778_ (.A(_09352_),
    .X(_09365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16779_ (.A1(_09284_),
    .A2(_09364_),
    .B1(\design_top.core0.REG2[4][5] ),
    .B2(_09365_),
    .X(_04853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16780_ (.A1(_09287_),
    .A2(_09364_),
    .B1(\design_top.core0.REG2[4][4] ),
    .B2(_09365_),
    .X(_04852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16781_ (.A1(_09288_),
    .A2(_09364_),
    .B1(\design_top.core0.REG2[4][3] ),
    .B2(_09365_),
    .X(_04851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16782_ (.A1(_09289_),
    .A2(_09364_),
    .B1(\design_top.core0.REG2[4][2] ),
    .B2(_09365_),
    .X(_04850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16783_ (.A1(_09290_),
    .A2(_09364_),
    .B1(\design_top.core0.REG2[4][1] ),
    .B2(_09365_),
    .X(_04849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16784_ (.A1(_09291_),
    .A2(_09350_),
    .B1(\design_top.core0.REG2[4][0] ),
    .B2(_09353_),
    .X(_04848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16785_ (.A(_09081_),
    .X(_09366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _16786_ (.A(_09292_),
    .B(_09200_),
    .C(_09083_),
    .D(_08779_),
    .X(_09367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16787_ (.A(_09367_),
    .X(_09368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16788_ (.A(_09368_),
    .X(_09369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16789_ (.A(_09369_),
    .X(_09370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16790_ (.A(_09368_),
    .Y(_09371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16791_ (.A(_09371_),
    .X(_09372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16792_ (.A(_09372_),
    .X(_09373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16793_ (.A1(_09366_),
    .A2(_09370_),
    .B1(\design_top.core0.REG2[3][31] ),
    .B2(_09373_),
    .X(_04847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16794_ (.A(_09095_),
    .X(_09374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16795_ (.A1(_09374_),
    .A2(_09370_),
    .B1(\design_top.core0.REG2[3][30] ),
    .B2(_09373_),
    .X(_04846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16796_ (.A(_09097_),
    .X(_09375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16797_ (.A1(_09375_),
    .A2(_09370_),
    .B1(\design_top.core0.REG2[3][29] ),
    .B2(_09373_),
    .X(_04845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16798_ (.A(_09099_),
    .X(_09376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16799_ (.A1(_09376_),
    .A2(_09370_),
    .B1(\design_top.core0.REG2[3][28] ),
    .B2(_09373_),
    .X(_04844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16800_ (.A(_09101_),
    .X(_09377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16801_ (.A1(_09377_),
    .A2(_09370_),
    .B1(\design_top.core0.REG2[3][27] ),
    .B2(_09373_),
    .X(_04843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16802_ (.A(_09103_),
    .X(_09378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16803_ (.A(_09369_),
    .X(_09379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16804_ (.A(_09372_),
    .X(_09380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16805_ (.A1(_09378_),
    .A2(_09379_),
    .B1(\design_top.core0.REG2[3][26] ),
    .B2(_09380_),
    .X(_04842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16806_ (.A(_09107_),
    .X(_09381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16807_ (.A1(_09381_),
    .A2(_09379_),
    .B1(\design_top.core0.REG2[3][25] ),
    .B2(_09380_),
    .X(_04841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16808_ (.A(_09109_),
    .X(_09382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16809_ (.A1(_09382_),
    .A2(_09379_),
    .B1(\design_top.core0.REG2[3][24] ),
    .B2(_09380_),
    .X(_04840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16810_ (.A(_09111_),
    .X(_09383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16811_ (.A1(_09383_),
    .A2(_09379_),
    .B1(\design_top.core0.REG2[3][23] ),
    .B2(_09380_),
    .X(_04839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16812_ (.A(_09113_),
    .X(_09384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16813_ (.A1(_09384_),
    .A2(_09379_),
    .B1(\design_top.core0.REG2[3][22] ),
    .B2(_09380_),
    .X(_04838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16814_ (.A(_09115_),
    .X(_09385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16815_ (.A(_09369_),
    .X(_09386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16816_ (.A(_09372_),
    .X(_09387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16817_ (.A1(_09385_),
    .A2(_09386_),
    .B1(\design_top.core0.REG2[3][21] ),
    .B2(_09387_),
    .X(_04837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16818_ (.A(_09119_),
    .X(_09388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16819_ (.A1(_09388_),
    .A2(_09386_),
    .B1(\design_top.core0.REG2[3][20] ),
    .B2(_09387_),
    .X(_04836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16820_ (.A(_09121_),
    .X(_09389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16821_ (.A1(_09389_),
    .A2(_09386_),
    .B1(\design_top.core0.REG2[3][19] ),
    .B2(_09387_),
    .X(_04835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16822_ (.A(_09123_),
    .X(_09390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16823_ (.A1(_09390_),
    .A2(_09386_),
    .B1(\design_top.core0.REG2[3][18] ),
    .B2(_09387_),
    .X(_04834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16824_ (.A(_09125_),
    .X(_09391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16825_ (.A1(_09391_),
    .A2(_09386_),
    .B1(\design_top.core0.REG2[3][17] ),
    .B2(_09387_),
    .X(_04833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16826_ (.A(_09127_),
    .X(_09392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16827_ (.A(_09368_),
    .X(_09393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16828_ (.A(_09371_),
    .X(_09394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16829_ (.A1(_09392_),
    .A2(_09393_),
    .B1(\design_top.core0.REG2[3][16] ),
    .B2(_09394_),
    .X(_04832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16830_ (.A(_09131_),
    .X(_09395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16831_ (.A1(_09395_),
    .A2(_09393_),
    .B1(\design_top.core0.REG2[3][15] ),
    .B2(_09394_),
    .X(_04831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16832_ (.A(_09133_),
    .X(_09396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16833_ (.A1(_09396_),
    .A2(_09393_),
    .B1(\design_top.core0.REG2[3][14] ),
    .B2(_09394_),
    .X(_04830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16834_ (.A1(\design_top.core0.REG2[3][13] ),
    .A2(_09369_),
    .B1(_09361_),
    .B2(_09372_),
    .X(_04829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16835_ (.A(_09136_),
    .X(_09397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16836_ (.A1(_09397_),
    .A2(_09393_),
    .B1(\design_top.core0.REG2[3][12] ),
    .B2(_09394_),
    .X(_04828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16837_ (.A(_09138_),
    .X(_09398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16838_ (.A1(_09398_),
    .A2(_09393_),
    .B1(\design_top.core0.REG2[3][11] ),
    .B2(_09394_),
    .X(_04827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16839_ (.A(_09140_),
    .X(_09399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16840_ (.A(_09368_),
    .X(_09400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16841_ (.A(_09371_),
    .X(_09401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16842_ (.A1(_09399_),
    .A2(_09400_),
    .B1(\design_top.core0.REG2[3][10] ),
    .B2(_09401_),
    .X(_04826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16843_ (.A(_09144_),
    .X(_09402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16844_ (.A1(_09402_),
    .A2(_09400_),
    .B1(\design_top.core0.REG2[3][9] ),
    .B2(_09401_),
    .X(_04825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16845_ (.A(_09146_),
    .X(_09403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16846_ (.A1(_09403_),
    .A2(_09400_),
    .B1(\design_top.core0.REG2[3][8] ),
    .B2(_09401_),
    .X(_04824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16847_ (.A(_09148_),
    .X(_09404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16848_ (.A1(_09404_),
    .A2(_09400_),
    .B1(\design_top.core0.REG2[3][7] ),
    .B2(_09401_),
    .X(_04823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16849_ (.A(_09150_),
    .X(_09405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16850_ (.A1(_09405_),
    .A2(_09400_),
    .B1(\design_top.core0.REG2[3][6] ),
    .B2(_09401_),
    .X(_04822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16851_ (.A(_09152_),
    .X(_09406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16852_ (.A(_09368_),
    .X(_09407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16853_ (.A(_09371_),
    .X(_09408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16854_ (.A1(_09406_),
    .A2(_09407_),
    .B1(\design_top.core0.REG2[3][5] ),
    .B2(_09408_),
    .X(_04821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16855_ (.A(_09156_),
    .X(_09409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16856_ (.A1(_09409_),
    .A2(_09407_),
    .B1(\design_top.core0.REG2[3][4] ),
    .B2(_09408_),
    .X(_04820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16857_ (.A(_09158_),
    .X(_09410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16858_ (.A1(_09410_),
    .A2(_09407_),
    .B1(\design_top.core0.REG2[3][3] ),
    .B2(_09408_),
    .X(_04819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16859_ (.A(_09160_),
    .X(_09411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16860_ (.A1(_09411_),
    .A2(_09407_),
    .B1(\design_top.core0.REG2[3][2] ),
    .B2(_09408_),
    .X(_04818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16861_ (.A(_09162_),
    .X(_09412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16862_ (.A1(_09412_),
    .A2(_09407_),
    .B1(\design_top.core0.REG2[3][1] ),
    .B2(_09408_),
    .X(_04817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16863_ (.A(_09164_),
    .X(_09413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16864_ (.A1(_09413_),
    .A2(_09369_),
    .B1(\design_top.core0.REG2[3][0] ),
    .B2(_09372_),
    .X(_04816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _16865_ (.A(_09292_),
    .B(_09200_),
    .C(_09083_),
    .D(_00860_),
    .X(_09414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16866_ (.A(_09414_),
    .X(_09415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16867_ (.A(_09415_),
    .X(_09416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16868_ (.A(_09416_),
    .X(_09417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16869_ (.A(_09415_),
    .Y(_09418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16870_ (.A(_09418_),
    .X(_09419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16871_ (.A(_09419_),
    .X(_09420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16872_ (.A1(_09366_),
    .A2(_09417_),
    .B1(\design_top.core0.REG2[2][31] ),
    .B2(_09420_),
    .X(_04815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16873_ (.A1(_09374_),
    .A2(_09417_),
    .B1(\design_top.core0.REG2[2][30] ),
    .B2(_09420_),
    .X(_04814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16874_ (.A1(_09375_),
    .A2(_09417_),
    .B1(\design_top.core0.REG2[2][29] ),
    .B2(_09420_),
    .X(_04813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16875_ (.A1(_09376_),
    .A2(_09417_),
    .B1(\design_top.core0.REG2[2][28] ),
    .B2(_09420_),
    .X(_04812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16876_ (.A1(_09377_),
    .A2(_09417_),
    .B1(\design_top.core0.REG2[2][27] ),
    .B2(_09420_),
    .X(_04811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16877_ (.A(_09416_),
    .X(_09421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16878_ (.A(_09419_),
    .X(_09422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16879_ (.A1(_09378_),
    .A2(_09421_),
    .B1(\design_top.core0.REG2[2][26] ),
    .B2(_09422_),
    .X(_04810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16880_ (.A1(_09381_),
    .A2(_09421_),
    .B1(\design_top.core0.REG2[2][25] ),
    .B2(_09422_),
    .X(_04809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16881_ (.A1(_09382_),
    .A2(_09421_),
    .B1(\design_top.core0.REG2[2][24] ),
    .B2(_09422_),
    .X(_04808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16882_ (.A1(_09383_),
    .A2(_09421_),
    .B1(\design_top.core0.REG2[2][23] ),
    .B2(_09422_),
    .X(_04807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16883_ (.A1(_09384_),
    .A2(_09421_),
    .B1(\design_top.core0.REG2[2][22] ),
    .B2(_09422_),
    .X(_04806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16884_ (.A(_09416_),
    .X(_09423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16885_ (.A(_09419_),
    .X(_09424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16886_ (.A1(_09385_),
    .A2(_09423_),
    .B1(\design_top.core0.REG2[2][21] ),
    .B2(_09424_),
    .X(_04805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16887_ (.A1(_09388_),
    .A2(_09423_),
    .B1(\design_top.core0.REG2[2][20] ),
    .B2(_09424_),
    .X(_04804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16888_ (.A1(_09389_),
    .A2(_09423_),
    .B1(\design_top.core0.REG2[2][19] ),
    .B2(_09424_),
    .X(_04803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16889_ (.A1(_09390_),
    .A2(_09423_),
    .B1(\design_top.core0.REG2[2][18] ),
    .B2(_09424_),
    .X(_04802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16890_ (.A1(_09391_),
    .A2(_09423_),
    .B1(\design_top.core0.REG2[2][17] ),
    .B2(_09424_),
    .X(_04801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16891_ (.A(_09415_),
    .X(_09425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16892_ (.A(_09418_),
    .X(_09426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16893_ (.A1(_09392_),
    .A2(_09425_),
    .B1(\design_top.core0.REG2[2][16] ),
    .B2(_09426_),
    .X(_04800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16894_ (.A1(_09395_),
    .A2(_09425_),
    .B1(\design_top.core0.REG2[2][15] ),
    .B2(_09426_),
    .X(_04799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16895_ (.A1(_09396_),
    .A2(_09425_),
    .B1(\design_top.core0.REG2[2][14] ),
    .B2(_09426_),
    .X(_04798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16896_ (.A1(\design_top.core0.REG2[2][13] ),
    .A2(_09416_),
    .B1(_09361_),
    .B2(_09419_),
    .X(_04797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16897_ (.A1(_09397_),
    .A2(_09425_),
    .B1(\design_top.core0.REG2[2][12] ),
    .B2(_09426_),
    .X(_04796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16898_ (.A1(_09398_),
    .A2(_09425_),
    .B1(\design_top.core0.REG2[2][11] ),
    .B2(_09426_),
    .X(_04795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16899_ (.A(_09415_),
    .X(_09427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16900_ (.A(_09418_),
    .X(_09428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16901_ (.A1(_09399_),
    .A2(_09427_),
    .B1(\design_top.core0.REG2[2][10] ),
    .B2(_09428_),
    .X(_04794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16902_ (.A1(_09402_),
    .A2(_09427_),
    .B1(\design_top.core0.REG2[2][9] ),
    .B2(_09428_),
    .X(_04793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16903_ (.A1(_09403_),
    .A2(_09427_),
    .B1(\design_top.core0.REG2[2][8] ),
    .B2(_09428_),
    .X(_04792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16904_ (.A1(_09404_),
    .A2(_09427_),
    .B1(\design_top.core0.REG2[2][7] ),
    .B2(_09428_),
    .X(_04791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16905_ (.A1(_09405_),
    .A2(_09427_),
    .B1(\design_top.core0.REG2[2][6] ),
    .B2(_09428_),
    .X(_04790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16906_ (.A(_09415_),
    .X(_09429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16907_ (.A(_09418_),
    .X(_09430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16908_ (.A1(_09406_),
    .A2(_09429_),
    .B1(\design_top.core0.REG2[2][5] ),
    .B2(_09430_),
    .X(_04789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16909_ (.A1(_09409_),
    .A2(_09429_),
    .B1(\design_top.core0.REG2[2][4] ),
    .B2(_09430_),
    .X(_04788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16910_ (.A1(_09410_),
    .A2(_09429_),
    .B1(\design_top.core0.REG2[2][3] ),
    .B2(_09430_),
    .X(_04787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16911_ (.A1(_09411_),
    .A2(_09429_),
    .B1(\design_top.core0.REG2[2][2] ),
    .B2(_09430_),
    .X(_04786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16912_ (.A1(_09412_),
    .A2(_09429_),
    .B1(\design_top.core0.REG2[2][1] ),
    .B2(_09430_),
    .X(_04785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16913_ (.A1(_09413_),
    .A2(_09416_),
    .B1(\design_top.core0.REG2[2][0] ),
    .B2(_09419_),
    .X(_04784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _16914_ (.A(_00861_),
    .B(_08780_),
    .C(_00863_),
    .D(_00862_),
    .X(_09431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16915_ (.A(_09431_),
    .X(_09432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16916_ (.A(_09432_),
    .X(_09433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16917_ (.A(_09433_),
    .X(_09434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16918_ (.A(_09432_),
    .Y(_09435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16919_ (.A(_09435_),
    .X(_09436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16920_ (.A(_09436_),
    .X(_09437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16921_ (.A1(_09366_),
    .A2(_09434_),
    .B1(\design_top.core0.REG2[1][31] ),
    .B2(_09437_),
    .X(_04783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16922_ (.A1(_09374_),
    .A2(_09434_),
    .B1(\design_top.core0.REG2[1][30] ),
    .B2(_09437_),
    .X(_04782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16923_ (.A1(_09375_),
    .A2(_09434_),
    .B1(\design_top.core0.REG2[1][29] ),
    .B2(_09437_),
    .X(_04781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16924_ (.A1(_09376_),
    .A2(_09434_),
    .B1(\design_top.core0.REG2[1][28] ),
    .B2(_09437_),
    .X(_04780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16925_ (.A1(_09377_),
    .A2(_09434_),
    .B1(\design_top.core0.REG2[1][27] ),
    .B2(_09437_),
    .X(_04779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16926_ (.A(_09433_),
    .X(_09438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16927_ (.A(_09436_),
    .X(_09439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16928_ (.A1(_09378_),
    .A2(_09438_),
    .B1(\design_top.core0.REG2[1][26] ),
    .B2(_09439_),
    .X(_04778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16929_ (.A1(_09381_),
    .A2(_09438_),
    .B1(\design_top.core0.REG2[1][25] ),
    .B2(_09439_),
    .X(_04777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16930_ (.A1(_09382_),
    .A2(_09438_),
    .B1(\design_top.core0.REG2[1][24] ),
    .B2(_09439_),
    .X(_04776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16931_ (.A1(_09383_),
    .A2(_09438_),
    .B1(\design_top.core0.REG2[1][23] ),
    .B2(_09439_),
    .X(_04775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16932_ (.A1(_09384_),
    .A2(_09438_),
    .B1(\design_top.core0.REG2[1][22] ),
    .B2(_09439_),
    .X(_04774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16933_ (.A(_09433_),
    .X(_09440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16934_ (.A(_09436_),
    .X(_09441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16935_ (.A1(_09385_),
    .A2(_09440_),
    .B1(\design_top.core0.REG2[1][21] ),
    .B2(_09441_),
    .X(_04773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16936_ (.A1(_09388_),
    .A2(_09440_),
    .B1(\design_top.core0.REG2[1][20] ),
    .B2(_09441_),
    .X(_04772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16937_ (.A1(_09389_),
    .A2(_09440_),
    .B1(\design_top.core0.REG2[1][19] ),
    .B2(_09441_),
    .X(_04771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16938_ (.A1(_09390_),
    .A2(_09440_),
    .B1(\design_top.core0.REG2[1][18] ),
    .B2(_09441_),
    .X(_04770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16939_ (.A1(_09391_),
    .A2(_09440_),
    .B1(\design_top.core0.REG2[1][17] ),
    .B2(_09441_),
    .X(_04769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16940_ (.A(_09432_),
    .X(_09442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16941_ (.A(_09435_),
    .X(_09443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16942_ (.A1(_09392_),
    .A2(_09442_),
    .B1(\design_top.core0.REG2[1][16] ),
    .B2(_09443_),
    .X(_04768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16943_ (.A1(_09395_),
    .A2(_09442_),
    .B1(\design_top.core0.REG2[1][15] ),
    .B2(_09443_),
    .X(_04767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16944_ (.A1(_09396_),
    .A2(_09442_),
    .B1(\design_top.core0.REG2[1][14] ),
    .B2(_09443_),
    .X(_04766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16945_ (.A1(\design_top.core0.REG2[1][13] ),
    .A2(_09433_),
    .B1(_09361_),
    .B2(_09436_),
    .X(_04765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16946_ (.A1(_09397_),
    .A2(_09442_),
    .B1(\design_top.core0.REG2[1][12] ),
    .B2(_09443_),
    .X(_04764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16947_ (.A1(_09398_),
    .A2(_09442_),
    .B1(\design_top.core0.REG2[1][11] ),
    .B2(_09443_),
    .X(_04763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16948_ (.A(_09432_),
    .X(_09444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16949_ (.A(_09435_),
    .X(_09445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16950_ (.A1(_09399_),
    .A2(_09444_),
    .B1(\design_top.core0.REG2[1][10] ),
    .B2(_09445_),
    .X(_04762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16951_ (.A1(_09402_),
    .A2(_09444_),
    .B1(\design_top.core0.REG2[1][9] ),
    .B2(_09445_),
    .X(_04761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16952_ (.A1(_09403_),
    .A2(_09444_),
    .B1(\design_top.core0.REG2[1][8] ),
    .B2(_09445_),
    .X(_04760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16953_ (.A1(_09404_),
    .A2(_09444_),
    .B1(\design_top.core0.REG2[1][7] ),
    .B2(_09445_),
    .X(_04759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16954_ (.A1(_09405_),
    .A2(_09444_),
    .B1(\design_top.core0.REG2[1][6] ),
    .B2(_09445_),
    .X(_04758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16955_ (.A(_09432_),
    .X(_09446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16956_ (.A(_09435_),
    .X(_09447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16957_ (.A1(_09406_),
    .A2(_09446_),
    .B1(\design_top.core0.REG2[1][5] ),
    .B2(_09447_),
    .X(_04757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16958_ (.A1(_09409_),
    .A2(_09446_),
    .B1(\design_top.core0.REG2[1][4] ),
    .B2(_09447_),
    .X(_04756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16959_ (.A1(_09410_),
    .A2(_09446_),
    .B1(\design_top.core0.REG2[1][3] ),
    .B2(_09447_),
    .X(_04755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16960_ (.A1(_09411_),
    .A2(_09446_),
    .B1(\design_top.core0.REG2[1][2] ),
    .B2(_09447_),
    .X(_04754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16961_ (.A1(_09412_),
    .A2(_09446_),
    .B1(\design_top.core0.REG2[1][1] ),
    .B2(_09447_),
    .X(_04753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16962_ (.A1(_09413_),
    .A2(_09433_),
    .B1(\design_top.core0.REG2[1][0] ),
    .B2(_09436_),
    .X(_04752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _16963_ (.A(_08782_),
    .B(_09087_),
    .C(_09083_),
    .D(_08779_),
    .X(_09448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16964_ (.A(_09448_),
    .X(_09449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16965_ (.A(_09449_),
    .X(_09450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16966_ (.A(_09450_),
    .X(_09451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _16967_ (.A(_09449_),
    .Y(_09452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16968_ (.A(_09452_),
    .X(_09453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16969_ (.A(_09453_),
    .X(_09454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16970_ (.A1(_09366_),
    .A2(_09451_),
    .B1(\design_top.core0.REG2[15][31] ),
    .B2(_09454_),
    .X(_04751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16971_ (.A1(_09374_),
    .A2(_09451_),
    .B1(\design_top.core0.REG2[15][30] ),
    .B2(_09454_),
    .X(_04750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16972_ (.A1(_09375_),
    .A2(_09451_),
    .B1(\design_top.core0.REG2[15][29] ),
    .B2(_09454_),
    .X(_04749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16973_ (.A1(_09376_),
    .A2(_09451_),
    .B1(\design_top.core0.REG2[15][28] ),
    .B2(_09454_),
    .X(_04748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16974_ (.A1(_09377_),
    .A2(_09451_),
    .B1(\design_top.core0.REG2[15][27] ),
    .B2(_09454_),
    .X(_04747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16975_ (.A(_09450_),
    .X(_09455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16976_ (.A(_09453_),
    .X(_09456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16977_ (.A1(_09378_),
    .A2(_09455_),
    .B1(\design_top.core0.REG2[15][26] ),
    .B2(_09456_),
    .X(_04746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16978_ (.A1(_09381_),
    .A2(_09455_),
    .B1(\design_top.core0.REG2[15][25] ),
    .B2(_09456_),
    .X(_04745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16979_ (.A1(_09382_),
    .A2(_09455_),
    .B1(\design_top.core0.REG2[15][24] ),
    .B2(_09456_),
    .X(_04744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16980_ (.A1(_09383_),
    .A2(_09455_),
    .B1(\design_top.core0.REG2[15][23] ),
    .B2(_09456_),
    .X(_04743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16981_ (.A1(_09384_),
    .A2(_09455_),
    .B1(\design_top.core0.REG2[15][22] ),
    .B2(_09456_),
    .X(_04742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16982_ (.A(_09450_),
    .X(_09457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16983_ (.A(_09453_),
    .X(_09458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16984_ (.A1(_09385_),
    .A2(_09457_),
    .B1(\design_top.core0.REG2[15][21] ),
    .B2(_09458_),
    .X(_04741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16985_ (.A1(_09388_),
    .A2(_09457_),
    .B1(\design_top.core0.REG2[15][20] ),
    .B2(_09458_),
    .X(_04740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16986_ (.A1(_09389_),
    .A2(_09457_),
    .B1(\design_top.core0.REG2[15][19] ),
    .B2(_09458_),
    .X(_04739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16987_ (.A1(_09390_),
    .A2(_09457_),
    .B1(\design_top.core0.REG2[15][18] ),
    .B2(_09458_),
    .X(_04738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16988_ (.A1(_09391_),
    .A2(_09457_),
    .B1(\design_top.core0.REG2[15][17] ),
    .B2(_09458_),
    .X(_04737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16989_ (.A(_09449_),
    .X(_09459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16990_ (.A(_09452_),
    .X(_09460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16991_ (.A1(_09392_),
    .A2(_09459_),
    .B1(\design_top.core0.REG2[15][16] ),
    .B2(_09460_),
    .X(_04736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16992_ (.A1(_09395_),
    .A2(_09459_),
    .B1(\design_top.core0.REG2[15][15] ),
    .B2(_09460_),
    .X(_04735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16993_ (.A1(_09396_),
    .A2(_09459_),
    .B1(\design_top.core0.REG2[15][14] ),
    .B2(_09460_),
    .X(_04734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _16994_ (.A1(\design_top.core0.REG2[15][13] ),
    .A2(_09450_),
    .B1(_09361_),
    .B2(_09453_),
    .X(_04733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16995_ (.A1(_09397_),
    .A2(_09459_),
    .B1(\design_top.core0.REG2[15][12] ),
    .B2(_09460_),
    .X(_04732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16996_ (.A1(_09398_),
    .A2(_09459_),
    .B1(\design_top.core0.REG2[15][11] ),
    .B2(_09460_),
    .X(_04731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16997_ (.A(_09449_),
    .X(_09461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _16998_ (.A(_09452_),
    .X(_09462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _16999_ (.A1(_09399_),
    .A2(_09461_),
    .B1(\design_top.core0.REG2[15][10] ),
    .B2(_09462_),
    .X(_04730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17000_ (.A1(_09402_),
    .A2(_09461_),
    .B1(\design_top.core0.REG2[15][9] ),
    .B2(_09462_),
    .X(_04729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17001_ (.A1(_09403_),
    .A2(_09461_),
    .B1(\design_top.core0.REG2[15][8] ),
    .B2(_09462_),
    .X(_04728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17002_ (.A1(_09404_),
    .A2(_09461_),
    .B1(\design_top.core0.REG2[15][7] ),
    .B2(_09462_),
    .X(_04727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17003_ (.A1(_09405_),
    .A2(_09461_),
    .B1(\design_top.core0.REG2[15][6] ),
    .B2(_09462_),
    .X(_04726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17004_ (.A(_09449_),
    .X(_09463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17005_ (.A(_09452_),
    .X(_09464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17006_ (.A1(_09406_),
    .A2(_09463_),
    .B1(\design_top.core0.REG2[15][5] ),
    .B2(_09464_),
    .X(_04725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17007_ (.A1(_09409_),
    .A2(_09463_),
    .B1(\design_top.core0.REG2[15][4] ),
    .B2(_09464_),
    .X(_04724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17008_ (.A1(_09410_),
    .A2(_09463_),
    .B1(\design_top.core0.REG2[15][3] ),
    .B2(_09464_),
    .X(_04723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17009_ (.A1(_09411_),
    .A2(_09463_),
    .B1(\design_top.core0.REG2[15][2] ),
    .B2(_09464_),
    .X(_04722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17010_ (.A1(_09412_),
    .A2(_09463_),
    .B1(\design_top.core0.REG2[15][1] ),
    .B2(_09464_),
    .X(_04721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17011_ (.A1(_09413_),
    .A2(_09450_),
    .B1(\design_top.core0.REG2[15][0] ),
    .B2(_09453_),
    .X(_04720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17012_ (.A1(_09032_),
    .A2(_07867_),
    .B1(_08150_),
    .B2(_09076_),
    .X(_09465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17013_ (.A(_09465_),
    .Y(_09466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17014_ (.A(_09466_),
    .X(_09467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17015_ (.A(_09465_),
    .X(_09468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17016_ (.A1(_00660_),
    .A2(_09467_),
    .B1(\design_top.MEM[6][7] ),
    .B2(_09468_),
    .X(_04719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17017_ (.A1(_00659_),
    .A2(_09467_),
    .B1(\design_top.MEM[6][6] ),
    .B2(_09468_),
    .X(_04718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17018_ (.A1(_00658_),
    .A2(_09467_),
    .B1(\design_top.MEM[6][5] ),
    .B2(_09468_),
    .X(_04717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17019_ (.A1(_00657_),
    .A2(_09467_),
    .B1(\design_top.MEM[6][4] ),
    .B2(_09468_),
    .X(_04716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17020_ (.A1(_00656_),
    .A2(_09467_),
    .B1(\design_top.MEM[6][3] ),
    .B2(_09468_),
    .X(_04715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17021_ (.A1(_00655_),
    .A2(_09466_),
    .B1(\design_top.MEM[6][2] ),
    .B2(_09465_),
    .X(_04714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17022_ (.A1(_00654_),
    .A2(_09466_),
    .B1(\design_top.MEM[6][1] ),
    .B2(_09465_),
    .X(_04713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17023_ (.A1(_00653_),
    .A2(_09466_),
    .B1(\design_top.MEM[6][0] ),
    .B2(_09465_),
    .X(_04712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17024_ (.A1(_08992_),
    .A2(_08170_),
    .B1(_08166_),
    .B2(_09076_),
    .X(_09469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17025_ (.A(_09469_),
    .Y(_09470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17026_ (.A(_09470_),
    .X(_09471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17027_ (.A(_09469_),
    .X(_09472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17028_ (.A1(_00652_),
    .A2(_09471_),
    .B1(\design_top.MEM[63][7] ),
    .B2(_09472_),
    .X(_04711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17029_ (.A1(_00651_),
    .A2(_09471_),
    .B1(\design_top.MEM[63][6] ),
    .B2(_09472_),
    .X(_04710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17030_ (.A1(_00650_),
    .A2(_09471_),
    .B1(\design_top.MEM[63][5] ),
    .B2(_09472_),
    .X(_04709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17031_ (.A1(_00649_),
    .A2(_09471_),
    .B1(\design_top.MEM[63][4] ),
    .B2(_09472_),
    .X(_04708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17032_ (.A1(_00648_),
    .A2(_09471_),
    .B1(\design_top.MEM[63][3] ),
    .B2(_09472_),
    .X(_04707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17033_ (.A1(_00647_),
    .A2(_09470_),
    .B1(\design_top.MEM[63][2] ),
    .B2(_09469_),
    .X(_04706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17034_ (.A1(_00646_),
    .A2(_09470_),
    .B1(\design_top.MEM[63][1] ),
    .B2(_09469_),
    .X(_04705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17035_ (.A1(_00645_),
    .A2(_09470_),
    .B1(\design_top.MEM[63][0] ),
    .B2(_09469_),
    .X(_04704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17036_ (.A1(_09032_),
    .A2(_08169_),
    .B1(_08193_),
    .B2(_09076_),
    .X(_09473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17037_ (.A(_09473_),
    .Y(_09474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17038_ (.A(_09474_),
    .X(_09475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17039_ (.A(_09473_),
    .X(_09476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17040_ (.A1(_00644_),
    .A2(_09475_),
    .B1(\design_top.MEM[62][7] ),
    .B2(_09476_),
    .X(_04703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17041_ (.A1(_00643_),
    .A2(_09475_),
    .B1(\design_top.MEM[62][6] ),
    .B2(_09476_),
    .X(_04702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17042_ (.A1(_00642_),
    .A2(_09475_),
    .B1(\design_top.MEM[62][5] ),
    .B2(_09476_),
    .X(_04701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17043_ (.A1(_00641_),
    .A2(_09475_),
    .B1(\design_top.MEM[62][4] ),
    .B2(_09476_),
    .X(_04700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17044_ (.A1(_00640_),
    .A2(_09475_),
    .B1(\design_top.MEM[62][3] ),
    .B2(_09476_),
    .X(_04699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17045_ (.A1(_00639_),
    .A2(_09474_),
    .B1(\design_top.MEM[62][2] ),
    .B2(_09473_),
    .X(_04698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17046_ (.A1(_00638_),
    .A2(_09474_),
    .B1(\design_top.MEM[62][1] ),
    .B2(_09473_),
    .X(_04697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17047_ (.A1(_00637_),
    .A2(_09474_),
    .B1(\design_top.MEM[62][0] ),
    .B2(_09473_),
    .X(_04696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17048_ (.A(_08789_),
    .X(_09477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _17049_ (.A(_09477_),
    .B(_09088_),
    .X(_09478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17050_ (.A(_09478_),
    .X(_09479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17051_ (.A(_09479_),
    .X(_09480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17052_ (.A(_09478_),
    .Y(_09481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17053_ (.A(_09481_),
    .X(_09482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17054_ (.A(_09482_),
    .X(_09483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17055_ (.A1(_09366_),
    .A2(_09480_),
    .B1(\design_top.core0.REG1[14][31] ),
    .B2(_09483_),
    .X(_04695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17056_ (.A1(_09374_),
    .A2(_09480_),
    .B1(\design_top.core0.REG1[14][30] ),
    .B2(_09483_),
    .X(_04694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17057_ (.A1(_09375_),
    .A2(_09480_),
    .B1(\design_top.core0.REG1[14][29] ),
    .B2(_09483_),
    .X(_04693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17058_ (.A1(_09376_),
    .A2(_09480_),
    .B1(\design_top.core0.REG1[14][28] ),
    .B2(_09483_),
    .X(_04692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17059_ (.A1(_09377_),
    .A2(_09480_),
    .B1(\design_top.core0.REG1[14][27] ),
    .B2(_09483_),
    .X(_04691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17060_ (.A(_09479_),
    .X(_09484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17061_ (.A(_09482_),
    .X(_09485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17062_ (.A1(_09378_),
    .A2(_09484_),
    .B1(\design_top.core0.REG1[14][26] ),
    .B2(_09485_),
    .X(_04690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17063_ (.A1(_09381_),
    .A2(_09484_),
    .B1(\design_top.core0.REG1[14][25] ),
    .B2(_09485_),
    .X(_04689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17064_ (.A1(_09382_),
    .A2(_09484_),
    .B1(\design_top.core0.REG1[14][24] ),
    .B2(_09485_),
    .X(_04688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17065_ (.A1(_09383_),
    .A2(_09484_),
    .B1(\design_top.core0.REG1[14][23] ),
    .B2(_09485_),
    .X(_04687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17066_ (.A1(_09384_),
    .A2(_09484_),
    .B1(\design_top.core0.REG1[14][22] ),
    .B2(_09485_),
    .X(_04686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17067_ (.A(_09479_),
    .X(_09486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17068_ (.A(_09482_),
    .X(_09487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17069_ (.A1(_09385_),
    .A2(_09486_),
    .B1(\design_top.core0.REG1[14][21] ),
    .B2(_09487_),
    .X(_04685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17070_ (.A1(_09388_),
    .A2(_09486_),
    .B1(\design_top.core0.REG1[14][20] ),
    .B2(_09487_),
    .X(_04684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17071_ (.A1(_09389_),
    .A2(_09486_),
    .B1(\design_top.core0.REG1[14][19] ),
    .B2(_09487_),
    .X(_04683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17072_ (.A1(_09390_),
    .A2(_09486_),
    .B1(\design_top.core0.REG1[14][18] ),
    .B2(_09487_),
    .X(_04682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17073_ (.A1(_09391_),
    .A2(_09486_),
    .B1(\design_top.core0.REG1[14][17] ),
    .B2(_09487_),
    .X(_04681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17074_ (.A(_09478_),
    .X(_09488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17075_ (.A(_09481_),
    .X(_09489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17076_ (.A1(_09392_),
    .A2(_09488_),
    .B1(\design_top.core0.REG1[14][16] ),
    .B2(_09489_),
    .X(_04680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17077_ (.A1(_09395_),
    .A2(_09488_),
    .B1(\design_top.core0.REG1[14][15] ),
    .B2(_09489_),
    .X(_04679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17078_ (.A1(_09396_),
    .A2(_09488_),
    .B1(\design_top.core0.REG1[14][14] ),
    .B2(_09489_),
    .X(_04678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17079_ (.A(_00045_),
    .X(_09490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17080_ (.A1(\design_top.core0.REG1[14][13] ),
    .A2(_09479_),
    .B1(_09490_),
    .B2(_09482_),
    .X(_04677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17081_ (.A1(_09397_),
    .A2(_09488_),
    .B1(\design_top.core0.REG1[14][12] ),
    .B2(_09489_),
    .X(_04676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17082_ (.A1(_09398_),
    .A2(_09488_),
    .B1(\design_top.core0.REG1[14][11] ),
    .B2(_09489_),
    .X(_04675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17083_ (.A(_09478_),
    .X(_09491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17084_ (.A(_09481_),
    .X(_09492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17085_ (.A1(_09399_),
    .A2(_09491_),
    .B1(\design_top.core0.REG1[14][10] ),
    .B2(_09492_),
    .X(_04674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17086_ (.A1(_09402_),
    .A2(_09491_),
    .B1(\design_top.core0.REG1[14][9] ),
    .B2(_09492_),
    .X(_04673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17087_ (.A1(_09403_),
    .A2(_09491_),
    .B1(\design_top.core0.REG1[14][8] ),
    .B2(_09492_),
    .X(_04672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17088_ (.A1(_09404_),
    .A2(_09491_),
    .B1(\design_top.core0.REG1[14][7] ),
    .B2(_09492_),
    .X(_04671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17089_ (.A1(_09405_),
    .A2(_09491_),
    .B1(\design_top.core0.REG1[14][6] ),
    .B2(_09492_),
    .X(_04670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17090_ (.A(_09478_),
    .X(_09493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17091_ (.A(_09481_),
    .X(_09494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17092_ (.A1(_09406_),
    .A2(_09493_),
    .B1(\design_top.core0.REG1[14][5] ),
    .B2(_09494_),
    .X(_04669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17093_ (.A1(_09409_),
    .A2(_09493_),
    .B1(\design_top.core0.REG1[14][4] ),
    .B2(_09494_),
    .X(_04668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17094_ (.A1(_09410_),
    .A2(_09493_),
    .B1(\design_top.core0.REG1[14][3] ),
    .B2(_09494_),
    .X(_04667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17095_ (.A1(_09411_),
    .A2(_09493_),
    .B1(\design_top.core0.REG1[14][2] ),
    .B2(_09494_),
    .X(_04666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17096_ (.A1(_09412_),
    .A2(_09493_),
    .B1(\design_top.core0.REG1[14][1] ),
    .B2(_09494_),
    .X(_04665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17097_ (.A1(_09413_),
    .A2(_09479_),
    .B1(\design_top.core0.REG1[14][0] ),
    .B2(_09482_),
    .X(_04664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17098_ (.A(_09081_),
    .X(_09495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _17099_ (.A(_09477_),
    .B(_09166_),
    .X(_09496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17100_ (.A(_09496_),
    .X(_09497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17101_ (.A(_09497_),
    .X(_09498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17102_ (.A(_09496_),
    .Y(_09499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17103_ (.A(_09499_),
    .X(_09500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17104_ (.A(_09500_),
    .X(_09501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17105_ (.A1(_09495_),
    .A2(_09498_),
    .B1(\design_top.core0.REG1[13][31] ),
    .B2(_09501_),
    .X(_04663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17106_ (.A(_09095_),
    .X(_09502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17107_ (.A1(_09502_),
    .A2(_09498_),
    .B1(\design_top.core0.REG1[13][30] ),
    .B2(_09501_),
    .X(_04662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17108_ (.A(_09097_),
    .X(_09503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17109_ (.A1(_09503_),
    .A2(_09498_),
    .B1(\design_top.core0.REG1[13][29] ),
    .B2(_09501_),
    .X(_04661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17110_ (.A(_09099_),
    .X(_09504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17111_ (.A1(_09504_),
    .A2(_09498_),
    .B1(\design_top.core0.REG1[13][28] ),
    .B2(_09501_),
    .X(_04660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17112_ (.A(_09101_),
    .X(_09505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17113_ (.A1(_09505_),
    .A2(_09498_),
    .B1(\design_top.core0.REG1[13][27] ),
    .B2(_09501_),
    .X(_04659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17114_ (.A(_09103_),
    .X(_09506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17115_ (.A(_09497_),
    .X(_09507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17116_ (.A(_09500_),
    .X(_09508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17117_ (.A1(_09506_),
    .A2(_09507_),
    .B1(\design_top.core0.REG1[13][26] ),
    .B2(_09508_),
    .X(_04658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17118_ (.A(_09107_),
    .X(_09509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17119_ (.A1(_09509_),
    .A2(_09507_),
    .B1(\design_top.core0.REG1[13][25] ),
    .B2(_09508_),
    .X(_04657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17120_ (.A(_09109_),
    .X(_09510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17121_ (.A1(_09510_),
    .A2(_09507_),
    .B1(\design_top.core0.REG1[13][24] ),
    .B2(_09508_),
    .X(_04656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17122_ (.A(_09111_),
    .X(_09511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17123_ (.A1(_09511_),
    .A2(_09507_),
    .B1(\design_top.core0.REG1[13][23] ),
    .B2(_09508_),
    .X(_04655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17124_ (.A(_09113_),
    .X(_09512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17125_ (.A1(_09512_),
    .A2(_09507_),
    .B1(\design_top.core0.REG1[13][22] ),
    .B2(_09508_),
    .X(_04654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17126_ (.A(_09115_),
    .X(_09513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17127_ (.A(_09497_),
    .X(_09514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17128_ (.A(_09500_),
    .X(_09515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17129_ (.A1(_09513_),
    .A2(_09514_),
    .B1(\design_top.core0.REG1[13][21] ),
    .B2(_09515_),
    .X(_04653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17130_ (.A(_09119_),
    .X(_09516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17131_ (.A1(_09516_),
    .A2(_09514_),
    .B1(\design_top.core0.REG1[13][20] ),
    .B2(_09515_),
    .X(_04652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17132_ (.A(_09121_),
    .X(_09517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17133_ (.A1(_09517_),
    .A2(_09514_),
    .B1(\design_top.core0.REG1[13][19] ),
    .B2(_09515_),
    .X(_04651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17134_ (.A(_09123_),
    .X(_09518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17135_ (.A1(_09518_),
    .A2(_09514_),
    .B1(\design_top.core0.REG1[13][18] ),
    .B2(_09515_),
    .X(_04650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17136_ (.A(_09125_),
    .X(_09519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17137_ (.A1(_09519_),
    .A2(_09514_),
    .B1(\design_top.core0.REG1[13][17] ),
    .B2(_09515_),
    .X(_04649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17138_ (.A(_09127_),
    .X(_09520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17139_ (.A(_09496_),
    .X(_09521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17140_ (.A(_09499_),
    .X(_09522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17141_ (.A1(_09520_),
    .A2(_09521_),
    .B1(\design_top.core0.REG1[13][16] ),
    .B2(_09522_),
    .X(_04648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17142_ (.A(_09131_),
    .X(_09523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17143_ (.A1(_09523_),
    .A2(_09521_),
    .B1(\design_top.core0.REG1[13][15] ),
    .B2(_09522_),
    .X(_04647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17144_ (.A(_09133_),
    .X(_09524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17145_ (.A1(_09524_),
    .A2(_09521_),
    .B1(\design_top.core0.REG1[13][14] ),
    .B2(_09522_),
    .X(_04646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17146_ (.A1(\design_top.core0.REG1[13][13] ),
    .A2(_09497_),
    .B1(_09490_),
    .B2(_09500_),
    .X(_04645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17147_ (.A(_09136_),
    .X(_09525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17148_ (.A1(_09525_),
    .A2(_09521_),
    .B1(\design_top.core0.REG1[13][12] ),
    .B2(_09522_),
    .X(_04644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17149_ (.A(_09138_),
    .X(_09526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17150_ (.A1(_09526_),
    .A2(_09521_),
    .B1(\design_top.core0.REG1[13][11] ),
    .B2(_09522_),
    .X(_04643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17151_ (.A(_09140_),
    .X(_09527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17152_ (.A(_09496_),
    .X(_09528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17153_ (.A(_09499_),
    .X(_09529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17154_ (.A1(_09527_),
    .A2(_09528_),
    .B1(\design_top.core0.REG1[13][10] ),
    .B2(_09529_),
    .X(_04642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17155_ (.A(_09144_),
    .X(_09530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17156_ (.A1(_09530_),
    .A2(_09528_),
    .B1(\design_top.core0.REG1[13][9] ),
    .B2(_09529_),
    .X(_04641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17157_ (.A(_09146_),
    .X(_09531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17158_ (.A1(_09531_),
    .A2(_09528_),
    .B1(\design_top.core0.REG1[13][8] ),
    .B2(_09529_),
    .X(_04640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17159_ (.A(_09148_),
    .X(_09532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17160_ (.A1(_09532_),
    .A2(_09528_),
    .B1(\design_top.core0.REG1[13][7] ),
    .B2(_09529_),
    .X(_04639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17161_ (.A(_09150_),
    .X(_09533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17162_ (.A1(_09533_),
    .A2(_09528_),
    .B1(\design_top.core0.REG1[13][6] ),
    .B2(_09529_),
    .X(_04638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17163_ (.A(_09152_),
    .X(_09534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17164_ (.A(_09496_),
    .X(_09535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17165_ (.A(_09499_),
    .X(_09536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17166_ (.A1(_09534_),
    .A2(_09535_),
    .B1(\design_top.core0.REG1[13][5] ),
    .B2(_09536_),
    .X(_04637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17167_ (.A(_09156_),
    .X(_09537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17168_ (.A1(_09537_),
    .A2(_09535_),
    .B1(\design_top.core0.REG1[13][4] ),
    .B2(_09536_),
    .X(_04636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17169_ (.A(_09158_),
    .X(_09538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17170_ (.A1(_09538_),
    .A2(_09535_),
    .B1(\design_top.core0.REG1[13][3] ),
    .B2(_09536_),
    .X(_04635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17171_ (.A(_09160_),
    .X(_09539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17172_ (.A1(_09539_),
    .A2(_09535_),
    .B1(\design_top.core0.REG1[13][2] ),
    .B2(_09536_),
    .X(_04634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17173_ (.A(_09162_),
    .X(_09540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17174_ (.A1(_09540_),
    .A2(_09535_),
    .B1(\design_top.core0.REG1[13][1] ),
    .B2(_09536_),
    .X(_04633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17175_ (.A(_09164_),
    .X(_09541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17176_ (.A1(_09541_),
    .A2(_09497_),
    .B1(\design_top.core0.REG1[13][0] ),
    .B2(_09500_),
    .X(_04632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _17177_ (.A(_09477_),
    .B(_09183_),
    .X(_09542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17178_ (.A(_09542_),
    .X(_09543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17179_ (.A(_09543_),
    .X(_09544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17180_ (.A(_09542_),
    .Y(_09545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17181_ (.A(_09545_),
    .X(_09546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17182_ (.A(_09546_),
    .X(_09547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17183_ (.A1(_09495_),
    .A2(_09544_),
    .B1(\design_top.core0.REG1[12][31] ),
    .B2(_09547_),
    .X(_04631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17184_ (.A1(_09502_),
    .A2(_09544_),
    .B1(\design_top.core0.REG1[12][30] ),
    .B2(_09547_),
    .X(_04630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17185_ (.A1(_09503_),
    .A2(_09544_),
    .B1(\design_top.core0.REG1[12][29] ),
    .B2(_09547_),
    .X(_04629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17186_ (.A1(_09504_),
    .A2(_09544_),
    .B1(\design_top.core0.REG1[12][28] ),
    .B2(_09547_),
    .X(_04628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17187_ (.A1(_09505_),
    .A2(_09544_),
    .B1(\design_top.core0.REG1[12][27] ),
    .B2(_09547_),
    .X(_04627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17188_ (.A(_09543_),
    .X(_09548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17189_ (.A(_09546_),
    .X(_09549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17190_ (.A1(_09506_),
    .A2(_09548_),
    .B1(\design_top.core0.REG1[12][26] ),
    .B2(_09549_),
    .X(_04626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17191_ (.A1(_09509_),
    .A2(_09548_),
    .B1(\design_top.core0.REG1[12][25] ),
    .B2(_09549_),
    .X(_04625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17192_ (.A1(_09510_),
    .A2(_09548_),
    .B1(\design_top.core0.REG1[12][24] ),
    .B2(_09549_),
    .X(_04624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17193_ (.A1(_09511_),
    .A2(_09548_),
    .B1(\design_top.core0.REG1[12][23] ),
    .B2(_09549_),
    .X(_04623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17194_ (.A1(_09512_),
    .A2(_09548_),
    .B1(\design_top.core0.REG1[12][22] ),
    .B2(_09549_),
    .X(_04622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17195_ (.A(_09543_),
    .X(_09550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17196_ (.A(_09546_),
    .X(_09551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17197_ (.A1(_09513_),
    .A2(_09550_),
    .B1(\design_top.core0.REG1[12][21] ),
    .B2(_09551_),
    .X(_04621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17198_ (.A1(_09516_),
    .A2(_09550_),
    .B1(\design_top.core0.REG1[12][20] ),
    .B2(_09551_),
    .X(_04620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17199_ (.A1(_09517_),
    .A2(_09550_),
    .B1(\design_top.core0.REG1[12][19] ),
    .B2(_09551_),
    .X(_04619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17200_ (.A1(_09518_),
    .A2(_09550_),
    .B1(\design_top.core0.REG1[12][18] ),
    .B2(_09551_),
    .X(_04618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17201_ (.A1(_09519_),
    .A2(_09550_),
    .B1(\design_top.core0.REG1[12][17] ),
    .B2(_09551_),
    .X(_04617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17202_ (.A(_09542_),
    .X(_09552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17203_ (.A(_09545_),
    .X(_09553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17204_ (.A1(_09520_),
    .A2(_09552_),
    .B1(\design_top.core0.REG1[12][16] ),
    .B2(_09553_),
    .X(_04616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17205_ (.A1(_09523_),
    .A2(_09552_),
    .B1(\design_top.core0.REG1[12][15] ),
    .B2(_09553_),
    .X(_04615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17206_ (.A1(_09524_),
    .A2(_09552_),
    .B1(\design_top.core0.REG1[12][14] ),
    .B2(_09553_),
    .X(_04614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17207_ (.A1(\design_top.core0.REG1[12][13] ),
    .A2(_09543_),
    .B1(_09490_),
    .B2(_09546_),
    .X(_04613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17208_ (.A1(_09525_),
    .A2(_09552_),
    .B1(\design_top.core0.REG1[12][12] ),
    .B2(_09553_),
    .X(_04612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17209_ (.A1(_09526_),
    .A2(_09552_),
    .B1(\design_top.core0.REG1[12][11] ),
    .B2(_09553_),
    .X(_04611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17210_ (.A(_09542_),
    .X(_09554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17211_ (.A(_09545_),
    .X(_09555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17212_ (.A1(_09527_),
    .A2(_09554_),
    .B1(\design_top.core0.REG1[12][10] ),
    .B2(_09555_),
    .X(_04610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17213_ (.A1(_09530_),
    .A2(_09554_),
    .B1(\design_top.core0.REG1[12][9] ),
    .B2(_09555_),
    .X(_04609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17214_ (.A1(_09531_),
    .A2(_09554_),
    .B1(\design_top.core0.REG1[12][8] ),
    .B2(_09555_),
    .X(_04608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17215_ (.A1(_09532_),
    .A2(_09554_),
    .B1(\design_top.core0.REG1[12][7] ),
    .B2(_09555_),
    .X(_04607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17216_ (.A1(_09533_),
    .A2(_09554_),
    .B1(\design_top.core0.REG1[12][6] ),
    .B2(_09555_),
    .X(_04606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17217_ (.A(_09542_),
    .X(_09556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17218_ (.A(_09545_),
    .X(_09557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17219_ (.A1(_09534_),
    .A2(_09556_),
    .B1(\design_top.core0.REG1[12][5] ),
    .B2(_09557_),
    .X(_04605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17220_ (.A1(_09537_),
    .A2(_09556_),
    .B1(\design_top.core0.REG1[12][4] ),
    .B2(_09557_),
    .X(_04604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17221_ (.A1(_09538_),
    .A2(_09556_),
    .B1(\design_top.core0.REG1[12][3] ),
    .B2(_09557_),
    .X(_04603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17222_ (.A1(_09539_),
    .A2(_09556_),
    .B1(\design_top.core0.REG1[12][2] ),
    .B2(_09557_),
    .X(_04602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17223_ (.A1(_09540_),
    .A2(_09556_),
    .B1(\design_top.core0.REG1[12][1] ),
    .B2(_09557_),
    .X(_04601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17224_ (.A1(_09541_),
    .A2(_09543_),
    .B1(\design_top.core0.REG1[12][0] ),
    .B2(_09546_),
    .X(_04600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _17225_ (.A(_09477_),
    .B(_09201_),
    .X(_09558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17226_ (.A(_09558_),
    .X(_09559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17227_ (.A(_09559_),
    .X(_09560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17228_ (.A(_09558_),
    .Y(_09561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17229_ (.A(_09561_),
    .X(_09562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17230_ (.A(_09562_),
    .X(_09563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17231_ (.A1(_09495_),
    .A2(_09560_),
    .B1(\design_top.core0.REG1[11][31] ),
    .B2(_09563_),
    .X(_04599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17232_ (.A1(_09502_),
    .A2(_09560_),
    .B1(\design_top.core0.REG1[11][30] ),
    .B2(_09563_),
    .X(_04598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17233_ (.A1(_09503_),
    .A2(_09560_),
    .B1(\design_top.core0.REG1[11][29] ),
    .B2(_09563_),
    .X(_04597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17234_ (.A1(_09504_),
    .A2(_09560_),
    .B1(\design_top.core0.REG1[11][28] ),
    .B2(_09563_),
    .X(_04596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17235_ (.A1(_09505_),
    .A2(_09560_),
    .B1(\design_top.core0.REG1[11][27] ),
    .B2(_09563_),
    .X(_04595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17236_ (.A(_09559_),
    .X(_09564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17237_ (.A(_09562_),
    .X(_09565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17238_ (.A1(_09506_),
    .A2(_09564_),
    .B1(\design_top.core0.REG1[11][26] ),
    .B2(_09565_),
    .X(_04594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17239_ (.A1(_09509_),
    .A2(_09564_),
    .B1(\design_top.core0.REG1[11][25] ),
    .B2(_09565_),
    .X(_04593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17240_ (.A1(_09510_),
    .A2(_09564_),
    .B1(\design_top.core0.REG1[11][24] ),
    .B2(_09565_),
    .X(_04592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17241_ (.A1(_09511_),
    .A2(_09564_),
    .B1(\design_top.core0.REG1[11][23] ),
    .B2(_09565_),
    .X(_04591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17242_ (.A1(_09512_),
    .A2(_09564_),
    .B1(\design_top.core0.REG1[11][22] ),
    .B2(_09565_),
    .X(_04590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17243_ (.A(_09559_),
    .X(_09566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17244_ (.A(_09562_),
    .X(_09567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17245_ (.A1(_09513_),
    .A2(_09566_),
    .B1(\design_top.core0.REG1[11][21] ),
    .B2(_09567_),
    .X(_04589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17246_ (.A1(_09516_),
    .A2(_09566_),
    .B1(\design_top.core0.REG1[11][20] ),
    .B2(_09567_),
    .X(_04588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17247_ (.A1(_09517_),
    .A2(_09566_),
    .B1(\design_top.core0.REG1[11][19] ),
    .B2(_09567_),
    .X(_04587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17248_ (.A1(_09518_),
    .A2(_09566_),
    .B1(\design_top.core0.REG1[11][18] ),
    .B2(_09567_),
    .X(_04586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17249_ (.A1(_09519_),
    .A2(_09566_),
    .B1(\design_top.core0.REG1[11][17] ),
    .B2(_09567_),
    .X(_04585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17250_ (.A(_09558_),
    .X(_09568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17251_ (.A(_09561_),
    .X(_09569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17252_ (.A1(_09520_),
    .A2(_09568_),
    .B1(\design_top.core0.REG1[11][16] ),
    .B2(_09569_),
    .X(_04584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17253_ (.A1(_09523_),
    .A2(_09568_),
    .B1(\design_top.core0.REG1[11][15] ),
    .B2(_09569_),
    .X(_04583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17254_ (.A1(_09524_),
    .A2(_09568_),
    .B1(\design_top.core0.REG1[11][14] ),
    .B2(_09569_),
    .X(_04582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17255_ (.A1(\design_top.core0.REG1[11][13] ),
    .A2(_09559_),
    .B1(_09490_),
    .B2(_09562_),
    .X(_04581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17256_ (.A1(_09525_),
    .A2(_09568_),
    .B1(\design_top.core0.REG1[11][12] ),
    .B2(_09569_),
    .X(_04580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17257_ (.A1(_09526_),
    .A2(_09568_),
    .B1(\design_top.core0.REG1[11][11] ),
    .B2(_09569_),
    .X(_04579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17258_ (.A(_09558_),
    .X(_09570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17259_ (.A(_09561_),
    .X(_09571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17260_ (.A1(_09527_),
    .A2(_09570_),
    .B1(\design_top.core0.REG1[11][10] ),
    .B2(_09571_),
    .X(_04578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17261_ (.A1(_09530_),
    .A2(_09570_),
    .B1(\design_top.core0.REG1[11][9] ),
    .B2(_09571_),
    .X(_04577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17262_ (.A1(_09531_),
    .A2(_09570_),
    .B1(\design_top.core0.REG1[11][8] ),
    .B2(_09571_),
    .X(_04576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17263_ (.A1(_09532_),
    .A2(_09570_),
    .B1(\design_top.core0.REG1[11][7] ),
    .B2(_09571_),
    .X(_04575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17264_ (.A1(_09533_),
    .A2(_09570_),
    .B1(\design_top.core0.REG1[11][6] ),
    .B2(_09571_),
    .X(_04574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17265_ (.A(_09558_),
    .X(_09572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17266_ (.A(_09561_),
    .X(_09573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17267_ (.A1(_09534_),
    .A2(_09572_),
    .B1(\design_top.core0.REG1[11][5] ),
    .B2(_09573_),
    .X(_04573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17268_ (.A1(_09537_),
    .A2(_09572_),
    .B1(\design_top.core0.REG1[11][4] ),
    .B2(_09573_),
    .X(_04572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17269_ (.A1(_09538_),
    .A2(_09572_),
    .B1(\design_top.core0.REG1[11][3] ),
    .B2(_09573_),
    .X(_04571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17270_ (.A1(_09539_),
    .A2(_09572_),
    .B1(\design_top.core0.REG1[11][2] ),
    .B2(_09573_),
    .X(_04570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17271_ (.A1(_09540_),
    .A2(_09572_),
    .B1(\design_top.core0.REG1[11][1] ),
    .B2(_09573_),
    .X(_04569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17272_ (.A1(_09541_),
    .A2(_09559_),
    .B1(\design_top.core0.REG1[11][0] ),
    .B2(_09562_),
    .X(_04568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17273_ (.A(_08789_),
    .X(_09574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _17274_ (.A(_09574_),
    .B(_09218_),
    .X(_09575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17275_ (.A(_09575_),
    .X(_09576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17276_ (.A(_09576_),
    .X(_09577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17277_ (.A(_09575_),
    .Y(_09578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17278_ (.A(_09578_),
    .X(_09579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17279_ (.A(_09579_),
    .X(_09580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17280_ (.A1(_09495_),
    .A2(_09577_),
    .B1(\design_top.core0.REG1[10][31] ),
    .B2(_09580_),
    .X(_04567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17281_ (.A1(_09502_),
    .A2(_09577_),
    .B1(\design_top.core0.REG1[10][30] ),
    .B2(_09580_),
    .X(_04566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17282_ (.A1(_09503_),
    .A2(_09577_),
    .B1(\design_top.core0.REG1[10][29] ),
    .B2(_09580_),
    .X(_04565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17283_ (.A1(_09504_),
    .A2(_09577_),
    .B1(\design_top.core0.REG1[10][28] ),
    .B2(_09580_),
    .X(_04564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17284_ (.A1(_09505_),
    .A2(_09577_),
    .B1(\design_top.core0.REG1[10][27] ),
    .B2(_09580_),
    .X(_04563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17285_ (.A(_09576_),
    .X(_09581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17286_ (.A(_09579_),
    .X(_09582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17287_ (.A1(_09506_),
    .A2(_09581_),
    .B1(\design_top.core0.REG1[10][26] ),
    .B2(_09582_),
    .X(_04562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17288_ (.A1(_09509_),
    .A2(_09581_),
    .B1(\design_top.core0.REG1[10][25] ),
    .B2(_09582_),
    .X(_04561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17289_ (.A1(_09510_),
    .A2(_09581_),
    .B1(\design_top.core0.REG1[10][24] ),
    .B2(_09582_),
    .X(_04560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17290_ (.A1(_09511_),
    .A2(_09581_),
    .B1(\design_top.core0.REG1[10][23] ),
    .B2(_09582_),
    .X(_04559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17291_ (.A1(_09512_),
    .A2(_09581_),
    .B1(\design_top.core0.REG1[10][22] ),
    .B2(_09582_),
    .X(_04558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17292_ (.A(_09576_),
    .X(_09583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17293_ (.A(_09579_),
    .X(_09584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17294_ (.A1(_09513_),
    .A2(_09583_),
    .B1(\design_top.core0.REG1[10][21] ),
    .B2(_09584_),
    .X(_04557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17295_ (.A1(_09516_),
    .A2(_09583_),
    .B1(\design_top.core0.REG1[10][20] ),
    .B2(_09584_),
    .X(_04556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17296_ (.A1(_09517_),
    .A2(_09583_),
    .B1(\design_top.core0.REG1[10][19] ),
    .B2(_09584_),
    .X(_04555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17297_ (.A1(_09518_),
    .A2(_09583_),
    .B1(\design_top.core0.REG1[10][18] ),
    .B2(_09584_),
    .X(_04554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17298_ (.A1(_09519_),
    .A2(_09583_),
    .B1(\design_top.core0.REG1[10][17] ),
    .B2(_09584_),
    .X(_04553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17299_ (.A(_09575_),
    .X(_09585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17300_ (.A(_09578_),
    .X(_09586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17301_ (.A1(_09520_),
    .A2(_09585_),
    .B1(\design_top.core0.REG1[10][16] ),
    .B2(_09586_),
    .X(_04552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17302_ (.A1(_09523_),
    .A2(_09585_),
    .B1(\design_top.core0.REG1[10][15] ),
    .B2(_09586_),
    .X(_04551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17303_ (.A1(_09524_),
    .A2(_09585_),
    .B1(\design_top.core0.REG1[10][14] ),
    .B2(_09586_),
    .X(_04550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17304_ (.A1(\design_top.core0.REG1[10][13] ),
    .A2(_09576_),
    .B1(_09490_),
    .B2(_09579_),
    .X(_04549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17305_ (.A1(_09525_),
    .A2(_09585_),
    .B1(\design_top.core0.REG1[10][12] ),
    .B2(_09586_),
    .X(_04548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17306_ (.A1(_09526_),
    .A2(_09585_),
    .B1(\design_top.core0.REG1[10][11] ),
    .B2(_09586_),
    .X(_04547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17307_ (.A(_09575_),
    .X(_09587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17308_ (.A(_09578_),
    .X(_09588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17309_ (.A1(_09527_),
    .A2(_09587_),
    .B1(\design_top.core0.REG1[10][10] ),
    .B2(_09588_),
    .X(_04546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17310_ (.A1(_09530_),
    .A2(_09587_),
    .B1(\design_top.core0.REG1[10][9] ),
    .B2(_09588_),
    .X(_04545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17311_ (.A1(_09531_),
    .A2(_09587_),
    .B1(\design_top.core0.REG1[10][8] ),
    .B2(_09588_),
    .X(_04544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17312_ (.A1(_09532_),
    .A2(_09587_),
    .B1(\design_top.core0.REG1[10][7] ),
    .B2(_09588_),
    .X(_04543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17313_ (.A1(_09533_),
    .A2(_09587_),
    .B1(\design_top.core0.REG1[10][6] ),
    .B2(_09588_),
    .X(_04542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17314_ (.A(_09575_),
    .X(_09589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17315_ (.A(_09578_),
    .X(_09590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17316_ (.A1(_09534_),
    .A2(_09589_),
    .B1(\design_top.core0.REG1[10][5] ),
    .B2(_09590_),
    .X(_04541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17317_ (.A1(_09537_),
    .A2(_09589_),
    .B1(\design_top.core0.REG1[10][4] ),
    .B2(_09590_),
    .X(_04540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17318_ (.A1(_09538_),
    .A2(_09589_),
    .B1(\design_top.core0.REG1[10][3] ),
    .B2(_09590_),
    .X(_04539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17319_ (.A1(_09539_),
    .A2(_09589_),
    .B1(\design_top.core0.REG1[10][2] ),
    .B2(_09590_),
    .X(_04538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17320_ (.A1(_09540_),
    .A2(_09589_),
    .B1(\design_top.core0.REG1[10][1] ),
    .B2(_09590_),
    .X(_04537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17321_ (.A1(_09541_),
    .A2(_09576_),
    .B1(\design_top.core0.REG1[10][0] ),
    .B2(_09579_),
    .X(_04536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17322_ (.A(\design_top.core0.REG1[0][31] ),
    .Y(_02664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _17323_ (.A(_09235_),
    .B(_09477_),
    .X(_09591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17324_ (.A(_09591_),
    .X(_09592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17325_ (.A(_09592_),
    .Y(_09593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _17326_ (.A(_02664_),
    .B(_09593_),
    .Y(_04535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17327_ (.A(_09592_),
    .X(_09594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17328_ (.A(\design_top.core0.REG1[0][30] ),
    .B(_09594_),
    .X(_04534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17329_ (.A(\design_top.core0.REG1[0][29] ),
    .B(_09594_),
    .X(_04533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17330_ (.A(\design_top.core0.REG1[0][28] ),
    .B(_09594_),
    .X(_04532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17331_ (.A(\design_top.core0.REG1[0][27] ),
    .B(_09594_),
    .X(_04531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17332_ (.A(\design_top.core0.REG1[0][26] ),
    .B(_09594_),
    .X(_04530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17333_ (.A(_09592_),
    .X(_09595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17334_ (.A(\design_top.core0.REG1[0][25] ),
    .B(_09595_),
    .X(_04529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17335_ (.A(\design_top.core0.REG1[0][24] ),
    .B(_09595_),
    .X(_04528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17336_ (.A(\design_top.core0.REG1[0][23] ),
    .B(_09595_),
    .X(_04527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17337_ (.A(\design_top.core0.REG1[0][22] ),
    .B(_09595_),
    .X(_04526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17338_ (.A(\design_top.core0.REG1[0][21] ),
    .B(_09595_),
    .X(_04525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17339_ (.A(_09592_),
    .X(_09596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17340_ (.A(\design_top.core0.REG1[0][20] ),
    .B(_09596_),
    .X(_04524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17341_ (.A(\design_top.core0.REG1[0][19] ),
    .B(_09596_),
    .X(_04523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17342_ (.A(\design_top.core0.REG1[0][18] ),
    .B(_09596_),
    .X(_04522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17343_ (.A(\design_top.core0.REG1[0][17] ),
    .B(_09596_),
    .X(_04521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17344_ (.A(\design_top.core0.REG1[0][16] ),
    .B(_09596_),
    .X(_04520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17345_ (.A(_09591_),
    .X(_09597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17346_ (.A(\design_top.core0.REG1[0][15] ),
    .B(_09597_),
    .X(_04519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17347_ (.A(\design_top.core0.REG1[0][14] ),
    .B(_09597_),
    .X(_04518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17348_ (.A(_00045_),
    .X(_09598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17349_ (.A1(\design_top.core0.REG1[0][13] ),
    .A2(_09592_),
    .B1(_09598_),
    .B2(_09593_),
    .X(_04517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17350_ (.A(\design_top.core0.REG1[0][12] ),
    .B(_09597_),
    .X(_04516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17351_ (.A(\design_top.core0.REG1[0][11] ),
    .B(_09597_),
    .X(_04515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17352_ (.A(\design_top.core0.REG1[0][10] ),
    .B(_09597_),
    .X(_04514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17353_ (.A(_09591_),
    .X(_09599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17354_ (.A(\design_top.core0.REG1[0][9] ),
    .B(_09599_),
    .X(_04513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17355_ (.A(\design_top.core0.REG1[0][8] ),
    .B(_09599_),
    .X(_04512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17356_ (.A(\design_top.core0.REG1[0][7] ),
    .B(_09599_),
    .X(_04511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17357_ (.A(\design_top.core0.REG1[0][6] ),
    .B(_09599_),
    .X(_04510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17358_ (.A(\design_top.core0.REG1[0][5] ),
    .B(_09599_),
    .X(_04509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17359_ (.A(_09591_),
    .X(_09600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17360_ (.A(\design_top.core0.REG1[0][4] ),
    .B(_09600_),
    .X(_04508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17361_ (.A(\design_top.core0.REG1[0][3] ),
    .B(_09600_),
    .X(_04507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17362_ (.A(\design_top.core0.REG1[0][2] ),
    .B(_09600_),
    .X(_04506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17363_ (.A(\design_top.core0.REG1[0][1] ),
    .B(_09600_),
    .X(_04505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _17364_ (.A(\design_top.core0.REG1[0][0] ),
    .B(_09600_),
    .X(_04504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _17365_ (.A(_09574_),
    .B(_09245_),
    .X(_09601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17366_ (.A(_09601_),
    .X(_09602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17367_ (.A(_09602_),
    .X(_09603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17368_ (.A(_09601_),
    .Y(_09604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17369_ (.A(_09604_),
    .X(_09605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17370_ (.A(_09605_),
    .X(_09606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17371_ (.A1(_09495_),
    .A2(_09603_),
    .B1(\design_top.core0.REG1[8][31] ),
    .B2(_09606_),
    .X(_04503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17372_ (.A1(_09502_),
    .A2(_09603_),
    .B1(\design_top.core0.REG1[8][30] ),
    .B2(_09606_),
    .X(_04502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17373_ (.A1(_09503_),
    .A2(_09603_),
    .B1(\design_top.core0.REG1[8][29] ),
    .B2(_09606_),
    .X(_04501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17374_ (.A1(_09504_),
    .A2(_09603_),
    .B1(\design_top.core0.REG1[8][28] ),
    .B2(_09606_),
    .X(_04500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17375_ (.A1(_09505_),
    .A2(_09603_),
    .B1(\design_top.core0.REG1[8][27] ),
    .B2(_09606_),
    .X(_04499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17376_ (.A(_09602_),
    .X(_09607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17377_ (.A(_09605_),
    .X(_09608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17378_ (.A1(_09506_),
    .A2(_09607_),
    .B1(\design_top.core0.REG1[8][26] ),
    .B2(_09608_),
    .X(_04498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17379_ (.A1(_09509_),
    .A2(_09607_),
    .B1(\design_top.core0.REG1[8][25] ),
    .B2(_09608_),
    .X(_04497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17380_ (.A1(_09510_),
    .A2(_09607_),
    .B1(\design_top.core0.REG1[8][24] ),
    .B2(_09608_),
    .X(_04496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17381_ (.A1(_09511_),
    .A2(_09607_),
    .B1(\design_top.core0.REG1[8][23] ),
    .B2(_09608_),
    .X(_04495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17382_ (.A1(_09512_),
    .A2(_09607_),
    .B1(\design_top.core0.REG1[8][22] ),
    .B2(_09608_),
    .X(_04494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17383_ (.A(_09602_),
    .X(_09609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17384_ (.A(_09605_),
    .X(_09610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17385_ (.A1(_09513_),
    .A2(_09609_),
    .B1(\design_top.core0.REG1[8][21] ),
    .B2(_09610_),
    .X(_04493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17386_ (.A1(_09516_),
    .A2(_09609_),
    .B1(\design_top.core0.REG1[8][20] ),
    .B2(_09610_),
    .X(_04492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17387_ (.A1(_09517_),
    .A2(_09609_),
    .B1(\design_top.core0.REG1[8][19] ),
    .B2(_09610_),
    .X(_04491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17388_ (.A1(_09518_),
    .A2(_09609_),
    .B1(\design_top.core0.REG1[8][18] ),
    .B2(_09610_),
    .X(_04490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17389_ (.A1(_09519_),
    .A2(_09609_),
    .B1(\design_top.core0.REG1[8][17] ),
    .B2(_09610_),
    .X(_04489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17390_ (.A(_09601_),
    .X(_09611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17391_ (.A(_09604_),
    .X(_09612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17392_ (.A1(_09520_),
    .A2(_09611_),
    .B1(\design_top.core0.REG1[8][16] ),
    .B2(_09612_),
    .X(_04488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17393_ (.A1(_09523_),
    .A2(_09611_),
    .B1(\design_top.core0.REG1[8][15] ),
    .B2(_09612_),
    .X(_04487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17394_ (.A1(_09524_),
    .A2(_09611_),
    .B1(\design_top.core0.REG1[8][14] ),
    .B2(_09612_),
    .X(_04486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17395_ (.A1(\design_top.core0.REG1[8][13] ),
    .A2(_09602_),
    .B1(_09598_),
    .B2(_09605_),
    .X(_04485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17396_ (.A1(_09525_),
    .A2(_09611_),
    .B1(\design_top.core0.REG1[8][12] ),
    .B2(_09612_),
    .X(_04484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17397_ (.A1(_09526_),
    .A2(_09611_),
    .B1(\design_top.core0.REG1[8][11] ),
    .B2(_09612_),
    .X(_04483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17398_ (.A(_09601_),
    .X(_09613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17399_ (.A(_09604_),
    .X(_09614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17400_ (.A1(_09527_),
    .A2(_09613_),
    .B1(\design_top.core0.REG1[8][10] ),
    .B2(_09614_),
    .X(_04482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17401_ (.A1(_09530_),
    .A2(_09613_),
    .B1(\design_top.core0.REG1[8][9] ),
    .B2(_09614_),
    .X(_04481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17402_ (.A1(_09531_),
    .A2(_09613_),
    .B1(\design_top.core0.REG1[8][8] ),
    .B2(_09614_),
    .X(_04480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17403_ (.A1(_09532_),
    .A2(_09613_),
    .B1(\design_top.core0.REG1[8][7] ),
    .B2(_09614_),
    .X(_04479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17404_ (.A1(_09533_),
    .A2(_09613_),
    .B1(\design_top.core0.REG1[8][6] ),
    .B2(_09614_),
    .X(_04478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17405_ (.A(_09601_),
    .X(_09615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17406_ (.A(_09604_),
    .X(_09616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17407_ (.A1(_09534_),
    .A2(_09615_),
    .B1(\design_top.core0.REG1[8][5] ),
    .B2(_09616_),
    .X(_04477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17408_ (.A1(_09537_),
    .A2(_09615_),
    .B1(\design_top.core0.REG1[8][4] ),
    .B2(_09616_),
    .X(_04476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17409_ (.A1(_09538_),
    .A2(_09615_),
    .B1(\design_top.core0.REG1[8][3] ),
    .B2(_09616_),
    .X(_04475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17410_ (.A1(_09539_),
    .A2(_09615_),
    .B1(\design_top.core0.REG1[8][2] ),
    .B2(_09616_),
    .X(_04474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17411_ (.A1(_09540_),
    .A2(_09615_),
    .B1(\design_top.core0.REG1[8][1] ),
    .B2(_09616_),
    .X(_04473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17412_ (.A1(_09541_),
    .A2(_09602_),
    .B1(\design_top.core0.REG1[8][0] ),
    .B2(_09605_),
    .X(_04472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17413_ (.A(_09081_),
    .X(_09617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _17414_ (.A(_09574_),
    .B(_09293_),
    .X(_09618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17415_ (.A(_09618_),
    .X(_09619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17416_ (.A(_09619_),
    .X(_09620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17417_ (.A(_09618_),
    .Y(_09621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17418_ (.A(_09621_),
    .X(_09622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17419_ (.A(_09622_),
    .X(_09623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17420_ (.A1(_09617_),
    .A2(_09620_),
    .B1(\design_top.core0.REG1[7][31] ),
    .B2(_09623_),
    .X(_04471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17421_ (.A(_09095_),
    .X(_09624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17422_ (.A1(_09624_),
    .A2(_09620_),
    .B1(\design_top.core0.REG1[7][30] ),
    .B2(_09623_),
    .X(_04470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17423_ (.A(_09097_),
    .X(_09625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17424_ (.A1(_09625_),
    .A2(_09620_),
    .B1(\design_top.core0.REG1[7][29] ),
    .B2(_09623_),
    .X(_04469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17425_ (.A(_09099_),
    .X(_09626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17426_ (.A1(_09626_),
    .A2(_09620_),
    .B1(\design_top.core0.REG1[7][28] ),
    .B2(_09623_),
    .X(_04468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17427_ (.A(_09101_),
    .X(_09627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17428_ (.A1(_09627_),
    .A2(_09620_),
    .B1(\design_top.core0.REG1[7][27] ),
    .B2(_09623_),
    .X(_04467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17429_ (.A(_09103_),
    .X(_09628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17430_ (.A(_09619_),
    .X(_09629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17431_ (.A(_09622_),
    .X(_09630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17432_ (.A1(_09628_),
    .A2(_09629_),
    .B1(\design_top.core0.REG1[7][26] ),
    .B2(_09630_),
    .X(_04466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17433_ (.A(_09107_),
    .X(_09631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17434_ (.A1(_09631_),
    .A2(_09629_),
    .B1(\design_top.core0.REG1[7][25] ),
    .B2(_09630_),
    .X(_04465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17435_ (.A(_09109_),
    .X(_09632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17436_ (.A1(_09632_),
    .A2(_09629_),
    .B1(\design_top.core0.REG1[7][24] ),
    .B2(_09630_),
    .X(_04464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17437_ (.A(_09111_),
    .X(_09633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17438_ (.A1(_09633_),
    .A2(_09629_),
    .B1(\design_top.core0.REG1[7][23] ),
    .B2(_09630_),
    .X(_04463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17439_ (.A(_09113_),
    .X(_09634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17440_ (.A1(_09634_),
    .A2(_09629_),
    .B1(\design_top.core0.REG1[7][22] ),
    .B2(_09630_),
    .X(_04462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17441_ (.A(_09115_),
    .X(_09635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17442_ (.A(_09619_),
    .X(_09636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17443_ (.A(_09622_),
    .X(_09637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17444_ (.A1(_09635_),
    .A2(_09636_),
    .B1(\design_top.core0.REG1[7][21] ),
    .B2(_09637_),
    .X(_04461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17445_ (.A(_09119_),
    .X(_09638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17446_ (.A1(_09638_),
    .A2(_09636_),
    .B1(\design_top.core0.REG1[7][20] ),
    .B2(_09637_),
    .X(_04460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17447_ (.A(_09121_),
    .X(_09639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17448_ (.A1(_09639_),
    .A2(_09636_),
    .B1(\design_top.core0.REG1[7][19] ),
    .B2(_09637_),
    .X(_04459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17449_ (.A(_09123_),
    .X(_09640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17450_ (.A1(_09640_),
    .A2(_09636_),
    .B1(\design_top.core0.REG1[7][18] ),
    .B2(_09637_),
    .X(_04458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17451_ (.A(_09125_),
    .X(_09641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17452_ (.A1(_09641_),
    .A2(_09636_),
    .B1(\design_top.core0.REG1[7][17] ),
    .B2(_09637_),
    .X(_04457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17453_ (.A(_09127_),
    .X(_09642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17454_ (.A(_09618_),
    .X(_09643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17455_ (.A(_09621_),
    .X(_09644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17456_ (.A1(_09642_),
    .A2(_09643_),
    .B1(\design_top.core0.REG1[7][16] ),
    .B2(_09644_),
    .X(_04456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17457_ (.A(_09131_),
    .X(_09645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17458_ (.A1(_09645_),
    .A2(_09643_),
    .B1(\design_top.core0.REG1[7][15] ),
    .B2(_09644_),
    .X(_04455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17459_ (.A(_09133_),
    .X(_09646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17460_ (.A1(_09646_),
    .A2(_09643_),
    .B1(\design_top.core0.REG1[7][14] ),
    .B2(_09644_),
    .X(_04454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17461_ (.A1(\design_top.core0.REG1[7][13] ),
    .A2(_09619_),
    .B1(_09598_),
    .B2(_09622_),
    .X(_04453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17462_ (.A(_09136_),
    .X(_09647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17463_ (.A1(_09647_),
    .A2(_09643_),
    .B1(\design_top.core0.REG1[7][12] ),
    .B2(_09644_),
    .X(_04452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17464_ (.A(_09138_),
    .X(_09648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17465_ (.A1(_09648_),
    .A2(_09643_),
    .B1(\design_top.core0.REG1[7][11] ),
    .B2(_09644_),
    .X(_04451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17466_ (.A(_09140_),
    .X(_09649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17467_ (.A(_09618_),
    .X(_09650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17468_ (.A(_09621_),
    .X(_09651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17469_ (.A1(_09649_),
    .A2(_09650_),
    .B1(\design_top.core0.REG1[7][10] ),
    .B2(_09651_),
    .X(_04450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17470_ (.A(_09144_),
    .X(_09652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17471_ (.A1(_09652_),
    .A2(_09650_),
    .B1(\design_top.core0.REG1[7][9] ),
    .B2(_09651_),
    .X(_04449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17472_ (.A(_09146_),
    .X(_09653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17473_ (.A1(_09653_),
    .A2(_09650_),
    .B1(\design_top.core0.REG1[7][8] ),
    .B2(_09651_),
    .X(_04448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17474_ (.A(_09148_),
    .X(_09654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17475_ (.A1(_09654_),
    .A2(_09650_),
    .B1(\design_top.core0.REG1[7][7] ),
    .B2(_09651_),
    .X(_04447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17476_ (.A(_09150_),
    .X(_09655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17477_ (.A1(_09655_),
    .A2(_09650_),
    .B1(\design_top.core0.REG1[7][6] ),
    .B2(_09651_),
    .X(_04446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17478_ (.A(_09152_),
    .X(_09656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17479_ (.A(_09618_),
    .X(_09657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17480_ (.A(_09621_),
    .X(_09658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17481_ (.A1(_09656_),
    .A2(_09657_),
    .B1(\design_top.core0.REG1[7][5] ),
    .B2(_09658_),
    .X(_04445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17482_ (.A(_09156_),
    .X(_09659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17483_ (.A1(_09659_),
    .A2(_09657_),
    .B1(\design_top.core0.REG1[7][4] ),
    .B2(_09658_),
    .X(_04444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17484_ (.A(_09158_),
    .X(_09660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17485_ (.A1(_09660_),
    .A2(_09657_),
    .B1(\design_top.core0.REG1[7][3] ),
    .B2(_09658_),
    .X(_04443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17486_ (.A(_09160_),
    .X(_09661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17487_ (.A1(_09661_),
    .A2(_09657_),
    .B1(\design_top.core0.REG1[7][2] ),
    .B2(_09658_),
    .X(_04442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17488_ (.A(_09162_),
    .X(_09662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17489_ (.A1(_09662_),
    .A2(_09657_),
    .B1(\design_top.core0.REG1[7][1] ),
    .B2(_09658_),
    .X(_04441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17490_ (.A(_09164_),
    .X(_09663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17491_ (.A1(_09663_),
    .A2(_09619_),
    .B1(\design_top.core0.REG1[7][0] ),
    .B2(_09622_),
    .X(_04440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _17492_ (.A(_09574_),
    .B(_09310_),
    .X(_09664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17493_ (.A(_09664_),
    .X(_09665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17494_ (.A(_09665_),
    .X(_09666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17495_ (.A(_09664_),
    .Y(_09667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17496_ (.A(_09667_),
    .X(_09668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17497_ (.A(_09668_),
    .X(_09669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17498_ (.A1(_09617_),
    .A2(_09666_),
    .B1(\design_top.core0.REG1[6][31] ),
    .B2(_09669_),
    .X(_04439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17499_ (.A1(_09624_),
    .A2(_09666_),
    .B1(\design_top.core0.REG1[6][30] ),
    .B2(_09669_),
    .X(_04438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17500_ (.A1(_09625_),
    .A2(_09666_),
    .B1(\design_top.core0.REG1[6][29] ),
    .B2(_09669_),
    .X(_04437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17501_ (.A1(_09626_),
    .A2(_09666_),
    .B1(\design_top.core0.REG1[6][28] ),
    .B2(_09669_),
    .X(_04436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17502_ (.A1(_09627_),
    .A2(_09666_),
    .B1(\design_top.core0.REG1[6][27] ),
    .B2(_09669_),
    .X(_04435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17503_ (.A(_09665_),
    .X(_09670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17504_ (.A(_09668_),
    .X(_09671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17505_ (.A1(_09628_),
    .A2(_09670_),
    .B1(\design_top.core0.REG1[6][26] ),
    .B2(_09671_),
    .X(_04434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17506_ (.A1(_09631_),
    .A2(_09670_),
    .B1(\design_top.core0.REG1[6][25] ),
    .B2(_09671_),
    .X(_04433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17507_ (.A1(_09632_),
    .A2(_09670_),
    .B1(\design_top.core0.REG1[6][24] ),
    .B2(_09671_),
    .X(_04432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17508_ (.A1(_09633_),
    .A2(_09670_),
    .B1(\design_top.core0.REG1[6][23] ),
    .B2(_09671_),
    .X(_04431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17509_ (.A1(_09634_),
    .A2(_09670_),
    .B1(\design_top.core0.REG1[6][22] ),
    .B2(_09671_),
    .X(_04430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17510_ (.A(_09665_),
    .X(_09672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17511_ (.A(_09668_),
    .X(_09673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17512_ (.A1(_09635_),
    .A2(_09672_),
    .B1(\design_top.core0.REG1[6][21] ),
    .B2(_09673_),
    .X(_04429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17513_ (.A1(_09638_),
    .A2(_09672_),
    .B1(\design_top.core0.REG1[6][20] ),
    .B2(_09673_),
    .X(_04428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17514_ (.A1(_09639_),
    .A2(_09672_),
    .B1(\design_top.core0.REG1[6][19] ),
    .B2(_09673_),
    .X(_04427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17515_ (.A1(_09640_),
    .A2(_09672_),
    .B1(\design_top.core0.REG1[6][18] ),
    .B2(_09673_),
    .X(_04426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17516_ (.A1(_09641_),
    .A2(_09672_),
    .B1(\design_top.core0.REG1[6][17] ),
    .B2(_09673_),
    .X(_04425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17517_ (.A(_09664_),
    .X(_09674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17518_ (.A(_09667_),
    .X(_09675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17519_ (.A1(_09642_),
    .A2(_09674_),
    .B1(\design_top.core0.REG1[6][16] ),
    .B2(_09675_),
    .X(_04424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17520_ (.A1(_09645_),
    .A2(_09674_),
    .B1(\design_top.core0.REG1[6][15] ),
    .B2(_09675_),
    .X(_04423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17521_ (.A1(_09646_),
    .A2(_09674_),
    .B1(\design_top.core0.REG1[6][14] ),
    .B2(_09675_),
    .X(_04422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17522_ (.A1(\design_top.core0.REG1[6][13] ),
    .A2(_09665_),
    .B1(_09598_),
    .B2(_09668_),
    .X(_04421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17523_ (.A1(_09647_),
    .A2(_09674_),
    .B1(\design_top.core0.REG1[6][12] ),
    .B2(_09675_),
    .X(_04420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17524_ (.A1(_09648_),
    .A2(_09674_),
    .B1(\design_top.core0.REG1[6][11] ),
    .B2(_09675_),
    .X(_04419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17525_ (.A(_09664_),
    .X(_09676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17526_ (.A(_09667_),
    .X(_09677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17527_ (.A1(_09649_),
    .A2(_09676_),
    .B1(\design_top.core0.REG1[6][10] ),
    .B2(_09677_),
    .X(_04418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17528_ (.A1(_09652_),
    .A2(_09676_),
    .B1(\design_top.core0.REG1[6][9] ),
    .B2(_09677_),
    .X(_04417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17529_ (.A1(_09653_),
    .A2(_09676_),
    .B1(\design_top.core0.REG1[6][8] ),
    .B2(_09677_),
    .X(_04416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17530_ (.A1(_09654_),
    .A2(_09676_),
    .B1(\design_top.core0.REG1[6][7] ),
    .B2(_09677_),
    .X(_04415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17531_ (.A1(_09655_),
    .A2(_09676_),
    .B1(\design_top.core0.REG1[6][6] ),
    .B2(_09677_),
    .X(_04414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17532_ (.A(_09664_),
    .X(_09678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17533_ (.A(_09667_),
    .X(_09679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17534_ (.A1(_09656_),
    .A2(_09678_),
    .B1(\design_top.core0.REG1[6][5] ),
    .B2(_09679_),
    .X(_04413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17535_ (.A1(_09659_),
    .A2(_09678_),
    .B1(\design_top.core0.REG1[6][4] ),
    .B2(_09679_),
    .X(_04412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17536_ (.A1(_09660_),
    .A2(_09678_),
    .B1(\design_top.core0.REG1[6][3] ),
    .B2(_09679_),
    .X(_04411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17537_ (.A1(_09661_),
    .A2(_09678_),
    .B1(\design_top.core0.REG1[6][2] ),
    .B2(_09679_),
    .X(_04410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17538_ (.A1(_09662_),
    .A2(_09678_),
    .B1(\design_top.core0.REG1[6][1] ),
    .B2(_09679_),
    .X(_04409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17539_ (.A1(_09663_),
    .A2(_09665_),
    .B1(\design_top.core0.REG1[6][0] ),
    .B2(_09668_),
    .X(_04408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17540_ (.A(_09010_),
    .X(_09680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17541_ (.A1(_09050_),
    .A2(_08169_),
    .B1(_08224_),
    .B2(_09680_),
    .X(_09681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17542_ (.A(_09681_),
    .Y(_09682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17543_ (.A(_09682_),
    .X(_09683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17544_ (.A(_09681_),
    .X(_09684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17545_ (.A1(_00636_),
    .A2(_09683_),
    .B1(\design_top.MEM[61][7] ),
    .B2(_09684_),
    .X(_04407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17546_ (.A1(_00635_),
    .A2(_09683_),
    .B1(\design_top.MEM[61][6] ),
    .B2(_09684_),
    .X(_04406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17547_ (.A1(_00634_),
    .A2(_09683_),
    .B1(\design_top.MEM[61][5] ),
    .B2(_09684_),
    .X(_04405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17548_ (.A1(_00633_),
    .A2(_09683_),
    .B1(\design_top.MEM[61][4] ),
    .B2(_09684_),
    .X(_04404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17549_ (.A1(_00632_),
    .A2(_09683_),
    .B1(\design_top.MEM[61][3] ),
    .B2(_09684_),
    .X(_04403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17550_ (.A1(_00631_),
    .A2(_09682_),
    .B1(\design_top.MEM[61][2] ),
    .B2(_09681_),
    .X(_04402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17551_ (.A1(_00630_),
    .A2(_09682_),
    .B1(\design_top.MEM[61][1] ),
    .B2(_09681_),
    .X(_04401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17552_ (.A1(_00629_),
    .A2(_09682_),
    .B1(\design_top.MEM[61][0] ),
    .B2(_09681_),
    .X(_04400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _17553_ (.A(_09574_),
    .B(_09327_),
    .X(_09685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17554_ (.A(_09685_),
    .X(_09686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17555_ (.A(_09686_),
    .X(_09687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17556_ (.A(_09685_),
    .Y(_09688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17557_ (.A(_09688_),
    .X(_09689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17558_ (.A(_09689_),
    .X(_09690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17559_ (.A1(_09617_),
    .A2(_09687_),
    .B1(\design_top.core0.REG1[5][31] ),
    .B2(_09690_),
    .X(_04399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17560_ (.A1(_09624_),
    .A2(_09687_),
    .B1(\design_top.core0.REG1[5][30] ),
    .B2(_09690_),
    .X(_04398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17561_ (.A1(_09625_),
    .A2(_09687_),
    .B1(\design_top.core0.REG1[5][29] ),
    .B2(_09690_),
    .X(_04397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17562_ (.A1(_09626_),
    .A2(_09687_),
    .B1(\design_top.core0.REG1[5][28] ),
    .B2(_09690_),
    .X(_04396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17563_ (.A1(_09627_),
    .A2(_09687_),
    .B1(\design_top.core0.REG1[5][27] ),
    .B2(_09690_),
    .X(_04395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17564_ (.A(_09686_),
    .X(_09691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17565_ (.A(_09689_),
    .X(_09692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17566_ (.A1(_09628_),
    .A2(_09691_),
    .B1(\design_top.core0.REG1[5][26] ),
    .B2(_09692_),
    .X(_04394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17567_ (.A1(_09631_),
    .A2(_09691_),
    .B1(\design_top.core0.REG1[5][25] ),
    .B2(_09692_),
    .X(_04393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17568_ (.A1(_09632_),
    .A2(_09691_),
    .B1(\design_top.core0.REG1[5][24] ),
    .B2(_09692_),
    .X(_04392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17569_ (.A1(_09633_),
    .A2(_09691_),
    .B1(\design_top.core0.REG1[5][23] ),
    .B2(_09692_),
    .X(_04391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17570_ (.A1(_09634_),
    .A2(_09691_),
    .B1(\design_top.core0.REG1[5][22] ),
    .B2(_09692_),
    .X(_04390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17571_ (.A(_09686_),
    .X(_09693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17572_ (.A(_09689_),
    .X(_09694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17573_ (.A1(_09635_),
    .A2(_09693_),
    .B1(\design_top.core0.REG1[5][21] ),
    .B2(_09694_),
    .X(_04389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17574_ (.A1(_09638_),
    .A2(_09693_),
    .B1(\design_top.core0.REG1[5][20] ),
    .B2(_09694_),
    .X(_04388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17575_ (.A1(_09639_),
    .A2(_09693_),
    .B1(\design_top.core0.REG1[5][19] ),
    .B2(_09694_),
    .X(_04387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17576_ (.A1(_09640_),
    .A2(_09693_),
    .B1(\design_top.core0.REG1[5][18] ),
    .B2(_09694_),
    .X(_04386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17577_ (.A1(_09641_),
    .A2(_09693_),
    .B1(\design_top.core0.REG1[5][17] ),
    .B2(_09694_),
    .X(_04385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17578_ (.A(_09685_),
    .X(_09695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17579_ (.A(_09688_),
    .X(_09696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17580_ (.A1(_09642_),
    .A2(_09695_),
    .B1(\design_top.core0.REG1[5][16] ),
    .B2(_09696_),
    .X(_04384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17581_ (.A1(_09645_),
    .A2(_09695_),
    .B1(\design_top.core0.REG1[5][15] ),
    .B2(_09696_),
    .X(_04383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17582_ (.A1(_09646_),
    .A2(_09695_),
    .B1(\design_top.core0.REG1[5][14] ),
    .B2(_09696_),
    .X(_04382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17583_ (.A1(\design_top.core0.REG1[5][13] ),
    .A2(_09686_),
    .B1(_09598_),
    .B2(_09689_),
    .X(_04381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17584_ (.A1(_09647_),
    .A2(_09695_),
    .B1(\design_top.core0.REG1[5][12] ),
    .B2(_09696_),
    .X(_04380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17585_ (.A1(_09648_),
    .A2(_09695_),
    .B1(\design_top.core0.REG1[5][11] ),
    .B2(_09696_),
    .X(_04379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17586_ (.A(_09685_),
    .X(_09697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17587_ (.A(_09688_),
    .X(_09698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17588_ (.A1(_09649_),
    .A2(_09697_),
    .B1(\design_top.core0.REG1[5][10] ),
    .B2(_09698_),
    .X(_04378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17589_ (.A1(_09652_),
    .A2(_09697_),
    .B1(\design_top.core0.REG1[5][9] ),
    .B2(_09698_),
    .X(_04377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17590_ (.A1(_09653_),
    .A2(_09697_),
    .B1(\design_top.core0.REG1[5][8] ),
    .B2(_09698_),
    .X(_04376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17591_ (.A1(_09654_),
    .A2(_09697_),
    .B1(\design_top.core0.REG1[5][7] ),
    .B2(_09698_),
    .X(_04375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17592_ (.A1(_09655_),
    .A2(_09697_),
    .B1(\design_top.core0.REG1[5][6] ),
    .B2(_09698_),
    .X(_04374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17593_ (.A(_09685_),
    .X(_09699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17594_ (.A(_09688_),
    .X(_09700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17595_ (.A1(_09656_),
    .A2(_09699_),
    .B1(\design_top.core0.REG1[5][5] ),
    .B2(_09700_),
    .X(_04373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17596_ (.A1(_09659_),
    .A2(_09699_),
    .B1(\design_top.core0.REG1[5][4] ),
    .B2(_09700_),
    .X(_04372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17597_ (.A1(_09660_),
    .A2(_09699_),
    .B1(\design_top.core0.REG1[5][3] ),
    .B2(_09700_),
    .X(_04371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17598_ (.A1(_09661_),
    .A2(_09699_),
    .B1(\design_top.core0.REG1[5][2] ),
    .B2(_09700_),
    .X(_04370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17599_ (.A1(_09662_),
    .A2(_09699_),
    .B1(\design_top.core0.REG1[5][1] ),
    .B2(_09700_),
    .X(_04369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17600_ (.A1(_09663_),
    .A2(_09686_),
    .B1(\design_top.core0.REG1[5][0] ),
    .B2(_09689_),
    .X(_04368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17601_ (.A(_08789_),
    .X(_09701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _17602_ (.A(_09701_),
    .B(_09348_),
    .X(_09702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17603_ (.A(_09702_),
    .X(_09703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17604_ (.A(_09703_),
    .X(_09704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17605_ (.A(_09702_),
    .Y(_09705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17606_ (.A(_09705_),
    .X(_09706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17607_ (.A(_09706_),
    .X(_09707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17608_ (.A1(_09617_),
    .A2(_09704_),
    .B1(\design_top.core0.REG1[4][31] ),
    .B2(_09707_),
    .X(_04367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17609_ (.A1(_09624_),
    .A2(_09704_),
    .B1(\design_top.core0.REG1[4][30] ),
    .B2(_09707_),
    .X(_04366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17610_ (.A1(_09625_),
    .A2(_09704_),
    .B1(\design_top.core0.REG1[4][29] ),
    .B2(_09707_),
    .X(_04365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17611_ (.A1(_09626_),
    .A2(_09704_),
    .B1(\design_top.core0.REG1[4][28] ),
    .B2(_09707_),
    .X(_04364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17612_ (.A1(_09627_),
    .A2(_09704_),
    .B1(\design_top.core0.REG1[4][27] ),
    .B2(_09707_),
    .X(_04363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17613_ (.A(_09703_),
    .X(_09708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17614_ (.A(_09706_),
    .X(_09709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17615_ (.A1(_09628_),
    .A2(_09708_),
    .B1(\design_top.core0.REG1[4][26] ),
    .B2(_09709_),
    .X(_04362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17616_ (.A1(_09631_),
    .A2(_09708_),
    .B1(\design_top.core0.REG1[4][25] ),
    .B2(_09709_),
    .X(_04361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17617_ (.A1(_09632_),
    .A2(_09708_),
    .B1(\design_top.core0.REG1[4][24] ),
    .B2(_09709_),
    .X(_04360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17618_ (.A1(_09633_),
    .A2(_09708_),
    .B1(\design_top.core0.REG1[4][23] ),
    .B2(_09709_),
    .X(_04359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17619_ (.A1(_09634_),
    .A2(_09708_),
    .B1(\design_top.core0.REG1[4][22] ),
    .B2(_09709_),
    .X(_04358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17620_ (.A(_09703_),
    .X(_09710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17621_ (.A(_09706_),
    .X(_09711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17622_ (.A1(_09635_),
    .A2(_09710_),
    .B1(\design_top.core0.REG1[4][21] ),
    .B2(_09711_),
    .X(_04357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17623_ (.A1(_09638_),
    .A2(_09710_),
    .B1(\design_top.core0.REG1[4][20] ),
    .B2(_09711_),
    .X(_04356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17624_ (.A1(_09639_),
    .A2(_09710_),
    .B1(\design_top.core0.REG1[4][19] ),
    .B2(_09711_),
    .X(_04355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17625_ (.A1(_09640_),
    .A2(_09710_),
    .B1(\design_top.core0.REG1[4][18] ),
    .B2(_09711_),
    .X(_04354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17626_ (.A1(_09641_),
    .A2(_09710_),
    .B1(\design_top.core0.REG1[4][17] ),
    .B2(_09711_),
    .X(_04353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17627_ (.A(_09702_),
    .X(_09712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17628_ (.A(_09705_),
    .X(_09713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17629_ (.A1(_09642_),
    .A2(_09712_),
    .B1(\design_top.core0.REG1[4][16] ),
    .B2(_09713_),
    .X(_04352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17630_ (.A1(_09645_),
    .A2(_09712_),
    .B1(\design_top.core0.REG1[4][15] ),
    .B2(_09713_),
    .X(_04351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17631_ (.A1(_09646_),
    .A2(_09712_),
    .B1(\design_top.core0.REG1[4][14] ),
    .B2(_09713_),
    .X(_04350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17632_ (.A(_00045_),
    .X(_09714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17633_ (.A1(\design_top.core0.REG1[4][13] ),
    .A2(_09703_),
    .B1(_09714_),
    .B2(_09706_),
    .X(_04349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17634_ (.A1(_09647_),
    .A2(_09712_),
    .B1(\design_top.core0.REG1[4][12] ),
    .B2(_09713_),
    .X(_04348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17635_ (.A1(_09648_),
    .A2(_09712_),
    .B1(\design_top.core0.REG1[4][11] ),
    .B2(_09713_),
    .X(_04347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17636_ (.A(_09702_),
    .X(_09715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17637_ (.A(_09705_),
    .X(_09716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17638_ (.A1(_09649_),
    .A2(_09715_),
    .B1(\design_top.core0.REG1[4][10] ),
    .B2(_09716_),
    .X(_04346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17639_ (.A1(_09652_),
    .A2(_09715_),
    .B1(\design_top.core0.REG1[4][9] ),
    .B2(_09716_),
    .X(_04345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17640_ (.A1(_09653_),
    .A2(_09715_),
    .B1(\design_top.core0.REG1[4][8] ),
    .B2(_09716_),
    .X(_04344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17641_ (.A1(_09654_),
    .A2(_09715_),
    .B1(\design_top.core0.REG1[4][7] ),
    .B2(_09716_),
    .X(_04343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17642_ (.A1(_09655_),
    .A2(_09715_),
    .B1(\design_top.core0.REG1[4][6] ),
    .B2(_09716_),
    .X(_04342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17643_ (.A(_09702_),
    .X(_09717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17644_ (.A(_09705_),
    .X(_09718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17645_ (.A1(_09656_),
    .A2(_09717_),
    .B1(\design_top.core0.REG1[4][5] ),
    .B2(_09718_),
    .X(_04341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17646_ (.A1(_09659_),
    .A2(_09717_),
    .B1(\design_top.core0.REG1[4][4] ),
    .B2(_09718_),
    .X(_04340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17647_ (.A1(_09660_),
    .A2(_09717_),
    .B1(\design_top.core0.REG1[4][3] ),
    .B2(_09718_),
    .X(_04339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17648_ (.A1(_09661_),
    .A2(_09717_),
    .B1(\design_top.core0.REG1[4][2] ),
    .B2(_09718_),
    .X(_04338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17649_ (.A1(_09662_),
    .A2(_09717_),
    .B1(\design_top.core0.REG1[4][1] ),
    .B2(_09718_),
    .X(_04337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17650_ (.A1(_09663_),
    .A2(_09703_),
    .B1(\design_top.core0.REG1[4][0] ),
    .B2(_09706_),
    .X(_04336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _17651_ (.A(_09701_),
    .B(_09367_),
    .X(_09719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17652_ (.A(_09719_),
    .X(_09720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17653_ (.A(_09720_),
    .X(_09721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17654_ (.A(_09719_),
    .Y(_09722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17655_ (.A(_09722_),
    .X(_09723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17656_ (.A(_09723_),
    .X(_09724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17657_ (.A1(_09617_),
    .A2(_09721_),
    .B1(\design_top.core0.REG1[3][31] ),
    .B2(_09724_),
    .X(_04335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17658_ (.A1(_09624_),
    .A2(_09721_),
    .B1(\design_top.core0.REG1[3][30] ),
    .B2(_09724_),
    .X(_04334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17659_ (.A1(_09625_),
    .A2(_09721_),
    .B1(\design_top.core0.REG1[3][29] ),
    .B2(_09724_),
    .X(_04333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17660_ (.A1(_09626_),
    .A2(_09721_),
    .B1(\design_top.core0.REG1[3][28] ),
    .B2(_09724_),
    .X(_04332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17661_ (.A1(_09627_),
    .A2(_09721_),
    .B1(\design_top.core0.REG1[3][27] ),
    .B2(_09724_),
    .X(_04331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17662_ (.A(_09720_),
    .X(_09725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17663_ (.A(_09723_),
    .X(_09726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17664_ (.A1(_09628_),
    .A2(_09725_),
    .B1(\design_top.core0.REG1[3][26] ),
    .B2(_09726_),
    .X(_04330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17665_ (.A1(_09631_),
    .A2(_09725_),
    .B1(\design_top.core0.REG1[3][25] ),
    .B2(_09726_),
    .X(_04329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17666_ (.A1(_09632_),
    .A2(_09725_),
    .B1(\design_top.core0.REG1[3][24] ),
    .B2(_09726_),
    .X(_04328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17667_ (.A1(_09633_),
    .A2(_09725_),
    .B1(\design_top.core0.REG1[3][23] ),
    .B2(_09726_),
    .X(_04327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17668_ (.A1(_09634_),
    .A2(_09725_),
    .B1(\design_top.core0.REG1[3][22] ),
    .B2(_09726_),
    .X(_04326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17669_ (.A(_09720_),
    .X(_09727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17670_ (.A(_09723_),
    .X(_09728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17671_ (.A1(_09635_),
    .A2(_09727_),
    .B1(\design_top.core0.REG1[3][21] ),
    .B2(_09728_),
    .X(_04325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17672_ (.A1(_09638_),
    .A2(_09727_),
    .B1(\design_top.core0.REG1[3][20] ),
    .B2(_09728_),
    .X(_04324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17673_ (.A1(_09639_),
    .A2(_09727_),
    .B1(\design_top.core0.REG1[3][19] ),
    .B2(_09728_),
    .X(_04323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17674_ (.A1(_09640_),
    .A2(_09727_),
    .B1(\design_top.core0.REG1[3][18] ),
    .B2(_09728_),
    .X(_04322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17675_ (.A1(_09641_),
    .A2(_09727_),
    .B1(\design_top.core0.REG1[3][17] ),
    .B2(_09728_),
    .X(_04321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17676_ (.A(_09719_),
    .X(_09729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17677_ (.A(_09722_),
    .X(_09730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17678_ (.A1(_09642_),
    .A2(_09729_),
    .B1(\design_top.core0.REG1[3][16] ),
    .B2(_09730_),
    .X(_04320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17679_ (.A1(_09645_),
    .A2(_09729_),
    .B1(\design_top.core0.REG1[3][15] ),
    .B2(_09730_),
    .X(_04319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17680_ (.A1(_09646_),
    .A2(_09729_),
    .B1(\design_top.core0.REG1[3][14] ),
    .B2(_09730_),
    .X(_04318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17681_ (.A1(\design_top.core0.REG1[3][13] ),
    .A2(_09720_),
    .B1(_09714_),
    .B2(_09723_),
    .X(_04317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17682_ (.A1(_09647_),
    .A2(_09729_),
    .B1(\design_top.core0.REG1[3][12] ),
    .B2(_09730_),
    .X(_04316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17683_ (.A1(_09648_),
    .A2(_09729_),
    .B1(\design_top.core0.REG1[3][11] ),
    .B2(_09730_),
    .X(_04315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17684_ (.A(_09719_),
    .X(_09731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17685_ (.A(_09722_),
    .X(_09732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17686_ (.A1(_09649_),
    .A2(_09731_),
    .B1(\design_top.core0.REG1[3][10] ),
    .B2(_09732_),
    .X(_04314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17687_ (.A1(_09652_),
    .A2(_09731_),
    .B1(\design_top.core0.REG1[3][9] ),
    .B2(_09732_),
    .X(_04313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17688_ (.A1(_09653_),
    .A2(_09731_),
    .B1(\design_top.core0.REG1[3][8] ),
    .B2(_09732_),
    .X(_04312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17689_ (.A1(_09654_),
    .A2(_09731_),
    .B1(\design_top.core0.REG1[3][7] ),
    .B2(_09732_),
    .X(_04311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17690_ (.A1(_09655_),
    .A2(_09731_),
    .B1(\design_top.core0.REG1[3][6] ),
    .B2(_09732_),
    .X(_04310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17691_ (.A(_09719_),
    .X(_09733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17692_ (.A(_09722_),
    .X(_09734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17693_ (.A1(_09656_),
    .A2(_09733_),
    .B1(\design_top.core0.REG1[3][5] ),
    .B2(_09734_),
    .X(_04309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17694_ (.A1(_09659_),
    .A2(_09733_),
    .B1(\design_top.core0.REG1[3][4] ),
    .B2(_09734_),
    .X(_04308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17695_ (.A1(_09660_),
    .A2(_09733_),
    .B1(\design_top.core0.REG1[3][3] ),
    .B2(_09734_),
    .X(_04307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17696_ (.A1(_09661_),
    .A2(_09733_),
    .B1(\design_top.core0.REG1[3][2] ),
    .B2(_09734_),
    .X(_04306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17697_ (.A1(_09662_),
    .A2(_09733_),
    .B1(\design_top.core0.REG1[3][1] ),
    .B2(_09734_),
    .X(_04305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17698_ (.A1(_09663_),
    .A2(_09720_),
    .B1(\design_top.core0.REG1[3][0] ),
    .B2(_09723_),
    .X(_04304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _17699_ (.A(_09701_),
    .B(_09414_),
    .X(_09735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17700_ (.A(_09735_),
    .X(_09736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17701_ (.A(_09736_),
    .X(_09737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17702_ (.A(_09735_),
    .Y(_09738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17703_ (.A(_09738_),
    .X(_09739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17704_ (.A(_09739_),
    .X(_09740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17705_ (.A1(_08800_),
    .A2(_09737_),
    .B1(\design_top.core0.REG1[2][31] ),
    .B2(_09740_),
    .X(_04303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17706_ (.A1(_08802_),
    .A2(_09737_),
    .B1(\design_top.core0.REG1[2][30] ),
    .B2(_09740_),
    .X(_04302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17707_ (.A1(_08804_),
    .A2(_09737_),
    .B1(\design_top.core0.REG1[2][29] ),
    .B2(_09740_),
    .X(_04301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17708_ (.A1(_08806_),
    .A2(_09737_),
    .B1(\design_top.core0.REG1[2][28] ),
    .B2(_09740_),
    .X(_04300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17709_ (.A1(_08809_),
    .A2(_09737_),
    .B1(\design_top.core0.REG1[2][27] ),
    .B2(_09740_),
    .X(_04299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17710_ (.A(_09736_),
    .X(_09741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17711_ (.A(_09739_),
    .X(_09742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17712_ (.A1(_08813_),
    .A2(_09741_),
    .B1(\design_top.core0.REG1[2][26] ),
    .B2(_09742_),
    .X(_04298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17713_ (.A1(_08815_),
    .A2(_09741_),
    .B1(\design_top.core0.REG1[2][25] ),
    .B2(_09742_),
    .X(_04297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17714_ (.A1(_08817_),
    .A2(_09741_),
    .B1(\design_top.core0.REG1[2][24] ),
    .B2(_09742_),
    .X(_04296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17715_ (.A1(_08819_),
    .A2(_09741_),
    .B1(\design_top.core0.REG1[2][23] ),
    .B2(_09742_),
    .X(_04295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17716_ (.A1(_08822_),
    .A2(_09741_),
    .B1(\design_top.core0.REG1[2][22] ),
    .B2(_09742_),
    .X(_04294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17717_ (.A(_09736_),
    .X(_09743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17718_ (.A(_09739_),
    .X(_09744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17719_ (.A1(_08826_),
    .A2(_09743_),
    .B1(\design_top.core0.REG1[2][21] ),
    .B2(_09744_),
    .X(_04293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17720_ (.A1(_08828_),
    .A2(_09743_),
    .B1(\design_top.core0.REG1[2][20] ),
    .B2(_09744_),
    .X(_04292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17721_ (.A1(_08830_),
    .A2(_09743_),
    .B1(\design_top.core0.REG1[2][19] ),
    .B2(_09744_),
    .X(_04291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17722_ (.A1(_08832_),
    .A2(_09743_),
    .B1(\design_top.core0.REG1[2][18] ),
    .B2(_09744_),
    .X(_04290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17723_ (.A1(_08835_),
    .A2(_09743_),
    .B1(\design_top.core0.REG1[2][17] ),
    .B2(_09744_),
    .X(_04289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17724_ (.A(_09735_),
    .X(_09745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17725_ (.A(_09738_),
    .X(_09746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17726_ (.A1(_08839_),
    .A2(_09745_),
    .B1(\design_top.core0.REG1[2][16] ),
    .B2(_09746_),
    .X(_04288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17727_ (.A1(_08841_),
    .A2(_09745_),
    .B1(\design_top.core0.REG1[2][15] ),
    .B2(_09746_),
    .X(_04287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17728_ (.A1(_08843_),
    .A2(_09745_),
    .B1(\design_top.core0.REG1[2][14] ),
    .B2(_09746_),
    .X(_04286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17729_ (.A1(\design_top.core0.REG1[2][13] ),
    .A2(_09736_),
    .B1(_09714_),
    .B2(_09739_),
    .X(_04285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17730_ (.A1(_08846_),
    .A2(_09745_),
    .B1(\design_top.core0.REG1[2][12] ),
    .B2(_09746_),
    .X(_04284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17731_ (.A1(_08849_),
    .A2(_09745_),
    .B1(\design_top.core0.REG1[2][11] ),
    .B2(_09746_),
    .X(_04283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17732_ (.A(_09735_),
    .X(_09747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17733_ (.A(_09738_),
    .X(_09748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17734_ (.A1(_08853_),
    .A2(_09747_),
    .B1(\design_top.core0.REG1[2][10] ),
    .B2(_09748_),
    .X(_04282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17735_ (.A1(_08855_),
    .A2(_09747_),
    .B1(\design_top.core0.REG1[2][9] ),
    .B2(_09748_),
    .X(_04281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17736_ (.A1(_08857_),
    .A2(_09747_),
    .B1(\design_top.core0.REG1[2][8] ),
    .B2(_09748_),
    .X(_04280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17737_ (.A1(_08859_),
    .A2(_09747_),
    .B1(\design_top.core0.REG1[2][7] ),
    .B2(_09748_),
    .X(_04279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17738_ (.A1(_08862_),
    .A2(_09747_),
    .B1(\design_top.core0.REG1[2][6] ),
    .B2(_09748_),
    .X(_04278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17739_ (.A(_09735_),
    .X(_09749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17740_ (.A(_09738_),
    .X(_09750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17741_ (.A1(_08866_),
    .A2(_09749_),
    .B1(\design_top.core0.REG1[2][5] ),
    .B2(_09750_),
    .X(_04277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17742_ (.A1(_08868_),
    .A2(_09749_),
    .B1(\design_top.core0.REG1[2][4] ),
    .B2(_09750_),
    .X(_04276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17743_ (.A1(_08870_),
    .A2(_09749_),
    .B1(\design_top.core0.REG1[2][3] ),
    .B2(_09750_),
    .X(_04275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17744_ (.A1(_08872_),
    .A2(_09749_),
    .B1(\design_top.core0.REG1[2][2] ),
    .B2(_09750_),
    .X(_04274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17745_ (.A1(_08874_),
    .A2(_09749_),
    .B1(\design_top.core0.REG1[2][1] ),
    .B2(_09750_),
    .X(_04273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17746_ (.A1(_08876_),
    .A2(_09736_),
    .B1(\design_top.core0.REG1[2][0] ),
    .B2(_09739_),
    .X(_04272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _17747_ (.A(_09701_),
    .B(_09431_),
    .X(_09751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17748_ (.A(_09751_),
    .X(_09752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17749_ (.A(_09752_),
    .X(_09753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17750_ (.A(_09751_),
    .Y(_09754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17751_ (.A(_09754_),
    .X(_09755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17752_ (.A(_09755_),
    .X(_09756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17753_ (.A1(_08800_),
    .A2(_09753_),
    .B1(\design_top.core0.REG1[1][31] ),
    .B2(_09756_),
    .X(_04271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17754_ (.A1(_08802_),
    .A2(_09753_),
    .B1(\design_top.core0.REG1[1][30] ),
    .B2(_09756_),
    .X(_04270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17755_ (.A1(_08804_),
    .A2(_09753_),
    .B1(\design_top.core0.REG1[1][29] ),
    .B2(_09756_),
    .X(_04269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17756_ (.A1(_08806_),
    .A2(_09753_),
    .B1(\design_top.core0.REG1[1][28] ),
    .B2(_09756_),
    .X(_04268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17757_ (.A1(_08809_),
    .A2(_09753_),
    .B1(\design_top.core0.REG1[1][27] ),
    .B2(_09756_),
    .X(_04267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17758_ (.A(_09752_),
    .X(_09757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17759_ (.A(_09755_),
    .X(_09758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17760_ (.A1(_08813_),
    .A2(_09757_),
    .B1(\design_top.core0.REG1[1][26] ),
    .B2(_09758_),
    .X(_04266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17761_ (.A1(_08815_),
    .A2(_09757_),
    .B1(\design_top.core0.REG1[1][25] ),
    .B2(_09758_),
    .X(_04265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17762_ (.A1(_08817_),
    .A2(_09757_),
    .B1(\design_top.core0.REG1[1][24] ),
    .B2(_09758_),
    .X(_04264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17763_ (.A1(_08819_),
    .A2(_09757_),
    .B1(\design_top.core0.REG1[1][23] ),
    .B2(_09758_),
    .X(_04263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17764_ (.A1(_08822_),
    .A2(_09757_),
    .B1(\design_top.core0.REG1[1][22] ),
    .B2(_09758_),
    .X(_04262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17765_ (.A(_09752_),
    .X(_09759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17766_ (.A(_09755_),
    .X(_09760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17767_ (.A1(_08826_),
    .A2(_09759_),
    .B1(\design_top.core0.REG1[1][21] ),
    .B2(_09760_),
    .X(_04261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17768_ (.A1(_08828_),
    .A2(_09759_),
    .B1(\design_top.core0.REG1[1][20] ),
    .B2(_09760_),
    .X(_04260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17769_ (.A1(_08830_),
    .A2(_09759_),
    .B1(\design_top.core0.REG1[1][19] ),
    .B2(_09760_),
    .X(_04259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17770_ (.A1(_08832_),
    .A2(_09759_),
    .B1(\design_top.core0.REG1[1][18] ),
    .B2(_09760_),
    .X(_04258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17771_ (.A1(_08835_),
    .A2(_09759_),
    .B1(\design_top.core0.REG1[1][17] ),
    .B2(_09760_),
    .X(_04257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17772_ (.A(_09751_),
    .X(_09761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17773_ (.A(_09754_),
    .X(_09762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17774_ (.A1(_08839_),
    .A2(_09761_),
    .B1(\design_top.core0.REG1[1][16] ),
    .B2(_09762_),
    .X(_04256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17775_ (.A1(_08841_),
    .A2(_09761_),
    .B1(\design_top.core0.REG1[1][15] ),
    .B2(_09762_),
    .X(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17776_ (.A1(_08843_),
    .A2(_09761_),
    .B1(\design_top.core0.REG1[1][14] ),
    .B2(_09762_),
    .X(_04254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17777_ (.A1(\design_top.core0.REG1[1][13] ),
    .A2(_09752_),
    .B1(_09714_),
    .B2(_09755_),
    .X(_04253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17778_ (.A1(_08846_),
    .A2(_09761_),
    .B1(\design_top.core0.REG1[1][12] ),
    .B2(_09762_),
    .X(_04252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17779_ (.A1(_08849_),
    .A2(_09761_),
    .B1(\design_top.core0.REG1[1][11] ),
    .B2(_09762_),
    .X(_04251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17780_ (.A(_09751_),
    .X(_09763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17781_ (.A(_09754_),
    .X(_09764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17782_ (.A1(_08853_),
    .A2(_09763_),
    .B1(\design_top.core0.REG1[1][10] ),
    .B2(_09764_),
    .X(_04250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17783_ (.A1(_08855_),
    .A2(_09763_),
    .B1(\design_top.core0.REG1[1][9] ),
    .B2(_09764_),
    .X(_04249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17784_ (.A1(_08857_),
    .A2(_09763_),
    .B1(\design_top.core0.REG1[1][8] ),
    .B2(_09764_),
    .X(_04248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17785_ (.A1(_08859_),
    .A2(_09763_),
    .B1(\design_top.core0.REG1[1][7] ),
    .B2(_09764_),
    .X(_04247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17786_ (.A1(_08862_),
    .A2(_09763_),
    .B1(\design_top.core0.REG1[1][6] ),
    .B2(_09764_),
    .X(_04246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17787_ (.A(_09751_),
    .X(_09765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17788_ (.A(_09754_),
    .X(_09766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17789_ (.A1(_08866_),
    .A2(_09765_),
    .B1(\design_top.core0.REG1[1][5] ),
    .B2(_09766_),
    .X(_04245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17790_ (.A1(_08868_),
    .A2(_09765_),
    .B1(\design_top.core0.REG1[1][4] ),
    .B2(_09766_),
    .X(_04244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17791_ (.A1(_08870_),
    .A2(_09765_),
    .B1(\design_top.core0.REG1[1][3] ),
    .B2(_09766_),
    .X(_04243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17792_ (.A1(_08872_),
    .A2(_09765_),
    .B1(\design_top.core0.REG1[1][2] ),
    .B2(_09766_),
    .X(_04242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17793_ (.A1(_08874_),
    .A2(_09765_),
    .B1(\design_top.core0.REG1[1][1] ),
    .B2(_09766_),
    .X(_04241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17794_ (.A1(_08876_),
    .A2(_09752_),
    .B1(\design_top.core0.REG1[1][0] ),
    .B2(_09755_),
    .X(_04240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _17795_ (.A(_09701_),
    .B(_09448_),
    .X(_09767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17796_ (.A(_09767_),
    .X(_09768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17797_ (.A(_09768_),
    .X(_09769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17798_ (.A(_09767_),
    .Y(_09770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17799_ (.A(_09770_),
    .X(_09771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17800_ (.A(_09771_),
    .X(_09772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17801_ (.A1(_08800_),
    .A2(_09769_),
    .B1(\design_top.core0.REG1[15][31] ),
    .B2(_09772_),
    .X(_04239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17802_ (.A1(_08802_),
    .A2(_09769_),
    .B1(\design_top.core0.REG1[15][30] ),
    .B2(_09772_),
    .X(_04238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17803_ (.A1(_08804_),
    .A2(_09769_),
    .B1(\design_top.core0.REG1[15][29] ),
    .B2(_09772_),
    .X(_04237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17804_ (.A1(_08806_),
    .A2(_09769_),
    .B1(\design_top.core0.REG1[15][28] ),
    .B2(_09772_),
    .X(_04236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17805_ (.A1(_08809_),
    .A2(_09769_),
    .B1(\design_top.core0.REG1[15][27] ),
    .B2(_09772_),
    .X(_04235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17806_ (.A(_09768_),
    .X(_09773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17807_ (.A(_09771_),
    .X(_09774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17808_ (.A1(_08813_),
    .A2(_09773_),
    .B1(\design_top.core0.REG1[15][26] ),
    .B2(_09774_),
    .X(_04234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17809_ (.A1(_08815_),
    .A2(_09773_),
    .B1(\design_top.core0.REG1[15][25] ),
    .B2(_09774_),
    .X(_04233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17810_ (.A1(_08817_),
    .A2(_09773_),
    .B1(\design_top.core0.REG1[15][24] ),
    .B2(_09774_),
    .X(_04232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17811_ (.A1(_08819_),
    .A2(_09773_),
    .B1(\design_top.core0.REG1[15][23] ),
    .B2(_09774_),
    .X(_04231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17812_ (.A1(_08822_),
    .A2(_09773_),
    .B1(\design_top.core0.REG1[15][22] ),
    .B2(_09774_),
    .X(_04230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17813_ (.A(_09768_),
    .X(_09775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17814_ (.A(_09771_),
    .X(_09776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17815_ (.A1(_08826_),
    .A2(_09775_),
    .B1(\design_top.core0.REG1[15][21] ),
    .B2(_09776_),
    .X(_04229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17816_ (.A1(_08828_),
    .A2(_09775_),
    .B1(\design_top.core0.REG1[15][20] ),
    .B2(_09776_),
    .X(_04228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17817_ (.A1(_08830_),
    .A2(_09775_),
    .B1(\design_top.core0.REG1[15][19] ),
    .B2(_09776_),
    .X(_04227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17818_ (.A1(_08832_),
    .A2(_09775_),
    .B1(\design_top.core0.REG1[15][18] ),
    .B2(_09776_),
    .X(_04226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17819_ (.A1(_08835_),
    .A2(_09775_),
    .B1(\design_top.core0.REG1[15][17] ),
    .B2(_09776_),
    .X(_04225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17820_ (.A(_09767_),
    .X(_09777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17821_ (.A(_09770_),
    .X(_09778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17822_ (.A1(_08839_),
    .A2(_09777_),
    .B1(\design_top.core0.REG1[15][16] ),
    .B2(_09778_),
    .X(_04224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17823_ (.A1(_08841_),
    .A2(_09777_),
    .B1(\design_top.core0.REG1[15][15] ),
    .B2(_09778_),
    .X(_04223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17824_ (.A1(_08843_),
    .A2(_09777_),
    .B1(\design_top.core0.REG1[15][14] ),
    .B2(_09778_),
    .X(_04222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17825_ (.A1(\design_top.core0.REG1[15][13] ),
    .A2(_09768_),
    .B1(_09714_),
    .B2(_09771_),
    .X(_04221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17826_ (.A1(_08846_),
    .A2(_09777_),
    .B1(\design_top.core0.REG1[15][12] ),
    .B2(_09778_),
    .X(_04220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17827_ (.A1(_08849_),
    .A2(_09777_),
    .B1(\design_top.core0.REG1[15][11] ),
    .B2(_09778_),
    .X(_04219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17828_ (.A(_09767_),
    .X(_09779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17829_ (.A(_09770_),
    .X(_09780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17830_ (.A1(_08853_),
    .A2(_09779_),
    .B1(\design_top.core0.REG1[15][10] ),
    .B2(_09780_),
    .X(_04218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17831_ (.A1(_08855_),
    .A2(_09779_),
    .B1(\design_top.core0.REG1[15][9] ),
    .B2(_09780_),
    .X(_04217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17832_ (.A1(_08857_),
    .A2(_09779_),
    .B1(\design_top.core0.REG1[15][8] ),
    .B2(_09780_),
    .X(_04216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17833_ (.A1(_08859_),
    .A2(_09779_),
    .B1(\design_top.core0.REG1[15][7] ),
    .B2(_09780_),
    .X(_04215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17834_ (.A1(_08862_),
    .A2(_09779_),
    .B1(\design_top.core0.REG1[15][6] ),
    .B2(_09780_),
    .X(_04214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17835_ (.A(_09767_),
    .X(_09781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17836_ (.A(_09770_),
    .X(_09782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17837_ (.A1(_08866_),
    .A2(_09781_),
    .B1(\design_top.core0.REG1[15][5] ),
    .B2(_09782_),
    .X(_04213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17838_ (.A1(_08868_),
    .A2(_09781_),
    .B1(\design_top.core0.REG1[15][4] ),
    .B2(_09782_),
    .X(_04212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17839_ (.A1(_08870_),
    .A2(_09781_),
    .B1(\design_top.core0.REG1[15][3] ),
    .B2(_09782_),
    .X(_04211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17840_ (.A1(_08872_),
    .A2(_09781_),
    .B1(\design_top.core0.REG1[15][2] ),
    .B2(_09782_),
    .X(_04210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17841_ (.A1(_08874_),
    .A2(_09781_),
    .B1(\design_top.core0.REG1[15][1] ),
    .B2(_09782_),
    .X(_04209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17842_ (.A1(_08876_),
    .A2(_09768_),
    .B1(\design_top.core0.REG1[15][0] ),
    .B2(_09771_),
    .X(_04208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17843_ (.A1(_10798_),
    .A2(_08169_),
    .B1(_08238_),
    .B2(_09680_),
    .X(_09783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17844_ (.A(_09783_),
    .Y(_09784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17845_ (.A(_09784_),
    .X(_09785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17846_ (.A(_09783_),
    .X(_09786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17847_ (.A1(_00628_),
    .A2(_09785_),
    .B1(\design_top.MEM[60][7] ),
    .B2(_09786_),
    .X(_04207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17848_ (.A1(_00627_),
    .A2(_09785_),
    .B1(\design_top.MEM[60][6] ),
    .B2(_09786_),
    .X(_04206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17849_ (.A1(_00626_),
    .A2(_09785_),
    .B1(\design_top.MEM[60][5] ),
    .B2(_09786_),
    .X(_04205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17850_ (.A1(_00625_),
    .A2(_09785_),
    .B1(\design_top.MEM[60][4] ),
    .B2(_09786_),
    .X(_04204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17851_ (.A1(_00624_),
    .A2(_09785_),
    .B1(\design_top.MEM[60][3] ),
    .B2(_09786_),
    .X(_04203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17852_ (.A1(_00623_),
    .A2(_09784_),
    .B1(\design_top.MEM[60][2] ),
    .B2(_09783_),
    .X(_04202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17853_ (.A1(_00622_),
    .A2(_09784_),
    .B1(\design_top.MEM[60][1] ),
    .B2(_09783_),
    .X(_04201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17854_ (.A1(_00621_),
    .A2(_09784_),
    .B1(\design_top.MEM[60][0] ),
    .B2(_09783_),
    .X(_04200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17855_ (.A1(_09050_),
    .A2(_07867_),
    .B1(_08252_),
    .B2(_09680_),
    .X(_09787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17856_ (.A(_09787_),
    .Y(_09788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17857_ (.A(_09788_),
    .X(_09789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17858_ (.A(_09787_),
    .X(_09790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17859_ (.A1(_00620_),
    .A2(_09789_),
    .B1(\design_top.MEM[5][7] ),
    .B2(_09790_),
    .X(_04199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17860_ (.A1(_00619_),
    .A2(_09789_),
    .B1(\design_top.MEM[5][6] ),
    .B2(_09790_),
    .X(_04198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17861_ (.A1(_00618_),
    .A2(_09789_),
    .B1(\design_top.MEM[5][5] ),
    .B2(_09790_),
    .X(_04197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17862_ (.A1(_00617_),
    .A2(_09789_),
    .B1(\design_top.MEM[5][4] ),
    .B2(_09790_),
    .X(_04196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17863_ (.A1(_00616_),
    .A2(_09789_),
    .B1(\design_top.MEM[5][3] ),
    .B2(_09790_),
    .X(_04195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17864_ (.A1(_00615_),
    .A2(_09788_),
    .B1(\design_top.MEM[5][2] ),
    .B2(_09787_),
    .X(_04194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17865_ (.A1(_00614_),
    .A2(_09788_),
    .B1(\design_top.MEM[5][1] ),
    .B2(_09787_),
    .X(_04193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17866_ (.A1(_00613_),
    .A2(_09788_),
    .B1(\design_top.MEM[5][0] ),
    .B2(_09787_),
    .X(_04192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17867_ (.A1(_10890_),
    .A2(_08269_),
    .B1(_08265_),
    .B2(_09680_),
    .X(_09791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17868_ (.A(_09791_),
    .Y(_09792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17869_ (.A(_09792_),
    .X(_09793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17870_ (.A(_09791_),
    .X(_09794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17871_ (.A1(_00612_),
    .A2(_09793_),
    .B1(\design_top.MEM[59][7] ),
    .B2(_09794_),
    .X(_04191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17872_ (.A1(_00611_),
    .A2(_09793_),
    .B1(\design_top.MEM[59][6] ),
    .B2(_09794_),
    .X(_04190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17873_ (.A1(_00610_),
    .A2(_09793_),
    .B1(\design_top.MEM[59][5] ),
    .B2(_09794_),
    .X(_04189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17874_ (.A1(_00609_),
    .A2(_09793_),
    .B1(\design_top.MEM[59][4] ),
    .B2(_09794_),
    .X(_04188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17875_ (.A1(_00608_),
    .A2(_09793_),
    .B1(\design_top.MEM[59][3] ),
    .B2(_09794_),
    .X(_04187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17876_ (.A1(_00607_),
    .A2(_09792_),
    .B1(\design_top.MEM[59][2] ),
    .B2(_09791_),
    .X(_04186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17877_ (.A1(_00606_),
    .A2(_09792_),
    .B1(\design_top.MEM[59][1] ),
    .B2(_09791_),
    .X(_04185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17878_ (.A1(_00605_),
    .A2(_09792_),
    .B1(\design_top.MEM[59][0] ),
    .B2(_09791_),
    .X(_04184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17879_ (.A1(_09032_),
    .A2(_08268_),
    .B1(_08281_),
    .B2(_09680_),
    .X(_09795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17880_ (.A(_09795_),
    .Y(_09796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17881_ (.A(_09796_),
    .X(_09797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17882_ (.A(_09795_),
    .X(_09798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17883_ (.A1(_00604_),
    .A2(_09797_),
    .B1(\design_top.MEM[58][7] ),
    .B2(_09798_),
    .X(_04183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17884_ (.A1(_00603_),
    .A2(_09797_),
    .B1(\design_top.MEM[58][6] ),
    .B2(_09798_),
    .X(_04182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17885_ (.A1(_00602_),
    .A2(_09797_),
    .B1(\design_top.MEM[58][5] ),
    .B2(_09798_),
    .X(_04181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17886_ (.A1(_00601_),
    .A2(_09797_),
    .B1(\design_top.MEM[58][4] ),
    .B2(_09798_),
    .X(_04180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17887_ (.A1(_00600_),
    .A2(_09797_),
    .B1(\design_top.MEM[58][3] ),
    .B2(_09798_),
    .X(_04179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17888_ (.A1(_00599_),
    .A2(_09796_),
    .B1(\design_top.MEM[58][2] ),
    .B2(_09795_),
    .X(_04178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17889_ (.A1(_00598_),
    .A2(_09796_),
    .B1(\design_top.MEM[58][1] ),
    .B2(_09795_),
    .X(_04177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17890_ (.A1(_00597_),
    .A2(_09796_),
    .B1(\design_top.MEM[58][0] ),
    .B2(_09795_),
    .X(_04176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17891_ (.A1(_09050_),
    .A2(_08268_),
    .B1(_08295_),
    .B2(_08756_),
    .X(_09799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17892_ (.A(_09799_),
    .Y(_09800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17893_ (.A(_09800_),
    .X(_09801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17894_ (.A(_09799_),
    .X(_09802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17895_ (.A1(_00596_),
    .A2(_09801_),
    .B1(\design_top.MEM[57][7] ),
    .B2(_09802_),
    .X(_04175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17896_ (.A1(_00595_),
    .A2(_09801_),
    .B1(\design_top.MEM[57][6] ),
    .B2(_09802_),
    .X(_04174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17897_ (.A1(_00594_),
    .A2(_09801_),
    .B1(\design_top.MEM[57][5] ),
    .B2(_09802_),
    .X(_04173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17898_ (.A1(_00593_),
    .A2(_09801_),
    .B1(\design_top.MEM[57][4] ),
    .B2(_09802_),
    .X(_04172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17899_ (.A1(_00592_),
    .A2(_09801_),
    .B1(\design_top.MEM[57][3] ),
    .B2(_09802_),
    .X(_04171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17900_ (.A1(_00591_),
    .A2(_09800_),
    .B1(\design_top.MEM[57][2] ),
    .B2(_09799_),
    .X(_04170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17901_ (.A1(_00590_),
    .A2(_09800_),
    .B1(\design_top.MEM[57][1] ),
    .B2(_09799_),
    .X(_04169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17902_ (.A1(_00589_),
    .A2(_09800_),
    .B1(\design_top.MEM[57][0] ),
    .B2(_09799_),
    .X(_04168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17903_ (.A1(_10798_),
    .A2(_08268_),
    .B1(_08308_),
    .B2(_08756_),
    .X(_09803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17904_ (.A(_09803_),
    .Y(_09804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17905_ (.A(_09804_),
    .X(_09805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17906_ (.A(_09803_),
    .X(_09806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17907_ (.A1(_00588_),
    .A2(_09805_),
    .B1(\design_top.MEM[56][7] ),
    .B2(_09806_),
    .X(_04167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17908_ (.A1(_00587_),
    .A2(_09805_),
    .B1(\design_top.MEM[56][6] ),
    .B2(_09806_),
    .X(_04166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17909_ (.A1(_00586_),
    .A2(_09805_),
    .B1(\design_top.MEM[56][5] ),
    .B2(_09806_),
    .X(_04165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17910_ (.A1(_00585_),
    .A2(_09805_),
    .B1(\design_top.MEM[56][4] ),
    .B2(_09806_),
    .X(_04164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17911_ (.A1(_00584_),
    .A2(_09805_),
    .B1(\design_top.MEM[56][3] ),
    .B2(_09806_),
    .X(_04163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17912_ (.A1(_00583_),
    .A2(_09804_),
    .B1(\design_top.MEM[56][2] ),
    .B2(_09803_),
    .X(_04162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17913_ (.A1(_00582_),
    .A2(_09804_),
    .B1(\design_top.MEM[56][1] ),
    .B2(_09803_),
    .X(_04161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17914_ (.A1(_00581_),
    .A2(_09804_),
    .B1(\design_top.MEM[56][0] ),
    .B2(_09803_),
    .X(_04160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _17915_ (.A1(_10890_),
    .A2(_07571_),
    .B1(_07624_),
    .B2(_08756_),
    .X(_09807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17916_ (.A(_09807_),
    .Y(_09808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17917_ (.A(_09808_),
    .X(_09809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17918_ (.A(_09807_),
    .X(_09810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17919_ (.A1(_00580_),
    .A2(_09809_),
    .B1(\design_top.MEM[55][7] ),
    .B2(_09810_),
    .X(_04159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17920_ (.A1(_00579_),
    .A2(_09809_),
    .B1(\design_top.MEM[55][6] ),
    .B2(_09810_),
    .X(_04158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17921_ (.A1(_00578_),
    .A2(_09809_),
    .B1(\design_top.MEM[55][5] ),
    .B2(_09810_),
    .X(_04157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17922_ (.A1(_00577_),
    .A2(_09809_),
    .B1(\design_top.MEM[55][4] ),
    .B2(_09810_),
    .X(_04156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17923_ (.A1(_00576_),
    .A2(_09809_),
    .B1(\design_top.MEM[55][3] ),
    .B2(_09810_),
    .X(_04155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17924_ (.A1(_00575_),
    .A2(_09808_),
    .B1(\design_top.MEM[55][2] ),
    .B2(_09807_),
    .X(_04154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17925_ (.A1(_00574_),
    .A2(_09808_),
    .B1(\design_top.MEM[55][1] ),
    .B2(_09807_),
    .X(_04153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17926_ (.A1(_00573_),
    .A2(_09808_),
    .B1(\design_top.MEM[55][0] ),
    .B2(_09807_),
    .X(_04152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17927_ (.A(_08325_),
    .Y(_09811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _17928_ (.A(_10823_),
    .B(_09811_),
    .X(_09812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _17929_ (.A(_02660_),
    .B(\design_top.DADDR[2] ),
    .C(_10828_),
    .X(_09813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _17930_ (.A(_09812_),
    .B(_09813_),
    .X(_09814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17931_ (.A(_09814_),
    .X(_09815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17932_ (.A(_09814_),
    .Y(_09816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17933_ (.A(_09816_),
    .X(_09817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17934_ (.A1(\design_top.GPIOFF[15] ),
    .A2(_09815_),
    .B1(\design_top.DATAO[31] ),
    .B2(_09817_),
    .X(_04151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17935_ (.A1(\design_top.GPIOFF[14] ),
    .A2(_09815_),
    .B1(\design_top.DATAO[30] ),
    .B2(_09817_),
    .X(_04150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17936_ (.A1(\design_top.GPIOFF[13] ),
    .A2(_09815_),
    .B1(\design_top.DATAO[29] ),
    .B2(_09817_),
    .X(_04149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17937_ (.A1(\design_top.GPIOFF[12] ),
    .A2(_09815_),
    .B1(\design_top.DATAO[28] ),
    .B2(_09817_),
    .X(_04148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17938_ (.A1(\design_top.GPIOFF[11] ),
    .A2(_09815_),
    .B1(\design_top.DATAO[27] ),
    .B2(_09817_),
    .X(_04147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17939_ (.A(_09814_),
    .X(_09818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17940_ (.A(_09816_),
    .X(_09819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17941_ (.A1(\design_top.GPIOFF[10] ),
    .A2(_09818_),
    .B1(\design_top.DATAO[26] ),
    .B2(_09819_),
    .X(_04146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17942_ (.A1(\design_top.GPIOFF[9] ),
    .A2(_09818_),
    .B1(\design_top.DATAO[25] ),
    .B2(_09819_),
    .X(_04145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17943_ (.A1(\design_top.GPIOFF[8] ),
    .A2(_09818_),
    .B1(\design_top.DATAO[24] ),
    .B2(_09819_),
    .X(_04144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17944_ (.A1(\design_top.GPIOFF[7] ),
    .A2(_09818_),
    .B1(\design_top.DATAO[23] ),
    .B2(_09819_),
    .X(_04143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17945_ (.A1(\design_top.GPIOFF[6] ),
    .A2(_09818_),
    .B1(\design_top.DATAO[22] ),
    .B2(_09819_),
    .X(_04142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17946_ (.A(_09814_),
    .X(_09820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17947_ (.A(_09816_),
    .X(_09821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17948_ (.A1(\design_top.GPIOFF[5] ),
    .A2(_09820_),
    .B1(\design_top.DATAO[21] ),
    .B2(_09821_),
    .X(_04141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17949_ (.A1(\design_top.GPIOFF[4] ),
    .A2(_09820_),
    .B1(\design_top.DATAO[20] ),
    .B2(_09821_),
    .X(_04140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17950_ (.A1(\design_top.GPIOFF[3] ),
    .A2(_09820_),
    .B1(\design_top.DATAO[19] ),
    .B2(_09821_),
    .X(_04139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17951_ (.A1(\design_top.GPIOFF[2] ),
    .A2(_09820_),
    .B1(\design_top.DATAO[18] ),
    .B2(_09821_),
    .X(_04138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17952_ (.A1(\design_top.GPIOFF[1] ),
    .A2(_09820_),
    .B1(\design_top.DATAO[17] ),
    .B2(_09821_),
    .X(_04137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17953_ (.A1(io_out[15]),
    .A2(_09814_),
    .B1(\design_top.DATAO[16] ),
    .B2(_09816_),
    .X(_04136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _17954_ (.A(_03200_),
    .B(_09813_),
    .X(_09822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17955_ (.A(_09822_),
    .X(_09823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _17956_ (.A(_09822_),
    .Y(_09824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17957_ (.A(_09824_),
    .X(_09825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17958_ (.A1(\design_top.LEDFF[15] ),
    .A2(_09823_),
    .B1(\design_top.DATAO[15] ),
    .B2(_09825_),
    .X(_04135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17959_ (.A1(\design_top.LEDFF[14] ),
    .A2(_09823_),
    .B1(\design_top.DATAO[14] ),
    .B2(_09825_),
    .X(_04134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17960_ (.A1(\design_top.LEDFF[13] ),
    .A2(_09823_),
    .B1(\design_top.DATAO[13] ),
    .B2(_09825_),
    .X(_04133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17961_ (.A1(\design_top.LEDFF[12] ),
    .A2(_09823_),
    .B1(\design_top.DATAO[12] ),
    .B2(_09825_),
    .X(_04132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17962_ (.A1(\design_top.LEDFF[11] ),
    .A2(_09823_),
    .B1(\design_top.DATAO[11] ),
    .B2(_09825_),
    .X(_04131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17963_ (.A(_09822_),
    .X(_09826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17964_ (.A(_09824_),
    .X(_09827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17965_ (.A1(\design_top.LEDFF[10] ),
    .A2(_09826_),
    .B1(\design_top.DATAO[10] ),
    .B2(_09827_),
    .X(_04130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17966_ (.A1(\design_top.LEDFF[9] ),
    .A2(_09826_),
    .B1(\design_top.DATAO[9] ),
    .B2(_09827_),
    .X(_04129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17967_ (.A1(\design_top.LEDFF[8] ),
    .A2(_09826_),
    .B1(\design_top.DATAO[8] ),
    .B2(_09827_),
    .X(_04128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17968_ (.A1(\design_top.LEDFF[7] ),
    .A2(_09826_),
    .B1(\design_top.DATAO[7] ),
    .B2(_09827_),
    .X(_04127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17969_ (.A1(\design_top.LEDFF[6] ),
    .A2(_09826_),
    .B1(\design_top.DATAO[6] ),
    .B2(_09827_),
    .X(_04126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17970_ (.A(_09822_),
    .X(_09828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17971_ (.A(_09824_),
    .X(_09829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17972_ (.A1(\design_top.LEDFF[5] ),
    .A2(_09828_),
    .B1(\design_top.DATAO[5] ),
    .B2(_09829_),
    .X(_04125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17973_ (.A1(\design_top.LEDFF[4] ),
    .A2(_09828_),
    .B1(\design_top.DATAO[4] ),
    .B2(_09829_),
    .X(_04124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17974_ (.A1(io_out[11]),
    .A2(_09828_),
    .B1(\design_top.DATAO[3] ),
    .B2(_09829_),
    .X(_04123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17975_ (.A1(io_out[10]),
    .A2(_09828_),
    .B1(\design_top.DATAO[2] ),
    .B2(_09829_),
    .X(_04122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17976_ (.A1(io_out[9]),
    .A2(_09828_),
    .B1(\design_top.DATAO[1] ),
    .B2(_09829_),
    .X(_04121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17977_ (.A1(io_out[8]),
    .A2(_09822_),
    .B1(\design_top.DATAO[0] ),
    .B2(_09824_),
    .X(_04120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17978_ (.A1(\design_top.ROMFF2[31] ),
    .A2(_08526_),
    .B1(\design_top.ROMFF[31] ),
    .B2(\design_top.HLT ),
    .X(_04119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17979_ (.A1(\design_top.ROMFF2[30] ),
    .A2(_08526_),
    .B1(\design_top.ROMFF[30] ),
    .B2(\design_top.HLT ),
    .X(_04118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17980_ (.A1(\design_top.ROMFF2[29] ),
    .A2(_08526_),
    .B1(\design_top.ROMFF[29] ),
    .B2(\design_top.HLT ),
    .X(_04117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17981_ (.A(_08473_),
    .X(_09830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17982_ (.A1(\design_top.ROMFF2[28] ),
    .A2(_08526_),
    .B1(\design_top.ROMFF[28] ),
    .B2(_09830_),
    .X(_04116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17983_ (.A(_08478_),
    .X(_09831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17984_ (.A1(\design_top.ROMFF2[27] ),
    .A2(_09831_),
    .B1(\design_top.ROMFF[27] ),
    .B2(_09830_),
    .X(_04115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17985_ (.A1(\design_top.ROMFF2[26] ),
    .A2(_09831_),
    .B1(\design_top.ROMFF[26] ),
    .B2(_09830_),
    .X(_04114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17986_ (.A1(\design_top.ROMFF2[25] ),
    .A2(_09831_),
    .B1(\design_top.ROMFF[25] ),
    .B2(_09830_),
    .X(_04113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17987_ (.A1(\design_top.ROMFF2[24] ),
    .A2(_09831_),
    .B1(\design_top.ROMFF[24] ),
    .B2(_09830_),
    .X(_04112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17988_ (.A(_08370_),
    .X(_09832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17989_ (.A(_09832_),
    .X(_09833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17990_ (.A1(\design_top.ROMFF2[23] ),
    .A2(_09831_),
    .B1(\design_top.ROMFF[23] ),
    .B2(_09833_),
    .X(_04111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17991_ (.A(_08438_),
    .X(_09834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17992_ (.A(_09834_),
    .X(_09835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17993_ (.A1(\design_top.ROMFF2[22] ),
    .A2(_09835_),
    .B1(\design_top.ROMFF[22] ),
    .B2(_09833_),
    .X(_04110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17994_ (.A1(\design_top.ROMFF2[21] ),
    .A2(_09835_),
    .B1(\design_top.ROMFF[21] ),
    .B2(_09833_),
    .X(_04109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17995_ (.A1(\design_top.ROMFF2[20] ),
    .A2(_09835_),
    .B1(\design_top.ROMFF[20] ),
    .B2(_09833_),
    .X(_04108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17996_ (.A1(\design_top.ROMFF2[19] ),
    .A2(_09835_),
    .B1(\design_top.ROMFF[19] ),
    .B2(_09833_),
    .X(_04107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17997_ (.A(_09832_),
    .X(_09836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _17998_ (.A1(\design_top.ROMFF2[18] ),
    .A2(_09835_),
    .B1(\design_top.ROMFF[18] ),
    .B2(_09836_),
    .X(_04106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _17999_ (.A(_09834_),
    .X(_09837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18000_ (.A1(\design_top.ROMFF2[17] ),
    .A2(_09837_),
    .B1(\design_top.ROMFF[17] ),
    .B2(_09836_),
    .X(_04105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18001_ (.A1(\design_top.ROMFF2[16] ),
    .A2(_09837_),
    .B1(\design_top.ROMFF[16] ),
    .B2(_09836_),
    .X(_04104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18002_ (.A1(\design_top.ROMFF2[15] ),
    .A2(_09837_),
    .B1(\design_top.ROMFF[15] ),
    .B2(_09836_),
    .X(_04103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18003_ (.A1(\design_top.ROMFF2[14] ),
    .A2(_09837_),
    .B1(\design_top.ROMFF[14] ),
    .B2(_09836_),
    .X(_04102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18004_ (.A(_09832_),
    .X(_09838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18005_ (.A1(\design_top.ROMFF2[13] ),
    .A2(_09837_),
    .B1(\design_top.ROMFF[13] ),
    .B2(_09838_),
    .X(_04101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18006_ (.A(_09834_),
    .X(_09839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18007_ (.A1(\design_top.ROMFF2[12] ),
    .A2(_09839_),
    .B1(\design_top.ROMFF[12] ),
    .B2(_09838_),
    .X(_04100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18008_ (.A1(\design_top.ROMFF2[11] ),
    .A2(_09839_),
    .B1(\design_top.ROMFF[11] ),
    .B2(_09838_),
    .X(_04099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18009_ (.A1(\design_top.ROMFF2[10] ),
    .A2(_09839_),
    .B1(\design_top.ROMFF[10] ),
    .B2(_09838_),
    .X(_04098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18010_ (.A1(\design_top.ROMFF2[9] ),
    .A2(_09839_),
    .B1(\design_top.ROMFF[9] ),
    .B2(_09838_),
    .X(_04097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18011_ (.A(_09832_),
    .X(_09840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18012_ (.A1(\design_top.ROMFF2[8] ),
    .A2(_09839_),
    .B1(\design_top.ROMFF[8] ),
    .B2(_09840_),
    .X(_04096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18013_ (.A(_09834_),
    .X(_09841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18014_ (.A1(\design_top.ROMFF2[7] ),
    .A2(_09841_),
    .B1(\design_top.ROMFF[7] ),
    .B2(_09840_),
    .X(_04095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18015_ (.A1(\design_top.ROMFF2[6] ),
    .A2(_09841_),
    .B1(\design_top.ROMFF[6] ),
    .B2(_09840_),
    .X(_04094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18016_ (.A1(\design_top.ROMFF2[5] ),
    .A2(_09841_),
    .B1(\design_top.ROMFF[5] ),
    .B2(_09840_),
    .X(_04093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18017_ (.A1(\design_top.ROMFF2[4] ),
    .A2(_09841_),
    .B1(\design_top.ROMFF[4] ),
    .B2(_09840_),
    .X(_04092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18018_ (.A(_09832_),
    .X(_09842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18019_ (.A1(\design_top.ROMFF2[3] ),
    .A2(_09841_),
    .B1(\design_top.ROMFF[3] ),
    .B2(_09842_),
    .X(_04091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18020_ (.A(_09834_),
    .X(_09843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18021_ (.A1(\design_top.ROMFF2[2] ),
    .A2(_09843_),
    .B1(\design_top.ROMFF[2] ),
    .B2(_09842_),
    .X(_04090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18022_ (.A1(\design_top.ROMFF2[1] ),
    .A2(_09843_),
    .B1(\design_top.ROMFF[1] ),
    .B2(_09842_),
    .X(_04089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18023_ (.A1(\design_top.ROMFF2[0] ),
    .A2(_09843_),
    .B1(\design_top.ROMFF[0] ),
    .B2(_09842_),
    .X(_04088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18024_ (.A1(\design_top.uart0.UART_XREQ ),
    .A2(_08619_),
    .B1(\design_top.uart0.UART_XACK ),
    .B2(_08620_),
    .X(_04087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18025_ (.A(\design_top.uart0.UART_RACK ),
    .Y(_09844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _18026_ (.A0(_09844_),
    .A1(\design_top.uart0.UART_RREQ ),
    .S(_08631_),
    .X(_04086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18027_ (.A(\design_top.uart0.UART_RXDFF[2] ),
    .X(_09845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _18028_ (.A(_08638_),
    .B(_08639_),
    .C(_08629_),
    .D(_08624_),
    .X(_09846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _18029_ (.A0(_09845_),
    .A1(\design_top.uart0.UART_RFIFO[7] ),
    .S(_09846_),
    .X(_04085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _18030_ (.A(_08641_),
    .B(_08639_),
    .C(_08629_),
    .D(_08623_),
    .X(_09847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _18031_ (.A0(_09845_),
    .A1(\design_top.uart0.UART_RFIFO[6] ),
    .S(_09847_),
    .X(_04084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18032_ (.A(_08628_),
    .X(_09848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _18033_ (.A(_08638_),
    .B(_08630_),
    .C(_09848_),
    .D(_08623_),
    .X(_09849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _18034_ (.A0(_09845_),
    .A1(\design_top.uart0.UART_RFIFO[5] ),
    .S(_09849_),
    .X(_04083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _18035_ (.A(_08629_),
    .B(_08624_),
    .C(_08641_),
    .D(_08630_),
    .X(_09850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _18036_ (.A0(_09845_),
    .A1(\design_top.uart0.UART_RFIFO[4] ),
    .S(_09850_),
    .X(_04082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _18037_ (.A(_08638_),
    .B(_08639_),
    .C(_09848_),
    .D(_08635_),
    .X(_09851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _18038_ (.A0(\design_top.uart0.UART_RXDFF[2] ),
    .A1(\design_top.uart0.UART_RFIFO[3] ),
    .S(_09851_),
    .X(_04081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _18039_ (.A(_08641_),
    .B(_08639_),
    .C(_09848_),
    .D(_08635_),
    .X(_09852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _18040_ (.A0(\design_top.uart0.UART_RXDFF[2] ),
    .A1(\design_top.uart0.UART_RFIFO[2] ),
    .S(_09852_),
    .X(_04080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _18041_ (.A(_08625_),
    .B(_08630_),
    .C(_09848_),
    .D(_08635_),
    .X(_09853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _18042_ (.A0(\design_top.uart0.UART_RXDFF[2] ),
    .A1(\design_top.uart0.UART_RFIFO[1] ),
    .S(_09853_),
    .X(_04079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _18043_ (.A(_08641_),
    .B(_08630_),
    .C(_09848_),
    .D(_08635_),
    .X(_09854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _18044_ (.A0(\design_top.uart0.UART_RXDFF[2] ),
    .A1(\design_top.uart0.UART_RFIFO[0] ),
    .S(_09854_),
    .X(_04078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18045_ (.A1(\design_top.core0.NXPC[31] ),
    .A2(_09843_),
    .B1(\design_top.core0.PC[31] ),
    .B2(_09842_),
    .X(_04077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18046_ (.A(_08370_),
    .X(_09855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18047_ (.A(_09855_),
    .X(_09856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18048_ (.A1(\design_top.core0.NXPC[30] ),
    .A2(_09843_),
    .B1(\design_top.core0.PC[30] ),
    .B2(_09856_),
    .X(_04076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18049_ (.A(_08438_),
    .X(_09857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18050_ (.A(_09857_),
    .X(_09858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18051_ (.A1(\design_top.core0.NXPC[29] ),
    .A2(_09858_),
    .B1(\design_top.core0.PC[29] ),
    .B2(_09856_),
    .X(_04075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18052_ (.A1(\design_top.core0.NXPC[28] ),
    .A2(_09858_),
    .B1(\design_top.core0.PC[28] ),
    .B2(_09856_),
    .X(_04074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18053_ (.A1(\design_top.core0.NXPC[27] ),
    .A2(_09858_),
    .B1(\design_top.core0.PC[27] ),
    .B2(_09856_),
    .X(_04073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18054_ (.A1(\design_top.core0.NXPC[26] ),
    .A2(_09858_),
    .B1(\design_top.core0.PC[26] ),
    .B2(_09856_),
    .X(_04072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18055_ (.A(_09855_),
    .X(_09859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18056_ (.A1(\design_top.core0.NXPC[25] ),
    .A2(_09858_),
    .B1(\design_top.core0.PC[25] ),
    .B2(_09859_),
    .X(_04071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18057_ (.A(_09857_),
    .X(_09860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18058_ (.A1(\design_top.core0.NXPC[24] ),
    .A2(_09860_),
    .B1(\design_top.core0.PC[24] ),
    .B2(_09859_),
    .X(_04070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18059_ (.A1(\design_top.core0.NXPC[23] ),
    .A2(_09860_),
    .B1(\design_top.core0.PC[23] ),
    .B2(_09859_),
    .X(_04069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18060_ (.A1(\design_top.core0.NXPC[22] ),
    .A2(_09860_),
    .B1(\design_top.core0.PC[22] ),
    .B2(_09859_),
    .X(_04068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18061_ (.A1(\design_top.core0.NXPC[21] ),
    .A2(_09860_),
    .B1(\design_top.core0.PC[21] ),
    .B2(_09859_),
    .X(_04067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18062_ (.A(_09855_),
    .X(_09861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18063_ (.A1(\design_top.core0.NXPC[20] ),
    .A2(_09860_),
    .B1(\design_top.core0.PC[20] ),
    .B2(_09861_),
    .X(_04066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18064_ (.A(_09857_),
    .X(_09862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18065_ (.A1(\design_top.core0.NXPC[19] ),
    .A2(_09862_),
    .B1(\design_top.core0.PC[19] ),
    .B2(_09861_),
    .X(_04065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18066_ (.A1(\design_top.core0.NXPC[18] ),
    .A2(_09862_),
    .B1(\design_top.core0.PC[18] ),
    .B2(_09861_),
    .X(_04064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18067_ (.A1(\design_top.core0.NXPC[17] ),
    .A2(_09862_),
    .B1(\design_top.core0.PC[17] ),
    .B2(_09861_),
    .X(_04063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18068_ (.A1(\design_top.core0.NXPC[16] ),
    .A2(_09862_),
    .B1(\design_top.core0.PC[16] ),
    .B2(_09861_),
    .X(_04062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18069_ (.A(_09855_),
    .X(_09863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18070_ (.A1(\design_top.core0.NXPC[15] ),
    .A2(_09862_),
    .B1(\design_top.core0.PC[15] ),
    .B2(_09863_),
    .X(_04061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18071_ (.A(_09857_),
    .X(_09864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18072_ (.A1(\design_top.core0.NXPC[14] ),
    .A2(_09864_),
    .B1(\design_top.core0.PC[14] ),
    .B2(_09863_),
    .X(_04060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18073_ (.A1(\design_top.core0.NXPC[13] ),
    .A2(_09864_),
    .B1(\design_top.core0.PC[13] ),
    .B2(_09863_),
    .X(_04059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18074_ (.A1(\design_top.core0.NXPC[12] ),
    .A2(_09864_),
    .B1(\design_top.core0.PC[12] ),
    .B2(_09863_),
    .X(_04058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18075_ (.A1(\design_top.core0.NXPC[11] ),
    .A2(_09864_),
    .B1(\design_top.core0.PC[11] ),
    .B2(_09863_),
    .X(_04057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18076_ (.A(_09855_),
    .X(_09865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18077_ (.A1(\design_top.core0.NXPC[10] ),
    .A2(_09864_),
    .B1(\design_top.core0.PC[10] ),
    .B2(_09865_),
    .X(_04056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18078_ (.A(_09857_),
    .X(_09866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18079_ (.A1(\design_top.core0.NXPC[9] ),
    .A2(_09866_),
    .B1(\design_top.core0.PC[9] ),
    .B2(_09865_),
    .X(_04055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18080_ (.A1(\design_top.core0.NXPC[8] ),
    .A2(_09866_),
    .B1(\design_top.core0.PC[8] ),
    .B2(_09865_),
    .X(_04054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18081_ (.A1(\design_top.core0.NXPC[7] ),
    .A2(_09866_),
    .B1(\design_top.core0.PC[7] ),
    .B2(_09865_),
    .X(_04053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18082_ (.A1(\design_top.core0.NXPC[6] ),
    .A2(_09866_),
    .B1(\design_top.core0.PC[6] ),
    .B2(_09865_),
    .X(_04052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18083_ (.A(_08370_),
    .X(_09867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18084_ (.A(_09867_),
    .X(_09868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18085_ (.A1(\design_top.core0.NXPC[5] ),
    .A2(_09866_),
    .B1(\design_top.core0.PC[5] ),
    .B2(_09868_),
    .X(_04051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18086_ (.A(_08438_),
    .X(_09869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18087_ (.A(_09869_),
    .X(_09870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18088_ (.A1(\design_top.core0.NXPC[4] ),
    .A2(_09870_),
    .B1(\design_top.core0.PC[4] ),
    .B2(_09868_),
    .X(_04050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18089_ (.A1(\design_top.core0.NXPC[3] ),
    .A2(_09870_),
    .B1(\design_top.core0.PC[3] ),
    .B2(_09868_),
    .X(_04049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18090_ (.A1(\design_top.core0.NXPC[2] ),
    .A2(_09870_),
    .B1(\design_top.core0.PC[2] ),
    .B2(_09868_),
    .X(_04048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18091_ (.A1(\design_top.core0.NXPC[1] ),
    .A2(_09870_),
    .B1(\design_top.core0.PC[1] ),
    .B2(_09868_),
    .X(_04047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18092_ (.A(_09867_),
    .X(_09871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18093_ (.A1(\design_top.core0.NXPC[0] ),
    .A2(_09870_),
    .B1(\design_top.core0.PC[0] ),
    .B2(_09871_),
    .X(_04046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18094_ (.A(_09869_),
    .X(_09872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18095_ (.A1(\design_top.IADDR[31] ),
    .A2(_09872_),
    .B1(\design_top.core0.NXPC[31] ),
    .B2(_09871_),
    .X(_04045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18096_ (.A1(\design_top.IADDR[30] ),
    .A2(_09872_),
    .B1(\design_top.core0.NXPC[30] ),
    .B2(_09871_),
    .X(_04044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18097_ (.A1(\design_top.IADDR[29] ),
    .A2(_09872_),
    .B1(\design_top.core0.NXPC[29] ),
    .B2(_09871_),
    .X(_04043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18098_ (.A1(\design_top.IADDR[28] ),
    .A2(_09872_),
    .B1(\design_top.core0.NXPC[28] ),
    .B2(_09871_),
    .X(_04042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18099_ (.A(_09867_),
    .X(_09873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18100_ (.A1(\design_top.IADDR[27] ),
    .A2(_09872_),
    .B1(\design_top.core0.NXPC[27] ),
    .B2(_09873_),
    .X(_04041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18101_ (.A(_09869_),
    .X(_09874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18102_ (.A1(\design_top.IADDR[26] ),
    .A2(_09874_),
    .B1(\design_top.core0.NXPC[26] ),
    .B2(_09873_),
    .X(_04040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18103_ (.A1(\design_top.IADDR[25] ),
    .A2(_09874_),
    .B1(\design_top.core0.NXPC[25] ),
    .B2(_09873_),
    .X(_04039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18104_ (.A1(\design_top.IADDR[24] ),
    .A2(_09874_),
    .B1(\design_top.core0.NXPC[24] ),
    .B2(_09873_),
    .X(_04038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18105_ (.A1(\design_top.IADDR[23] ),
    .A2(_09874_),
    .B1(\design_top.core0.NXPC[23] ),
    .B2(_09873_),
    .X(_04037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18106_ (.A(_09867_),
    .X(_09875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18107_ (.A1(\design_top.IADDR[22] ),
    .A2(_09874_),
    .B1(\design_top.core0.NXPC[22] ),
    .B2(_09875_),
    .X(_04036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18108_ (.A(_09869_),
    .X(_09876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18109_ (.A1(\design_top.IADDR[21] ),
    .A2(_09876_),
    .B1(\design_top.core0.NXPC[21] ),
    .B2(_09875_),
    .X(_04035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18110_ (.A1(\design_top.IADDR[20] ),
    .A2(_09876_),
    .B1(\design_top.core0.NXPC[20] ),
    .B2(_09875_),
    .X(_04034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18111_ (.A1(\design_top.IADDR[19] ),
    .A2(_09876_),
    .B1(\design_top.core0.NXPC[19] ),
    .B2(_09875_),
    .X(_04033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18112_ (.A1(\design_top.IADDR[18] ),
    .A2(_09876_),
    .B1(\design_top.core0.NXPC[18] ),
    .B2(_09875_),
    .X(_04032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18113_ (.A(_09867_),
    .X(_09877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18114_ (.A1(\design_top.IADDR[17] ),
    .A2(_09876_),
    .B1(\design_top.core0.NXPC[17] ),
    .B2(_09877_),
    .X(_04031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18115_ (.A(_09869_),
    .X(_09878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18116_ (.A1(\design_top.IADDR[16] ),
    .A2(_09878_),
    .B1(\design_top.core0.NXPC[16] ),
    .B2(_09877_),
    .X(_04030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18117_ (.A1(\design_top.IADDR[15] ),
    .A2(_09878_),
    .B1(\design_top.core0.NXPC[15] ),
    .B2(_09877_),
    .X(_04029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18118_ (.A1(\design_top.IADDR[14] ),
    .A2(_09878_),
    .B1(\design_top.core0.NXPC[14] ),
    .B2(_09877_),
    .X(_04028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18119_ (.A1(\design_top.IADDR[13] ),
    .A2(_09878_),
    .B1(\design_top.core0.NXPC[13] ),
    .B2(_09877_),
    .X(_04027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18120_ (.A(_08353_),
    .X(_09879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18121_ (.A1(\design_top.IADDR[12] ),
    .A2(_09878_),
    .B1(\design_top.core0.NXPC[12] ),
    .B2(_09879_),
    .X(_04026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18122_ (.A(_08439_),
    .X(_09880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18123_ (.A1(\design_top.IADDR[11] ),
    .A2(_09880_),
    .B1(\design_top.core0.NXPC[11] ),
    .B2(_09879_),
    .X(_04025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18124_ (.A1(\design_top.IADDR[10] ),
    .A2(_09880_),
    .B1(\design_top.core0.NXPC[10] ),
    .B2(_09879_),
    .X(_04024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18125_ (.A1(\design_top.IADDR[9] ),
    .A2(_09880_),
    .B1(\design_top.core0.NXPC[9] ),
    .B2(_09879_),
    .X(_04023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18126_ (.A1(\design_top.IADDR[8] ),
    .A2(_09880_),
    .B1(\design_top.core0.NXPC[8] ),
    .B2(_09879_),
    .X(_04022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18127_ (.A(_08353_),
    .X(_09881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18128_ (.A1(\design_top.IADDR[7] ),
    .A2(_09880_),
    .B1(\design_top.core0.NXPC[7] ),
    .B2(_09881_),
    .X(_04021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18129_ (.A(_08439_),
    .X(_09882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18130_ (.A1(\design_top.IADDR[6] ),
    .A2(_09882_),
    .B1(\design_top.core0.NXPC[6] ),
    .B2(_09881_),
    .X(_04020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18131_ (.A1(\design_top.IADDR[5] ),
    .A2(_09882_),
    .B1(\design_top.core0.NXPC[5] ),
    .B2(_09881_),
    .X(_04019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18132_ (.A1(_08525_),
    .A2(_09882_),
    .B1(\design_top.core0.NXPC[4] ),
    .B2(_09881_),
    .X(_04018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18133_ (.A1(io_out[19]),
    .A2(_09882_),
    .B1(\design_top.core0.NXPC[3] ),
    .B2(_09881_),
    .X(_04017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18134_ (.A1(io_out[18]),
    .A2(_09882_),
    .B1(\design_top.core0.NXPC[2] ),
    .B2(_08489_),
    .X(_04016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18135_ (.A1(io_out[17]),
    .A2(_08431_),
    .B1(\design_top.core0.NXPC[1] ),
    .B2(_08489_),
    .X(_04015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18136_ (.A1(io_out[16]),
    .A2(_08431_),
    .B1(\design_top.core0.NXPC[0] ),
    .B2(_08489_),
    .X(_04014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18137_ (.A(_08783_),
    .X(_09883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18138_ (.A(_09883_),
    .X(_09884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18139_ (.A(_09884_),
    .X(_09885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18140_ (.A(_09883_),
    .Y(_09886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18141_ (.A(_09886_),
    .X(_09887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18142_ (.A(_09887_),
    .X(_09888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18143_ (.A1(_09885_),
    .A2(_08800_),
    .B1(\design_top.core0.REG2[9][31] ),
    .B2(_09888_),
    .X(_04013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18144_ (.A1(_09885_),
    .A2(_08802_),
    .B1(\design_top.core0.REG2[9][30] ),
    .B2(_09888_),
    .X(_04012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18145_ (.A1(_09885_),
    .A2(_08804_),
    .B1(\design_top.core0.REG2[9][29] ),
    .B2(_09888_),
    .X(_04011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18146_ (.A1(_09885_),
    .A2(_08806_),
    .B1(\design_top.core0.REG2[9][28] ),
    .B2(_09888_),
    .X(_04010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18147_ (.A1(_09885_),
    .A2(_08809_),
    .B1(\design_top.core0.REG2[9][27] ),
    .B2(_09888_),
    .X(_04009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18148_ (.A(_09884_),
    .X(_09889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18149_ (.A(_09887_),
    .X(_09890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18150_ (.A1(_09889_),
    .A2(_08813_),
    .B1(\design_top.core0.REG2[9][26] ),
    .B2(_09890_),
    .X(_04008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18151_ (.A1(_09889_),
    .A2(_08815_),
    .B1(\design_top.core0.REG2[9][25] ),
    .B2(_09890_),
    .X(_04007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18152_ (.A1(_09889_),
    .A2(_08817_),
    .B1(\design_top.core0.REG2[9][24] ),
    .B2(_09890_),
    .X(_04006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18153_ (.A1(_09889_),
    .A2(_08819_),
    .B1(\design_top.core0.REG2[9][23] ),
    .B2(_09890_),
    .X(_04005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18154_ (.A1(_09889_),
    .A2(_08822_),
    .B1(\design_top.core0.REG2[9][22] ),
    .B2(_09890_),
    .X(_04004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18155_ (.A(_09884_),
    .X(_09891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18156_ (.A(_09887_),
    .X(_09892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18157_ (.A1(_09891_),
    .A2(_08826_),
    .B1(\design_top.core0.REG2[9][21] ),
    .B2(_09892_),
    .X(_04003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18158_ (.A1(_09891_),
    .A2(_08828_),
    .B1(\design_top.core0.REG2[9][20] ),
    .B2(_09892_),
    .X(_04002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18159_ (.A1(_09891_),
    .A2(_08830_),
    .B1(\design_top.core0.REG2[9][19] ),
    .B2(_09892_),
    .X(_04001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18160_ (.A1(_09891_),
    .A2(_08832_),
    .B1(\design_top.core0.REG2[9][18] ),
    .B2(_09892_),
    .X(_04000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18161_ (.A1(_09891_),
    .A2(_08835_),
    .B1(\design_top.core0.REG2[9][17] ),
    .B2(_09892_),
    .X(_03999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18162_ (.A(_09883_),
    .X(_09893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18163_ (.A(_09886_),
    .X(_09894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18164_ (.A1(_09893_),
    .A2(_08839_),
    .B1(\design_top.core0.REG2[9][16] ),
    .B2(_09894_),
    .X(_03998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18165_ (.A1(_09893_),
    .A2(_08841_),
    .B1(\design_top.core0.REG2[9][15] ),
    .B2(_09894_),
    .X(_03997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18166_ (.A1(_09893_),
    .A2(_08843_),
    .B1(\design_top.core0.REG2[9][14] ),
    .B2(_09894_),
    .X(_03996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18167_ (.A1(\design_top.core0.REG2[9][13] ),
    .A2(_09884_),
    .B1(_08844_),
    .B2(_09887_),
    .X(_03995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18168_ (.A1(_09893_),
    .A2(_08846_),
    .B1(\design_top.core0.REG2[9][12] ),
    .B2(_09894_),
    .X(_03994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18169_ (.A1(_09893_),
    .A2(_08849_),
    .B1(\design_top.core0.REG2[9][11] ),
    .B2(_09894_),
    .X(_03993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18170_ (.A(_09883_),
    .X(_09895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18171_ (.A(_09886_),
    .X(_09896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18172_ (.A1(_09895_),
    .A2(_08853_),
    .B1(\design_top.core0.REG2[9][10] ),
    .B2(_09896_),
    .X(_03992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18173_ (.A1(_09895_),
    .A2(_08855_),
    .B1(\design_top.core0.REG2[9][9] ),
    .B2(_09896_),
    .X(_03991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18174_ (.A1(_09895_),
    .A2(_08857_),
    .B1(\design_top.core0.REG2[9][8] ),
    .B2(_09896_),
    .X(_03990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18175_ (.A1(_09895_),
    .A2(_08859_),
    .B1(\design_top.core0.REG2[9][7] ),
    .B2(_09896_),
    .X(_03989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18176_ (.A1(_09895_),
    .A2(_08862_),
    .B1(\design_top.core0.REG2[9][6] ),
    .B2(_09896_),
    .X(_03988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18177_ (.A(_09883_),
    .X(_09897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18178_ (.A(_09886_),
    .X(_09898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18179_ (.A1(_09897_),
    .A2(_08866_),
    .B1(\design_top.core0.REG2[9][5] ),
    .B2(_09898_),
    .X(_03987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18180_ (.A1(_09897_),
    .A2(_08868_),
    .B1(\design_top.core0.REG2[9][4] ),
    .B2(_09898_),
    .X(_03986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18181_ (.A1(_09897_),
    .A2(_08870_),
    .B1(\design_top.core0.REG2[9][3] ),
    .B2(_09898_),
    .X(_03985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18182_ (.A1(_09897_),
    .A2(_08872_),
    .B1(\design_top.core0.REG2[9][2] ),
    .B2(_09898_),
    .X(_03984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18183_ (.A1(_09897_),
    .A2(_08874_),
    .B1(\design_top.core0.REG2[9][1] ),
    .B2(_09898_),
    .X(_03983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18184_ (.A1(_09884_),
    .A2(_08876_),
    .B1(\design_top.core0.REG2[9][0] ),
    .B2(_09887_),
    .X(_03982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3b_2 _18185_ (.A_N(\design_top.DACK[1] ),
    .B(\design_top.DACK[0] ),
    .C(io_out[12]),
    .X(_09899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _18186_ (.A(_02857_),
    .B(\design_top.DADDR[3] ),
    .C(_10827_),
    .X(_09900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18187_ (.A(_09900_),
    .Y(_09901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _18188_ (.A1(\design_top.DADDR[2] ),
    .A2(_09899_),
    .A3(_09901_),
    .B1(_08347_),
    .X(_09902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _18189_ (.A0(\design_top.uart0.UART_RACK ),
    .A1(\design_top.uart0.UART_RREQ ),
    .S(_09902_),
    .X(_03981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _18190_ (.A(_08369_),
    .B(_10596_),
    .C(_02651_),
    .D(_09900_),
    .X(_09903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18191_ (.A(_09903_),
    .X(_09904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2ai_2 _18192_ (.A1_N(\design_top.uart0.UART_XREQ ),
    .A2_N(_09904_),
    .B1(\design_top.uart0.UART_XACK ),
    .B2(_09904_),
    .Y(_03980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _18193_ (.A0(\design_top.DATAO[15] ),
    .A1(\design_top.uart0.UART_XFIFO[7] ),
    .S(_09904_),
    .X(_03979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _18194_ (.A0(\design_top.DATAO[14] ),
    .A1(\design_top.uart0.UART_XFIFO[6] ),
    .S(_09904_),
    .X(_03978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _18195_ (.A0(\design_top.DATAO[13] ),
    .A1(\design_top.uart0.UART_XFIFO[5] ),
    .S(_09904_),
    .X(_03977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18196_ (.A(_09903_),
    .X(_09905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _18197_ (.A0(\design_top.DATAO[12] ),
    .A1(\design_top.uart0.UART_XFIFO[4] ),
    .S(_09905_),
    .X(_03976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _18198_ (.A0(\design_top.DATAO[11] ),
    .A1(\design_top.uart0.UART_XFIFO[3] ),
    .S(_09905_),
    .X(_03975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _18199_ (.A0(\design_top.DATAO[10] ),
    .A1(\design_top.uart0.UART_XFIFO[2] ),
    .S(_09905_),
    .X(_03974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _18200_ (.A0(\design_top.DATAO[9] ),
    .A1(\design_top.uart0.UART_XFIFO[1] ),
    .S(_09905_),
    .X(_03973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _18201_ (.A0(\design_top.DATAO[8] ),
    .A1(\design_top.uart0.UART_XFIFO[0] ),
    .S(_09905_),
    .X(_03972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18202_ (.A(_10824_),
    .X(_09906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18203_ (.A(_09906_),
    .X(_02855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18204_ (.A(_09811_),
    .X(_09907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18205_ (.A(_09907_),
    .X(_02850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18206_ (.A(_09812_),
    .X(_09908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18207_ (.A(_09908_),
    .Y(_03273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18208_ (.A(_08751_),
    .X(_09909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18209_ (.A(_09909_),
    .X(_09910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18210_ (.A(_10959_),
    .B(_09910_),
    .Y(_03265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18211_ (.A(_10886_),
    .B(_09910_),
    .Y(_03266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18212_ (.A(_10825_),
    .X(_09911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18213_ (.A(_09911_),
    .Y(_02866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18214_ (.A(_03077_),
    .Y(_09912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18215_ (.A(_10825_),
    .X(_02867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18216_ (.A(_09912_),
    .B(_02867_),
    .Y(_03267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18217_ (.A(\design_top.core0.FCT3[2] ),
    .X(_09913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18218_ (.A(\design_top.core0.FCT3[0] ),
    .Y(_09914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18219_ (.A(_08502_),
    .B(_09914_),
    .X(_09915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18220_ (.A(_09915_),
    .X(_02849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18221_ (.A(_09913_),
    .B(_02849_),
    .Y(_02847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18222_ (.A(_03012_),
    .Y(_09916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18223_ (.A(_09916_),
    .B(_02850_),
    .Y(_03268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18224_ (.A(_10596_),
    .Y(io_out[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18225_ (.A(_08751_),
    .X(_09917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18226_ (.A(_09917_),
    .X(_09918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18227_ (.A(_11041_),
    .B(_09918_),
    .Y(_03261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18228_ (.A(_11020_),
    .B(_09910_),
    .Y(_03262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18229_ (.A(_11001_),
    .B(_09910_),
    .Y(_03263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18230_ (.A(_10981_),
    .B(_09910_),
    .Y(_03264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18231_ (.A(_11165_),
    .B(_09918_),
    .Y(_03257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18232_ (.A(_11150_),
    .B(_09918_),
    .Y(_03258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18233_ (.A(_11131_),
    .B(_09918_),
    .Y(_03259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18234_ (.A(_10784_),
    .B(_09918_),
    .Y(_03260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18235_ (.A(_09917_),
    .X(_09919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18236_ (.A(_11257_),
    .B(_09919_),
    .Y(_03253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18237_ (.A(_11240_),
    .B(_09919_),
    .Y(_03254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18238_ (.A(_11226_),
    .B(_09919_),
    .Y(_03255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18239_ (.A(_11192_),
    .B(_09919_),
    .Y(_03256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18240_ (.A(_09917_),
    .X(_09920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18241_ (.A(_11355_),
    .B(_09920_),
    .Y(_03248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18242_ (.A(_11342_),
    .B(_09920_),
    .Y(_03249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18243_ (.A(_11277_),
    .B(_09919_),
    .Y(_03250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18244_ (.A(_11287_),
    .B(_09920_),
    .Y(_03251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18245_ (.A(_11106_),
    .B(_09920_),
    .Y(_03252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18246_ (.A(_09917_),
    .X(_09921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18247_ (.A(_07505_),
    .B(_09921_),
    .Y(_03243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18248_ (.A(_07472_),
    .B(_09921_),
    .Y(_03244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18249_ (.A(_07956_),
    .B(_09921_),
    .Y(_03245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18250_ (.A(_07442_),
    .B(_09921_),
    .Y(_03246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18251_ (.A(_11327_),
    .B(_09920_),
    .Y(_03247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18252_ (.A(_09917_),
    .X(_09922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18253_ (.A(_07602_),
    .B(_09922_),
    .Y(_03237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18254_ (.A(_07567_),
    .B(_09922_),
    .Y(_03238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18255_ (.A(_07577_),
    .B(_09922_),
    .Y(_03239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18256_ (.A(_07643_),
    .B(_09921_),
    .Y(_03240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18257_ (.A(_07528_),
    .B(_09922_),
    .Y(_03241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18258_ (.A(_07516_),
    .B(_09922_),
    .Y(_03242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18259_ (.A(_08751_),
    .X(_09923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18260_ (.A(_09923_),
    .X(_09924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18261_ (.A(_07703_),
    .B(_09924_),
    .Y(_03235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18262_ (.A(_07698_),
    .B(_09924_),
    .Y(_03236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18263_ (.A(_09923_),
    .X(_09925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18264_ (.A(_07781_),
    .B(_09925_),
    .Y(_03231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18265_ (.A(_07772_),
    .B(_09924_),
    .Y(_03232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18266_ (.A(_07751_),
    .B(_09924_),
    .Y(_03233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18267_ (.A(_07728_),
    .B(_09924_),
    .Y(_03234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18268_ (.A(_09923_),
    .X(_09926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18269_ (.A(_07906_),
    .B(_09926_),
    .Y(_03226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18270_ (.A(_07864_),
    .B(_09925_),
    .Y(_03227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18271_ (.A(_07851_),
    .B(_09925_),
    .Y(_03228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18272_ (.A(_07828_),
    .B(_09925_),
    .Y(_03229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18273_ (.A(_07822_),
    .B(_09925_),
    .Y(_03230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18274_ (.A(_07451_),
    .B(_09926_),
    .Y(_03223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18275_ (.A(_07930_),
    .B(_09926_),
    .Y(_03224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18276_ (.A(_07559_),
    .B(_09926_),
    .Y(_03225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18277_ (.A(_09923_),
    .X(_09927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18278_ (.A(_07671_),
    .B(_09927_),
    .Y(_03219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18279_ (.A(_08019_),
    .B(_09927_),
    .Y(_03220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18280_ (.A(_07978_),
    .B(_09927_),
    .Y(_03221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18281_ (.A(_07973_),
    .B(_09926_),
    .Y(_03222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18282_ (.A(_08068_),
    .B(_09927_),
    .Y(_03217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18283_ (.A(_08044_),
    .B(_09927_),
    .Y(_03218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18284_ (.A(_09923_),
    .X(_09928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18285_ (.A(_08166_),
    .B(_09928_),
    .Y(_03211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18286_ (.A(_08150_),
    .B(_09928_),
    .Y(_03212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18287_ (.A(_08134_),
    .B(_09928_),
    .Y(_03213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18288_ (.A(_08120_),
    .B(_09928_),
    .Y(_03214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18289_ (.A(_08103_),
    .B(_09928_),
    .Y(_03215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18290_ (.A(_08751_),
    .X(_09929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18291_ (.A(_08238_),
    .B(_09929_),
    .Y(_03208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18292_ (.A(_08224_),
    .B(_09929_),
    .Y(_03209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18293_ (.A(_08193_),
    .B(_09929_),
    .Y(_03210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18294_ (.A(_08295_),
    .B(_09909_),
    .Y(_03204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18295_ (.A(_08281_),
    .B(_09909_),
    .Y(_03205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18296_ (.A(_08265_),
    .B(_09929_),
    .Y(_03206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18297_ (.A(_08252_),
    .B(_09929_),
    .Y(_03207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18298_ (.A(_07624_),
    .B(_09909_),
    .Y(_03202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18299_ (.A(_08308_),
    .B(_09909_),
    .Y(_03203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18300_ (.A1_N(\design_top.IACK[7] ),
    .A2_N(\design_top.IREQ[7] ),
    .B1(\design_top.IACK[7] ),
    .B2(\design_top.IREQ[7] ),
    .X(_03198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18301_ (.A(\design_top.IDATA[20] ),
    .Y(_09930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18302_ (.A(_08362_),
    .X(_09931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor4_2 _18303_ (.A(_09930_),
    .B(_00009_),
    .C(_00008_),
    .D(_09931_),
    .Y(_00700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18304_ (.A(_08362_),
    .X(_09932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18305_ (.A(_08402_),
    .B(_09932_),
    .Y(_00701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18306_ (.A(_08397_),
    .B(_09932_),
    .Y(_00704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18307_ (.A(_08394_),
    .B(_09932_),
    .Y(_00707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18308_ (.A(_08392_),
    .B(_09932_),
    .Y(_00711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18309_ (.A(_08390_),
    .B(_09932_),
    .Y(_00714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18310_ (.A(_08362_),
    .X(_09933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18311_ (.A(_08388_),
    .B(_09933_),
    .Y(_00717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18312_ (.A(_08383_),
    .B(_09933_),
    .Y(_00720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18313_ (.A(_08381_),
    .B(_09933_),
    .Y(_00723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18314_ (.A(_08377_),
    .B(_09933_),
    .Y(_00726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18315_ (.A(_08372_),
    .B(_09933_),
    .Y(_00729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18316_ (.A(_08362_),
    .X(_09934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18317_ (.A(_08351_),
    .B(_09934_),
    .Y(_00732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _18318_ (.A(\design_top.IDATA[12] ),
    .B(_09934_),
    .X(_00735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _18319_ (.A(\design_top.IDATA[13] ),
    .B(_09934_),
    .X(_00738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _18320_ (.A(\design_top.IDATA[14] ),
    .B(_09934_),
    .X(_00740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _18321_ (.A(\design_top.IDATA[15] ),
    .B(_09934_),
    .X(_00742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _18322_ (.A(\design_top.IDATA[16] ),
    .B(_09931_),
    .X(_00744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _18323_ (.A(\design_top.IDATA[17] ),
    .B(_09931_),
    .X(_00746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _18324_ (.A(\design_top.IDATA[18] ),
    .B(_09931_),
    .X(_00748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _18325_ (.A(_03936_),
    .B(_09931_),
    .X(_00750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18326_ (.A(_09930_),
    .B(_03914_),
    .Y(_00752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _18327_ (.A1(_02643_),
    .A2(_10822_),
    .B1(_10712_),
    .C1(_10714_),
    .X(_09935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18328_ (.A(_09935_),
    .X(_09936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18329_ (.A(_09936_),
    .Y(_00754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18330_ (.A(_09907_),
    .X(_09937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _18331_ (.A(_03134_),
    .B(_09937_),
    .C(_02855_),
    .X(_00755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18332_ (.A(_03134_),
    .Y(_09938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18333_ (.A(_08325_),
    .X(_09939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18334_ (.A(_09939_),
    .X(_09940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18335_ (.A(_09938_),
    .B(_09940_),
    .Y(_00756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _18336_ (.A(_03127_),
    .B(_09937_),
    .C(_02855_),
    .X(_00758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18337_ (.A(_03127_),
    .Y(_09941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18338_ (.A(_09941_),
    .X(_09942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18339_ (.A(_09942_),
    .B(_09940_),
    .Y(_00759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18340_ (.A(_09811_),
    .X(_09943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _18341_ (.A(_03119_),
    .B(_09943_),
    .C(_02855_),
    .X(_00761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18342_ (.A(_03119_),
    .Y(_09944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18343_ (.A(_09944_),
    .B(_09940_),
    .Y(_00762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _18344_ (.A(_03110_),
    .B(_09943_),
    .C(_02855_),
    .X(_00764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18345_ (.A(_03110_),
    .Y(_09945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18346_ (.A(_09945_),
    .B(_09940_),
    .Y(_00765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _18347_ (.A(_03102_),
    .B(_09943_),
    .C(_09906_),
    .X(_00767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18348_ (.A(_03102_),
    .Y(_09946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18349_ (.A(_09946_),
    .B(_09940_),
    .Y(_00768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _18350_ (.A(_03093_),
    .B(_09943_),
    .C(_09906_),
    .X(_00770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18351_ (.A(_03093_),
    .Y(_09947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18352_ (.A(_09947_),
    .X(_09948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18353_ (.A(_09939_),
    .X(_09949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18354_ (.A(_09948_),
    .B(_09949_),
    .Y(_00771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _18355_ (.A(_03086_),
    .B(_09943_),
    .C(_09906_),
    .X(_00773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18356_ (.A(_03086_),
    .Y(_09950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18357_ (.A(_09950_),
    .X(_09951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18358_ (.A(_09951_),
    .B(_09949_),
    .Y(_00774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _18359_ (.A(_03077_),
    .B(_09907_),
    .C(_09906_),
    .X(_00776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18360_ (.A(_09912_),
    .B(_09949_),
    .Y(_00777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18361_ (.A(\design_top.core0.NXPC[31] ),
    .Y(_00779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18362_ (.A(_08555_),
    .X(_03183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18363_ (.A(_08554_),
    .X(_03181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18364_ (.A(_08536_),
    .X(_03179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18365_ (.A(_08534_),
    .X(_03177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18366_ (.A(_08572_),
    .X(_03171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18367_ (.A(_08594_),
    .X(_03169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18368_ (.A(_08591_),
    .Y(_03168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _18369_ (.A(_08590_),
    .B(_03062_),
    .Y(_03064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18370_ (.A(_08584_),
    .X(_09952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18371_ (.A(_09952_),
    .Y(_03166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _18372_ (.A(_02827_),
    .B(_03078_),
    .Y(_03080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18373_ (.A(_08581_),
    .Y(_03165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _18374_ (.A(_10691_),
    .B(_03094_),
    .Y(_03096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18375_ (.A(_08582_),
    .X(_03164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18376_ (.A(_08587_),
    .Y(_03163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _18377_ (.A(_03111_),
    .B(_02659_),
    .Y(_03113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18378_ (.A(_03128_),
    .X(_09953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _18379_ (.A(_09953_),
    .B(_02641_),
    .Y(_00781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18380_ (.A1(_00688_),
    .A2(_02646_),
    .B1(_08575_),
    .B2(_02649_),
    .X(_09954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18381_ (.A(_09954_),
    .Y(_03162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18382_ (.A(_08578_),
    .Y(_03129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18383_ (.A(_08558_),
    .Y(_03188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18384_ (.A(_02903_),
    .B(_10606_),
    .Y(_02904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _18385_ (.A(_03178_),
    .B(_03177_),
    .C(_03180_),
    .D(_03179_),
    .X(_09955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18386_ (.A(_08544_),
    .X(_01560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _18387_ (.A(_03175_),
    .B(_03174_),
    .C(_01560_),
    .D(_03176_),
    .X(_09956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _18388_ (.A(_03172_),
    .B(_03171_),
    .C(_08565_),
    .D(_03173_),
    .X(_09957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _18389_ (.A(_03168_),
    .B(_03167_),
    .C(_03170_),
    .D(_03169_),
    .X(_09958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18390_ (.A(_08579_),
    .X(_01269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18391_ (.A(_08570_),
    .Y(_01079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18392_ (.A(_03135_),
    .Y(_09959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18393_ (.A(_09959_),
    .B(_03162_),
    .X(_09960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18394_ (.A(_09960_),
    .X(_00938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _18395_ (.A1(_03129_),
    .A2(_00938_),
    .B1(_00781_),
    .X(_09961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18396_ (.A1(_08575_),
    .A2(_02633_),
    .B1(_00688_),
    .B2(_02630_),
    .X(_09962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18397_ (.A(_09962_),
    .Y(_03114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18398_ (.A(_08569_),
    .B(_03114_),
    .X(_09963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18399_ (.A(_09963_),
    .X(_01078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _18400_ (.A1(_01079_),
    .A2(_09961_),
    .B1(_01078_),
    .X(_09964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _18401_ (.A1(_03163_),
    .A2(_09964_),
    .B1(_03113_),
    .X(_09965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _18402_ (.A(_03165_),
    .B(_03164_),
    .C(_09965_),
    .X(_09966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _18403_ (.A1(_03096_),
    .A2(_01181_),
    .B1(_03095_),
    .X(_09967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18404_ (.A(_03087_),
    .B(_10696_),
    .Y(_03088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _18405_ (.A1(_01268_),
    .A2(_09967_),
    .B1(_03088_),
    .C1(_03079_),
    .X(_09968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o311a_2 _18406_ (.A1(_01269_),
    .A2(_03166_),
    .A3(_09966_),
    .B1(_03080_),
    .C1(_09968_),
    .X(_09969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18407_ (.A(_08588_),
    .Y(_03047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _18408_ (.A1(_03064_),
    .A2(_01337_),
    .B1(_03063_),
    .Y(_09970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18409_ (.A(_08593_),
    .B(_09970_),
    .Y(_09971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _18410_ (.A1(_03047_),
    .A2(_03056_),
    .A3(_09971_),
    .B1(_03048_),
    .X(_09972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18411_ (.A(_03030_),
    .B(_08567_),
    .Y(_03031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _18412_ (.A1(_03032_),
    .A2(_01428_),
    .B1(_03031_),
    .X(_09973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18413_ (.A(_03022_),
    .B(_10664_),
    .Y(_03023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18414_ (.A(_03013_),
    .B(_10657_),
    .Y(_03014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _18415_ (.A1(_01476_),
    .A2(_09973_),
    .B1(_03023_),
    .C1(_03014_),
    .X(_09974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _18416_ (.A1(_09957_),
    .A2(_09972_),
    .B1(_03015_),
    .C1(_09974_),
    .X(_09975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _18417_ (.A1(_09957_),
    .A2(_09958_),
    .A3(_09969_),
    .B1(_09975_),
    .X(_09976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18418_ (.A(_02979_),
    .B(_08541_),
    .Y(_02980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18419_ (.A(_02996_),
    .B(_08539_),
    .Y(_02997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _18420_ (.A1(_02998_),
    .A2(_01517_),
    .B1(_02997_),
    .Y(_09977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18421_ (.A(_08543_),
    .B(_09977_),
    .Y(_09978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _18422_ (.A1(_02989_),
    .A2(_02980_),
    .A3(_09978_),
    .B1(_02981_),
    .X(_09979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18423_ (.A(_02962_),
    .B(_08531_),
    .Y(_02963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _18424_ (.A1(_02964_),
    .A2(_01601_),
    .B1(_02963_),
    .X(_09980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18425_ (.A(_08529_),
    .Y(_02946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18426_ (.A(_02954_),
    .B(_10635_),
    .Y(_02955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _18427_ (.A1(_01643_),
    .A2(_09980_),
    .B1(_02946_),
    .C1(_02955_),
    .X(_09981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _18428_ (.A1(_09955_),
    .A2(_09979_),
    .B1(_02947_),
    .C1(_09981_),
    .X(_09982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _18429_ (.A1(_09955_),
    .A2(_09956_),
    .A3(_09976_),
    .B1(_09982_),
    .X(_09983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _18430_ (.A(_03182_),
    .B(_08554_),
    .C(_03184_),
    .D(_03183_),
    .X(_09984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18431_ (.A(_02911_),
    .B(_08549_),
    .Y(_02912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18432_ (.A(_02920_),
    .B(_10619_),
    .Y(_02921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18433_ (.A(_02928_),
    .B(_08551_),
    .Y(_02929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _18434_ (.A1(_02930_),
    .A2(_01683_),
    .B1(_02929_),
    .X(_09985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _18435_ (.A1(_02921_),
    .A2(_09985_),
    .B1(_02913_),
    .C1(_01725_),
    .X(_09986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18436_ (.A1(_09983_),
    .A2(_09984_),
    .B1(_02912_),
    .B2(_09986_),
    .X(_09987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18437_ (.A(_02904_),
    .B(_09987_),
    .X(_09988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18438_ (.A(_02894_),
    .B(_08559_),
    .Y(_02895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _18439_ (.A1(_02896_),
    .A2(_01766_),
    .A3(_09988_),
    .B1(_02895_),
    .X(_09989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _18440_ (.A1(_03187_),
    .A2(_09989_),
    .B1(_02887_),
    .X(_09990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18441_ (.A1_N(_03188_),
    .A2_N(_09990_),
    .B1(_03188_),
    .B2(_09990_),
    .X(_00782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18442_ (.A(_08475_),
    .B(_08492_),
    .Y(_00783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18443_ (.A(_10598_),
    .X(_02879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18444_ (.A1_N(_03139_),
    .A2_N(_02879_),
    .B1(_03139_),
    .B2(_10598_),
    .X(_09991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18445_ (.A(_10604_),
    .X(_02897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18446_ (.A(_03141_),
    .Y(_09992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18447_ (.A1(_03141_),
    .A2(_02897_),
    .B1(_09992_),
    .B2(_10606_),
    .X(_09993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18448_ (.A(_10760_),
    .X(_02888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18449_ (.A(_03140_),
    .Y(_09994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18450_ (.A1(_03140_),
    .A2(_02888_),
    .B1(_09994_),
    .B2(_08559_),
    .X(_09995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18451_ (.A(_03143_),
    .Y(_09996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18452_ (.A1(_03143_),
    .A2(_10756_),
    .B1(_09996_),
    .B2(_10619_),
    .X(_09997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18453_ (.A(_03142_),
    .Y(_09998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18454_ (.A(_09998_),
    .B(_08549_),
    .Y(_09999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _18455_ (.A1(_09998_),
    .A2(_08549_),
    .B1(_09999_),
    .X(_10000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18456_ (.A(_09997_),
    .B(_10000_),
    .X(_10001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18457_ (.A(_03144_),
    .Y(_10002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18458_ (.A(_03145_),
    .Y(_10003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18459_ (.A1(_10003_),
    .A2(_08553_),
    .B1(_10002_),
    .B2(_08551_),
    .X(_10004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _18460_ (.A1(_10002_),
    .A2(_08551_),
    .B1(_10004_),
    .Y(_10005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18461_ (.A(_10633_),
    .X(_10006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18462_ (.A(_03147_),
    .Y(_10007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18463_ (.A1(_03147_),
    .A2(_10006_),
    .B1(_10007_),
    .B2(_10635_),
    .X(_10008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18464_ (.A(_03146_),
    .Y(_10009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18465_ (.A(_10638_),
    .X(_10010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18466_ (.A(_10009_),
    .B(_10010_),
    .Y(_10011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _18467_ (.A1(_10009_),
    .A2(_10010_),
    .B1(_10011_),
    .X(_10012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18468_ (.A(_10008_),
    .B(_10012_),
    .X(_10013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18469_ (.A(_03148_),
    .Y(_10014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18470_ (.A(_03149_),
    .Y(_10015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18471_ (.A1(_10015_),
    .A2(_08533_),
    .B1(_10014_),
    .B2(_08531_),
    .X(_10016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _18472_ (.A1(_10014_),
    .A2(_08531_),
    .B1(_10016_),
    .Y(_10017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18473_ (.A1(_10015_),
    .A2(_08533_),
    .B1(_03149_),
    .B2(_10624_),
    .X(_10018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18474_ (.A1(_03148_),
    .A2(_10628_),
    .B1(_10014_),
    .B2(_08531_),
    .X(_10019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _18475_ (.A(_10018_),
    .B(_10019_),
    .C(_10013_),
    .X(_10020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18476_ (.A(_10644_),
    .X(_10021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18477_ (.A(_03151_),
    .Y(_10022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18478_ (.A1(_03151_),
    .A2(_10021_),
    .B1(_10022_),
    .B2(_02761_),
    .X(_10023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18479_ (.A(_03150_),
    .Y(_10024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18480_ (.A(_10024_),
    .B(_08541_),
    .Y(_10025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _18481_ (.A1(_10024_),
    .A2(_08541_),
    .B1(_10025_),
    .X(_10026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18482_ (.A(_10023_),
    .B(_10026_),
    .X(_10027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18483_ (.A(_03152_),
    .Y(_10028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18484_ (.A(_03153_),
    .Y(_10029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18485_ (.A1(_10029_),
    .A2(_08546_),
    .B1(_10028_),
    .B2(_08539_),
    .X(_10030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _18486_ (.A1(_10028_),
    .A2(_08539_),
    .B1(_10030_),
    .Y(_10031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18487_ (.A(_10736_),
    .X(_10032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18488_ (.A(_10032_),
    .X(_03007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _18489_ (.A1(_03154_),
    .A2(_10032_),
    .B1(_03155_),
    .C1(_10734_),
    .X(_10033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18490_ (.A(_03155_),
    .Y(_10034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18491_ (.A1(_03155_),
    .A2(_10734_),
    .B1(_10034_),
    .B2(_10664_),
    .X(_10035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18492_ (.A1_N(_03154_),
    .A2_N(_10032_),
    .B1(_03154_),
    .B2(_10032_),
    .X(_10036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18493_ (.A(_10035_),
    .B(_10036_),
    .X(_10037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18494_ (.A(_03156_),
    .Y(_10038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _18495_ (.A1(_03156_),
    .A2(_10667_),
    .B1(_03157_),
    .B2(_10670_),
    .Y(_10039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _18496_ (.A1(_10038_),
    .A2(_08567_),
    .B1(_10039_),
    .Y(_10040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18497_ (.A(_10037_),
    .B(_10040_),
    .X(_10041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18498_ (.A(_10667_),
    .X(_03024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18499_ (.A1(_10038_),
    .A2(_08567_),
    .B1(_03156_),
    .B2(_03024_),
    .X(_10042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18500_ (.A(_10670_),
    .X(_10043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18501_ (.A1_N(_03157_),
    .A2_N(_10043_),
    .B1(_03157_),
    .B2(_10043_),
    .X(_10044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18502_ (.A(_10699_),
    .X(_00809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18503_ (.A(_03111_),
    .X(_10045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18504_ (.A(_08586_),
    .Y(_03105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _18505_ (.A1(_03111_),
    .A2(_08586_),
    .B1(_03113_),
    .X(_10046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18506_ (.A(_08576_),
    .Y(_03122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18507_ (.A(_09959_),
    .B(_02650_),
    .Y(_10047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18508_ (.A1(_03128_),
    .A2(_03122_),
    .B1(_08577_),
    .B2(_10047_),
    .X(_10048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _18509_ (.A1(_03120_),
    .A2(_09962_),
    .B1(_01078_),
    .X(_10049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18510_ (.A1(_03120_),
    .A2(_03114_),
    .B1(_10048_),
    .B2(_10049_),
    .X(_10050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18511_ (.A1(_10045_),
    .A2(_03105_),
    .B1(_10046_),
    .B2(_10050_),
    .X(_10051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _18512_ (.A1(_03103_),
    .A2(_10694_),
    .A3(_08581_),
    .B1(_00811_),
    .B2(_03094_),
    .X(_10052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18513_ (.A1(_03087_),
    .A2(_03081_),
    .B1(_08580_),
    .B2(_10052_),
    .X(_10053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18514_ (.A(_09952_),
    .B(_10053_),
    .X(_10054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _18515_ (.A1(_00809_),
    .A2(_03078_),
    .B1(_08585_),
    .B2(_10051_),
    .C1(_10054_),
    .X(_10055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18516_ (.A(_10727_),
    .X(_03065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _18517_ (.A1(_03071_),
    .A2(_03065_),
    .A3(_08591_),
    .B1(_00805_),
    .B2(_03062_),
    .X(_10056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18518_ (.A1(_03055_),
    .A2(_03049_),
    .B1(_08595_),
    .B2(_10056_),
    .X(_10057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18519_ (.A(_08589_),
    .B(_10057_),
    .X(_10058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _18520_ (.A1(_00803_),
    .A2(_03046_),
    .B1(_08596_),
    .B2(_10055_),
    .C1(_10058_),
    .X(_10059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _18521_ (.A(_10042_),
    .B(_10044_),
    .C(_10037_),
    .D(_10059_),
    .X(_10060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2111a_2 _18522_ (.A1(_03154_),
    .A2(_03007_),
    .B1(_10033_),
    .C1(_10041_),
    .D1(_10060_),
    .X(_10061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18523_ (.A1(_10029_),
    .A2(_08546_),
    .B1(_03153_),
    .B2(_10740_),
    .X(_10062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18524_ (.A1(_03152_),
    .A2(_10743_),
    .B1(_10028_),
    .B2(_08539_),
    .X(_10063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _18525_ (.A(_10062_),
    .B(_10063_),
    .C(_10027_),
    .X(_10064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18526_ (.A(_10654_),
    .X(_02973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _18527_ (.A1(_03151_),
    .A2(_10021_),
    .A3(_10025_),
    .B1(_03150_),
    .B2(_02973_),
    .X(_10065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _18528_ (.A1(_10027_),
    .A2(_10031_),
    .B1(_10061_),
    .B2(_10064_),
    .C1(_10065_),
    .X(_10066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _18529_ (.A1(_03147_),
    .A2(_10006_),
    .A3(_10011_),
    .B1(_03146_),
    .B2(_02939_),
    .X(_10067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _18530_ (.A1(_10013_),
    .A2(_10017_),
    .B1(_10020_),
    .B2(_10066_),
    .C1(_10067_),
    .X(_10068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18531_ (.A1(_03145_),
    .A2(_10613_),
    .B1(_10003_),
    .B2(_08553_),
    .X(_10069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18532_ (.A(_10609_),
    .X(_02922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18533_ (.A1(_03144_),
    .A2(_02922_),
    .B1(_10002_),
    .B2(_08551_),
    .X(_10070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _18534_ (.A(_10069_),
    .B(_10070_),
    .C(_10001_),
    .X(_10071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18535_ (.A(_10756_),
    .X(_02914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18536_ (.A(_10617_),
    .X(_02905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _18537_ (.A1(_03143_),
    .A2(_02914_),
    .A3(_09999_),
    .B1(_03142_),
    .B2(_02905_),
    .X(_10072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _18538_ (.A1(_10001_),
    .A2(_10005_),
    .B1(_10068_),
    .B2(_10071_),
    .C1(_10072_),
    .X(_10073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18539_ (.A1(_09992_),
    .A2(_10606_),
    .B1(_09994_),
    .B2(_08559_),
    .X(_10074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _18540_ (.A1(_09994_),
    .A2(_08559_),
    .B1(_10074_),
    .Y(_10075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _18541_ (.A1(_09993_),
    .A2(_09995_),
    .A3(_10073_),
    .B1(_10075_),
    .X(_10076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _18542_ (.A1(_03139_),
    .A2(_02879_),
    .B1(_09991_),
    .B2(_10076_),
    .Y(_10077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18543_ (.A(_10764_),
    .X(_10078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18544_ (.A(_03138_),
    .Y(_10079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18545_ (.A(_10078_),
    .B(_10079_),
    .Y(_10080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _18546_ (.A1(_10078_),
    .A2(_10079_),
    .B1(_10080_),
    .Y(_10081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18547_ (.A1_N(_10077_),
    .A2_N(_10081_),
    .B1(_10077_),
    .B2(_10081_),
    .X(_00784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18548_ (.A(\design_top.core0.REG1[14][31] ),
    .Y(_02681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18549_ (.A(_03135_),
    .X(_10082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18550_ (.A(_02684_),
    .X(_10083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18551_ (.A(_10082_),
    .B(_10083_),
    .X(_00820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18552_ (.A(_09953_),
    .B(_00820_),
    .X(_00821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18553_ (.A(_03120_),
    .X(_10084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18554_ (.A(_10084_),
    .X(_10085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18555_ (.A(_10085_),
    .B(_00821_),
    .X(_00822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18556_ (.A(_10045_),
    .X(_10086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18557_ (.A(_10086_),
    .B(_00822_),
    .X(_00823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18558_ (.A(_03103_),
    .X(_10087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18559_ (.A(_10087_),
    .X(_10088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18560_ (.A(_10088_),
    .B(_00823_),
    .X(_00824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18561_ (.A(\design_top.core0.REG1[15][31] ),
    .Y(_02682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _18562_ (.A(\design_top.core0.FCT3[1] ),
    .B(_09914_),
    .C(_08599_),
    .X(_10089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18563_ (.A(_10089_),
    .X(_10090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18564_ (.A(_10090_),
    .X(_00827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _18565_ (.A(_08502_),
    .B(\design_top.core0.FCT3[0] ),
    .C(_08599_),
    .X(_10091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18566_ (.A(_10091_),
    .X(_10092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18567_ (.A(_10092_),
    .X(_00828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _18568_ (.A(_00826_),
    .B(_00827_),
    .C(_00828_),
    .X(_00829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18569_ (.A(\design_top.RAMFF[31] ),
    .Y(_00832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18570_ (.A(\design_top.XADDR[2] ),
    .B(\design_top.XADDR[3] ),
    .Y(_00833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18571_ (.A(\design_top.IOMUX[3][31] ),
    .Y(_10093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18572_ (.A(\design_top.XADDR[2] ),
    .Y(_00994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18573_ (.A(\design_top.XADDR[3] ),
    .Y(_10094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18574_ (.A(_00994_),
    .B(_10094_),
    .X(_10095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18575_ (.A(_10095_),
    .X(_10096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18576_ (.A(_10096_),
    .X(_10097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18577_ (.A(\design_top.GPIOFF[15] ),
    .Y(_10098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18578_ (.A(\design_top.XADDR[2] ),
    .B(_10094_),
    .X(_10099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18579_ (.A(_10099_),
    .X(_10100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18580_ (.A(_10100_),
    .X(_10101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18581_ (.A1(_10093_),
    .A2(_10097_),
    .B1(_10098_),
    .B2(_10101_),
    .X(_00834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18582_ (.A(\design_top.RAMFF[15] ),
    .Y(_00837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18583_ (.A(\design_top.IOMUX[3][15] ),
    .Y(_10102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18584_ (.A(_10095_),
    .X(_10103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18585_ (.A(\design_top.LEDFF[15] ),
    .Y(_10104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18586_ (.A(_10099_),
    .X(_10105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18587_ (.A(_00994_),
    .B(\design_top.XADDR[3] ),
    .Y(_10106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18588_ (.A(_10106_),
    .X(_10107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _18589_ (.A(\design_top.uart0.UART_RFIFO[7] ),
    .B(_10107_),
    .Y(_10108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _18590_ (.A1(_10102_),
    .A2(_10103_),
    .B1(_10104_),
    .B2(_10105_),
    .C1(_10108_),
    .X(_00838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _18591_ (.A(_09913_),
    .B(_09915_),
    .C(_00840_),
    .X(_00841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18592_ (.A(\design_top.RAMFF[23] ),
    .Y(_00843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18593_ (.A(\design_top.IOMUX[3][23] ),
    .Y(_10109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18594_ (.A(\design_top.GPIOFF[7] ),
    .Y(_10110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18595_ (.A1(_10109_),
    .A2(_10097_),
    .B1(_10110_),
    .B2(_10101_),
    .X(_00844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18596_ (.A(\design_top.RAMFF[7] ),
    .Y(_00846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18597_ (.A(\design_top.IOMUX[3][7] ),
    .Y(_10111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18598_ (.A(\design_top.LEDFF[7] ),
    .Y(_10112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18599_ (.A1(_10111_),
    .A2(_10097_),
    .B1(_10112_),
    .B2(_10101_),
    .X(_00847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _18600_ (.A(_09913_),
    .B(_02854_),
    .C(_00851_),
    .X(_00852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _18601_ (.A(_10590_),
    .B(_10591_),
    .C(\design_top.core0.XLUI ),
    .X(_00854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18602_ (.A(\design_top.core0.REG1[13][31] ),
    .Y(_02680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _18603_ (.A(_10590_),
    .B(_10591_),
    .C(\design_top.core0.XAUIPC ),
    .X(_00857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18604_ (.A(\design_top.core0.PC[30] ),
    .Y(_10113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18605_ (.A1(\design_top.core0.SIMM[30] ),
    .A2(\design_top.core0.PC[30] ),
    .B1(_02690_),
    .B2(_10113_),
    .X(_10114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18606_ (.A(_10600_),
    .B(\design_top.core0.PC[29] ),
    .Y(_10115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18607_ (.A(_10605_),
    .B(\design_top.core0.PC[28] ),
    .Y(_10116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18608_ (.A(\design_top.core0.PC[27] ),
    .Y(_10117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18609_ (.A(_10620_),
    .X(_02714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18610_ (.A(\design_top.core0.PC[26] ),
    .Y(_10118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _18611_ (.A1(_02708_),
    .A2(_10117_),
    .B1(_02714_),
    .C1(_10118_),
    .X(_10119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18612_ (.A1(\design_top.core0.SIMM[27] ),
    .A2(\design_top.core0.PC[27] ),
    .B1(_02708_),
    .B2(_10117_),
    .X(_10120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18613_ (.A1(\design_top.core0.SIMM[26] ),
    .A2(\design_top.core0.PC[26] ),
    .B1(_02714_),
    .B2(_10118_),
    .X(_10121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18614_ (.A(_10120_),
    .B(_10121_),
    .X(_10122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18615_ (.A1(_08457_),
    .A2(\design_top.core0.PC[25] ),
    .B1(_08460_),
    .B2(\design_top.core0.PC[24] ),
    .X(_10123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _18616_ (.A1(_08457_),
    .A2(\design_top.core0.PC[25] ),
    .B1(_10123_),
    .Y(_10124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18617_ (.A(_10122_),
    .B(_10124_),
    .X(_10125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18618_ (.A1_N(_08457_),
    .A2_N(\design_top.core0.PC[25] ),
    .B1(_08457_),
    .B2(\design_top.core0.PC[25] ),
    .X(_10126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18619_ (.A(_10126_),
    .Y(_10127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18620_ (.A1_N(_08460_),
    .A2_N(\design_top.core0.PC[24] ),
    .B1(_08460_),
    .B2(\design_top.core0.PC[24] ),
    .X(_10128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18621_ (.A(_10128_),
    .Y(_10129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18622_ (.A(_10653_),
    .B(\design_top.core0.PC[19] ),
    .X(_10130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _18623_ (.A1(_10653_),
    .A2(\design_top.core0.PC[19] ),
    .B1_N(_10130_),
    .X(_10131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18624_ (.A(_10131_),
    .Y(_10132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18625_ (.A(\design_top.core0.PC[18] ),
    .Y(_10133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18626_ (.A1(_02762_),
    .A2(_10133_),
    .B1(\design_top.core0.SIMM[18] ),
    .B2(\design_top.core0.PC[18] ),
    .X(_10134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18627_ (.A1_N(_08466_),
    .A2_N(\design_top.core0.PC[17] ),
    .B1(_08466_),
    .B2(\design_top.core0.PC[17] ),
    .X(_10135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18628_ (.A1_N(_08467_),
    .A2_N(\design_top.core0.PC[16] ),
    .B1(_08467_),
    .B2(\design_top.core0.PC[16] ),
    .X(_10136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and4_2 _18629_ (.A(_10132_),
    .B(_10134_),
    .C(_10135_),
    .D(_10136_),
    .X(_10137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18630_ (.A1_N(_08462_),
    .A2_N(\design_top.core0.PC[21] ),
    .B1(_08462_),
    .B2(\design_top.core0.PC[21] ),
    .X(_10138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18631_ (.A(_10138_),
    .Y(_10139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18632_ (.A(\design_top.core0.PC[20] ),
    .Y(_10140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18633_ (.A1(_02750_),
    .A2(_10140_),
    .B1(_10625_),
    .B2(\design_top.core0.PC[20] ),
    .X(_10141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18634_ (.A(_10141_),
    .Y(_10142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18635_ (.A(\design_top.core0.PC[22] ),
    .Y(_10143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18636_ (.A1(_10634_),
    .A2(\design_top.core0.PC[22] ),
    .B1(_02738_),
    .B2(_10143_),
    .X(_10144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18637_ (.A(\design_top.core0.PC[23] ),
    .Y(_10145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18638_ (.A1(_10750_),
    .A2(\design_top.core0.PC[23] ),
    .B1(_02732_),
    .B2(_10145_),
    .X(_10146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor4_2 _18639_ (.A(_10139_),
    .B(_10142_),
    .C(_10144_),
    .D(_10146_),
    .Y(_10147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18640_ (.A(_10688_),
    .B(\design_top.core0.PC[11] ),
    .X(_10148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _18641_ (.A1(_10688_),
    .A2(\design_top.core0.PC[11] ),
    .B1_N(_10148_),
    .X(_10149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18642_ (.A(_10149_),
    .Y(_10150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18643_ (.A(\design_top.core0.PC[10] ),
    .Y(_10151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18644_ (.A1(_02810_),
    .A2(_10151_),
    .B1(\design_top.core0.SIMM[10] ),
    .B2(\design_top.core0.PC[10] ),
    .X(_10152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18645_ (.A1_N(_08437_),
    .A2_N(\design_top.core0.PC[9] ),
    .B1(_08437_),
    .B2(\design_top.core0.PC[9] ),
    .X(_10153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18646_ (.A1_N(_08441_),
    .A2_N(\design_top.core0.PC[8] ),
    .B1(_08441_),
    .B2(\design_top.core0.PC[8] ),
    .X(_10154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and4_2 _18647_ (.A(_10150_),
    .B(_10152_),
    .C(_10153_),
    .D(_10154_),
    .X(_10155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18648_ (.A1_N(_08472_),
    .A2_N(\design_top.core0.PC[13] ),
    .B1(_08472_),
    .B2(\design_top.core0.PC[13] ),
    .X(_10156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18649_ (.A(_10156_),
    .Y(_10157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18650_ (.A(\design_top.core0.PC[12] ),
    .Y(_10158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18651_ (.A1(_02798_),
    .A2(_10158_),
    .B1(_10671_),
    .B2(\design_top.core0.PC[12] ),
    .X(_10159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18652_ (.A(_10159_),
    .Y(_10160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18653_ (.A(\design_top.core0.PC[14] ),
    .Y(_10161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18654_ (.A1(_10663_),
    .A2(\design_top.core0.PC[14] ),
    .B1(_02786_),
    .B2(_10161_),
    .X(_10162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18655_ (.A(\design_top.core0.PC[15] ),
    .Y(_10163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18656_ (.A1(_10735_),
    .A2(\design_top.core0.PC[15] ),
    .B1(_02780_),
    .B2(_10163_),
    .X(_10164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor4_2 _18657_ (.A(_10157_),
    .B(_10160_),
    .C(_10162_),
    .D(_10164_),
    .Y(_10165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18658_ (.A1_N(_08443_),
    .A2_N(\design_top.core0.PC[7] ),
    .B1(_08443_),
    .B2(\design_top.core0.PC[7] ),
    .X(_10166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18659_ (.A1_N(_08444_),
    .A2_N(\design_top.core0.PC[6] ),
    .B1(_08444_),
    .B2(\design_top.core0.PC[6] ),
    .X(_10167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18660_ (.A1_N(_08445_),
    .A2_N(\design_top.core0.PC[5] ),
    .B1(_08445_),
    .B2(\design_top.core0.PC[5] ),
    .X(_10168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18661_ (.A1_N(_08447_),
    .A2_N(\design_top.core0.PC[4] ),
    .B1(_08447_),
    .B2(\design_top.core0.PC[4] ),
    .X(_10169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18662_ (.A(_10702_),
    .B(\design_top.core0.PC[3] ),
    .Y(_10170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18663_ (.A(_10706_),
    .B(\design_top.core0.PC[2] ),
    .Y(_10171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18664_ (.A1_N(_10709_),
    .A2_N(\design_top.core0.PC[1] ),
    .B1(_10709_),
    .B2(\design_top.core0.PC[1] ),
    .X(_10172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18665_ (.A(\design_top.core0.PC[0] ),
    .Y(_10173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18666_ (.A(_10710_),
    .B(_10173_),
    .Y(_10174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18667_ (.A1(_10709_),
    .A2(\design_top.core0.PC[1] ),
    .B1(_10172_),
    .B2(_10174_),
    .X(_10175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18668_ (.A(_10175_),
    .Y(_10176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18669_ (.A1_N(_10706_),
    .A2_N(\design_top.core0.PC[2] ),
    .B1(_10171_),
    .B2(_10176_),
    .X(_10177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2ai_2 _18670_ (.A1_N(_10702_),
    .A2_N(\design_top.core0.PC[3] ),
    .B1(_10170_),
    .B2(_10177_),
    .Y(_10178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18671_ (.A(_08445_),
    .B(\design_top.core0.PC[5] ),
    .X(_10179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a32o_2 _18672_ (.A1(_08447_),
    .A2(\design_top.core0.PC[4] ),
    .A3(_10179_),
    .B1(_08445_),
    .B2(\design_top.core0.PC[5] ),
    .X(_10180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _18673_ (.A1(_10168_),
    .A2(_10169_),
    .A3(_10178_),
    .B1(_10180_),
    .X(_10181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18674_ (.A(_08443_),
    .B(\design_top.core0.PC[7] ),
    .X(_10182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a32o_2 _18675_ (.A1(_08444_),
    .A2(\design_top.core0.PC[6] ),
    .A3(_10182_),
    .B1(_08443_),
    .B2(\design_top.core0.PC[7] ),
    .X(_10183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _18676_ (.A1(_10166_),
    .A2(_10167_),
    .A3(_10181_),
    .B1(_10183_),
    .X(_10184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18677_ (.A1(_08437_),
    .A2(\design_top.core0.PC[9] ),
    .B1(_08441_),
    .B2(\design_top.core0.PC[8] ),
    .X(_10185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _18678_ (.A1(_08437_),
    .A2(\design_top.core0.PC[9] ),
    .B1(_10185_),
    .X(_10186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a32o_2 _18679_ (.A1(\design_top.core0.SIMM[10] ),
    .A2(\design_top.core0.PC[10] ),
    .A3(_10148_),
    .B1(_10688_),
    .B2(\design_top.core0.PC[11] ),
    .X(_10187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _18680_ (.A1(_10150_),
    .A2(_10152_),
    .A3(_10186_),
    .B1(_10187_),
    .X(_10188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18681_ (.A1(_08472_),
    .A2(\design_top.core0.PC[13] ),
    .B1(_10671_),
    .B2(\design_top.core0.PC[12] ),
    .X(_10189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _18682_ (.A1(_08472_),
    .A2(\design_top.core0.PC[13] ),
    .B1(_10189_),
    .X(_10190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _18683_ (.A1(_10156_),
    .A2(_10159_),
    .A3(_10188_),
    .B1(_10190_),
    .X(_10191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _18684_ (.A1(_10663_),
    .A2(\design_top.core0.PC[14] ),
    .B1(_10191_),
    .X(_10192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18685_ (.A1(_10663_),
    .A2(\design_top.core0.PC[14] ),
    .B1(_10735_),
    .B2(\design_top.core0.PC[15] ),
    .X(_10193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18686_ (.A1(_10735_),
    .A2(\design_top.core0.PC[15] ),
    .B1(_10192_),
    .B2(_10193_),
    .X(_10194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _18687_ (.A1(_10155_),
    .A2(_10165_),
    .A3(_10184_),
    .B1(_10194_),
    .X(_10195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18688_ (.A1(_08466_),
    .A2(\design_top.core0.PC[17] ),
    .B1(_08467_),
    .B2(\design_top.core0.PC[16] ),
    .X(_10196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _18689_ (.A1(_08466_),
    .A2(\design_top.core0.PC[17] ),
    .B1(_10196_),
    .X(_10197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a32o_2 _18690_ (.A1(\design_top.core0.SIMM[18] ),
    .A2(\design_top.core0.PC[18] ),
    .A3(_10130_),
    .B1(_10653_),
    .B2(\design_top.core0.PC[19] ),
    .X(_10198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _18691_ (.A1(_10132_),
    .A2(_10134_),
    .A3(_10197_),
    .B1(_10198_),
    .X(_10199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18692_ (.A1(_08462_),
    .A2(\design_top.core0.PC[21] ),
    .B1(_10625_),
    .B2(\design_top.core0.PC[20] ),
    .X(_10200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _18693_ (.A1(_08462_),
    .A2(\design_top.core0.PC[21] ),
    .B1(_10200_),
    .X(_10201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _18694_ (.A1(_10138_),
    .A2(_10141_),
    .A3(_10199_),
    .B1(_10201_),
    .X(_10202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _18695_ (.A1(_10634_),
    .A2(\design_top.core0.PC[22] ),
    .B1(_10202_),
    .X(_10203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18696_ (.A1(_10634_),
    .A2(\design_top.core0.PC[22] ),
    .B1(_10750_),
    .B2(\design_top.core0.PC[23] ),
    .X(_10204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18697_ (.A1(_10750_),
    .A2(\design_top.core0.PC[23] ),
    .B1(_10203_),
    .B2(_10204_),
    .X(_10205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _18698_ (.A1(_10137_),
    .A2(_10147_),
    .A3(_10195_),
    .B1(_10205_),
    .X(_10206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18699_ (.A(_10206_),
    .Y(_10207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _18700_ (.A(_10127_),
    .B(_10129_),
    .C(_10122_),
    .D(_10207_),
    .X(_10208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2111a_2 _18701_ (.A1(_02708_),
    .A2(_10117_),
    .B1(_10119_),
    .C1(_10125_),
    .D1(_10208_),
    .X(_10209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18702_ (.A1_N(_10605_),
    .A2_N(\design_top.core0.PC[28] ),
    .B1(_10116_),
    .B2(_10209_),
    .X(_10210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18703_ (.A1_N(_10600_),
    .A2_N(\design_top.core0.PC[29] ),
    .B1(_10115_),
    .B2(_10210_),
    .X(_10211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _18704_ (.A1(_02690_),
    .A2(_10113_),
    .B1(_10114_),
    .B2(_10211_),
    .Y(_10212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18705_ (.A1_N(_00780_),
    .A2_N(\design_top.core0.PC[31] ),
    .B1(_00780_),
    .B2(\design_top.core0.PC[31] ),
    .X(_10213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18706_ (.A1_N(_10212_),
    .A2_N(_10213_),
    .B1(_10212_),
    .B2(_10213_),
    .X(_00858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18707_ (.A(_09935_),
    .X(_02856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18708_ (.A(_09938_),
    .B(_02856_),
    .Y(_00864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18709_ (.A(_03070_),
    .Y(_10214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18710_ (.A(_10214_),
    .B(_09949_),
    .Y(_00865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18711_ (.A(_09942_),
    .B(_02856_),
    .Y(_00867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18712_ (.A(_03061_),
    .Y(_10215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18713_ (.A(_10215_),
    .B(_09949_),
    .Y(_00868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18714_ (.A(_09944_),
    .B(_02856_),
    .Y(_00870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18715_ (.A(_03054_),
    .Y(_10216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18716_ (.A(_09939_),
    .X(_10217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18717_ (.A(_10216_),
    .B(_10217_),
    .Y(_00871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18718_ (.A(_09945_),
    .B(_02856_),
    .Y(_00873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18719_ (.A(_03045_),
    .Y(_10218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18720_ (.A(_10218_),
    .B(_10217_),
    .Y(_00874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18721_ (.A(_09946_),
    .B(_09936_),
    .Y(_00876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18722_ (.A(_03038_),
    .Y(_10219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18723_ (.A(_10219_),
    .B(_10217_),
    .Y(_00877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18724_ (.A(_09948_),
    .B(_09936_),
    .Y(_00879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18725_ (.A(_03029_),
    .Y(_10220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18726_ (.A(_10220_),
    .B(_10217_),
    .Y(_00880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18727_ (.A(_09951_),
    .B(_09936_),
    .Y(_00882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18728_ (.A(_03021_),
    .Y(_10221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18729_ (.A(_10221_),
    .B(_10217_),
    .Y(_00883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18730_ (.A(_09912_),
    .B(_09936_),
    .Y(_00885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18731_ (.A(_09916_),
    .B(_09939_),
    .Y(_00886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18732_ (.A(_09812_),
    .X(_02864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18733_ (.A(_09938_),
    .B(_02864_),
    .Y(_00888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18734_ (.A(_09938_),
    .B(_02850_),
    .Y(_00889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18735_ (.A(_09942_),
    .B(_02864_),
    .Y(_00891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18736_ (.A(_09942_),
    .B(_02850_),
    .Y(_00892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18737_ (.A(_09944_),
    .B(_02864_),
    .Y(_00894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18738_ (.A(_09944_),
    .B(_02850_),
    .Y(_00895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18739_ (.A(_09945_),
    .B(_02864_),
    .Y(_00897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18740_ (.A(_09907_),
    .X(_10222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18741_ (.A(_09945_),
    .B(_10222_),
    .Y(_00898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18742_ (.A(_09946_),
    .B(_09908_),
    .Y(_00900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18743_ (.A(_09946_),
    .B(_10222_),
    .Y(_00901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18744_ (.A(_09948_),
    .B(_09908_),
    .Y(_00903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18745_ (.A(_09948_),
    .B(_10222_),
    .Y(_00904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18746_ (.A(_09951_),
    .B(_09908_),
    .Y(_00906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18747_ (.A(_09951_),
    .B(_10222_),
    .Y(_00907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18748_ (.A(_09912_),
    .B(_09908_),
    .Y(_00909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18749_ (.A(_09912_),
    .B(_10222_),
    .Y(_00910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18750_ (.A(_09938_),
    .B(_02867_),
    .Y(_00912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18751_ (.A(_09907_),
    .X(_10223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18752_ (.A(_10214_),
    .B(_10223_),
    .Y(_00913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18753_ (.A(_09942_),
    .B(_02867_),
    .Y(_00915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18754_ (.A(_10215_),
    .B(_10223_),
    .Y(_00916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18755_ (.A(_09944_),
    .B(_02867_),
    .Y(_00918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18756_ (.A(_10216_),
    .B(_10223_),
    .Y(_00919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18757_ (.A(_09945_),
    .B(_09911_),
    .Y(_00921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18758_ (.A(_10218_),
    .B(_10223_),
    .Y(_00922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18759_ (.A(_09946_),
    .B(_09911_),
    .Y(_00924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18760_ (.A(_10219_),
    .B(_10223_),
    .Y(_00925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18761_ (.A(_09948_),
    .B(_09911_),
    .Y(_00927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18762_ (.A(_10220_),
    .B(_09937_),
    .Y(_00928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18763_ (.A(_09951_),
    .B(_09911_),
    .Y(_00930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18764_ (.A(_10221_),
    .B(_09937_),
    .Y(_00931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18765_ (.A(\design_top.core0.RESMODE[1] ),
    .Y(_10224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18766_ (.A(_08669_),
    .B(_10224_),
    .Y(_00933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18767_ (.A(_03195_),
    .Y(_00935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18768_ (.A(_10590_),
    .B(_10591_),
    .Y(_00936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18769_ (.A(\design_top.core0.NXPC[0] ),
    .Y(_00937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _18770_ (.A(_10082_),
    .B(_09954_),
    .Y(_00939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18771_ (.A(_10082_),
    .B(_03162_),
    .X(_00941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18772_ (.A(_09953_),
    .B(_00941_),
    .X(_00942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18773_ (.A(_10085_),
    .B(_00942_),
    .X(_00943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18774_ (.A(_10086_),
    .B(_00943_),
    .X(_00944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18775_ (.A(_10088_),
    .B(_00944_),
    .X(_00945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18776_ (.A(_00976_),
    .X(_00977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18777_ (.A(\design_top.RAMFF[0] ),
    .Y(_00984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18778_ (.A1_N(\design_top.uart0.UART_XACK ),
    .A2_N(\design_top.uart0.UART_XREQ ),
    .B1(\design_top.uart0.UART_XACK ),
    .B2(\design_top.uart0.UART_XREQ ),
    .X(_00985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18779_ (.A(\design_top.IOMUX[3][0] ),
    .Y(_10225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18780_ (.A(io_out[8]),
    .Y(_10226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _18781_ (.A(_00994_),
    .B(\design_top.XADDR[3] ),
    .C(_00985_),
    .X(_10227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _18782_ (.A1(_10225_),
    .A2(_10103_),
    .B1(_10226_),
    .B2(_10105_),
    .C1(_10227_),
    .X(_00986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18783_ (.A(\design_top.RAMFF[16] ),
    .Y(_00988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18784_ (.A(\design_top.IOMUX[3][16] ),
    .Y(_10228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18785_ (.A(io_out[15]),
    .Y(_10229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18786_ (.A1(_10228_),
    .A2(_10097_),
    .B1(_10229_),
    .B2(_10101_),
    .X(_00989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18787_ (.A(\design_top.RAMFF[24] ),
    .Y(_00993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18788_ (.A(\design_top.IOMUX[3][24] ),
    .Y(_10230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18789_ (.A(\design_top.GPIOFF[8] ),
    .Y(_10231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18790_ (.A1(_10230_),
    .A2(_10097_),
    .B1(_10231_),
    .B2(_10101_),
    .X(_00995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18791_ (.A(\design_top.RAMFF[8] ),
    .Y(_00998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18792_ (.A(\design_top.IOMUX[3][8] ),
    .Y(_10232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18793_ (.A(\design_top.LEDFF[8] ),
    .Y(_10233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _18794_ (.A(\design_top.uart0.UART_RFIFO[0] ),
    .B(_10107_),
    .Y(_10234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _18795_ (.A1(_10232_),
    .A2(_10103_),
    .B1(_10233_),
    .B2(_10105_),
    .C1(_10234_),
    .X(_00999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _18796_ (.A1(_02643_),
    .A2(_10173_),
    .B1(_10174_),
    .X(_01007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18797_ (.A(\design_top.core0.REG1[12][31] ),
    .Y(_02679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18798_ (.A(\design_top.core0.NXPC[1] ),
    .Y(_01009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a32o_2 _18799_ (.A1(_10082_),
    .A2(_09954_),
    .A3(_08578_),
    .B1(_03129_),
    .B2(_00938_),
    .X(_01011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18800_ (.A1_N(_08578_),
    .A2_N(_10047_),
    .B1(_08578_),
    .B2(_10047_),
    .X(_01012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18801_ (.A(\design_top.core0.REG1[11][31] ),
    .Y(_02677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18802_ (.A(_09953_),
    .B(_00815_),
    .X(_01013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18803_ (.A(_10085_),
    .B(_01013_),
    .X(_01014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18804_ (.A(_10086_),
    .B(_01014_),
    .X(_01015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18805_ (.A(_10088_),
    .B(_01015_),
    .X(_01016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18806_ (.A(\design_top.core0.REG1[10][31] ),
    .Y(_02676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _18807_ (.A(_01050_),
    .B(_00827_),
    .C(_00828_),
    .X(_01051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18808_ (.A(\design_top.RAMFF[1] ),
    .Y(_01054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18809_ (.A(\design_top.IOMUX[3][1] ),
    .Y(_10235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18810_ (.A(_10095_),
    .X(_10236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18811_ (.A(io_out[9]),
    .Y(_10237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18812_ (.A(_10099_),
    .X(_10238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _18813_ (.A1(\design_top.uart0.UART_RREQ ),
    .A2(\design_top.uart0.UART_RACK ),
    .B1(_10106_),
    .Y(_10239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _18814_ (.A1(\design_top.uart0.UART_RREQ ),
    .A2(\design_top.uart0.UART_RACK ),
    .B1(_10239_),
    .X(_10240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _18815_ (.A1(_10235_),
    .A2(_10236_),
    .B1(_10237_),
    .B2(_10238_),
    .C1(_10240_),
    .X(_01055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18816_ (.A(\design_top.RAMFF[17] ),
    .Y(_01057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18817_ (.A(\design_top.IOMUX[3][17] ),
    .Y(_10241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18818_ (.A(_10096_),
    .X(_10242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18819_ (.A(\design_top.GPIOFF[1] ),
    .Y(_10243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18820_ (.A(_10100_),
    .X(_10244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18821_ (.A1(_10241_),
    .A2(_10242_),
    .B1(_10243_),
    .B2(_10244_),
    .X(_01058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18822_ (.A(\design_top.RAMFF[25] ),
    .Y(_01062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18823_ (.A(\design_top.IOMUX[3][25] ),
    .Y(_10245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18824_ (.A(\design_top.GPIOFF[9] ),
    .Y(_10246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18825_ (.A1(_10245_),
    .A2(_10242_),
    .B1(_10246_),
    .B2(_10244_),
    .X(_01063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18826_ (.A(\design_top.RAMFF[9] ),
    .Y(_01066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18827_ (.A(\design_top.IOMUX[3][9] ),
    .Y(_10247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18828_ (.A(\design_top.LEDFF[9] ),
    .Y(_10248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _18829_ (.A(\design_top.uart0.UART_RFIFO[1] ),
    .B(_10107_),
    .Y(_10249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _18830_ (.A1(_10247_),
    .A2(_10236_),
    .B1(_10248_),
    .B2(_10238_),
    .C1(_10249_),
    .X(_01067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18831_ (.A(\design_top.core0.REG1[8][31] ),
    .Y(_02674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2ai_2 _18832_ (.A1_N(_10172_),
    .A2_N(_10174_),
    .B1(_10172_),
    .B2(_10174_),
    .Y(_01075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18833_ (.A(\design_top.core0.REG1[9][31] ),
    .Y(_02675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18834_ (.A(\design_top.core0.NXPC[2] ),
    .Y(_01077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18835_ (.A1_N(_01079_),
    .A2_N(_09961_),
    .B1(_01079_),
    .B2(_09961_),
    .X(_01080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18836_ (.A1_N(_10048_),
    .A2_N(_10049_),
    .B1(_10048_),
    .B2(_10049_),
    .X(_01081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18837_ (.A(_10085_),
    .B(_01083_),
    .X(_01084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18838_ (.A(_10086_),
    .B(_01084_),
    .X(_01085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18839_ (.A(_10088_),
    .B(_01085_),
    .X(_01086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18840_ (.A(_09953_),
    .B(_00972_),
    .X(_01098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18841_ (.A(\design_top.core0.REG1[7][31] ),
    .Y(_02672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _18842_ (.A(_01105_),
    .B(_00827_),
    .C(_00828_),
    .X(_01106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18843_ (.A(\design_top.RAMFF[2] ),
    .Y(_01109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18844_ (.A(\design_top.IOMUX[3][2] ),
    .Y(_10250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18845_ (.A(io_out[10]),
    .Y(_10251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18846_ (.A1(_10250_),
    .A2(_10242_),
    .B1(_10251_),
    .B2(_10244_),
    .X(_01110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18847_ (.A(\design_top.RAMFF[18] ),
    .Y(_01112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18848_ (.A(\design_top.IOMUX[3][18] ),
    .Y(_10252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18849_ (.A(\design_top.GPIOFF[2] ),
    .Y(_10253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18850_ (.A1(_10252_),
    .A2(_10242_),
    .B1(_10253_),
    .B2(_10244_),
    .X(_01113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18851_ (.A(\design_top.RAMFF[26] ),
    .Y(_01118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18852_ (.A(\design_top.IOMUX[3][26] ),
    .Y(_10254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18853_ (.A(\design_top.GPIOFF[10] ),
    .Y(_10255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18854_ (.A1(_10254_),
    .A2(_10242_),
    .B1(_10255_),
    .B2(_10244_),
    .X(_01119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18855_ (.A(\design_top.RAMFF[10] ),
    .Y(_01121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18856_ (.A(\design_top.IOMUX[3][10] ),
    .Y(_10256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18857_ (.A(\design_top.LEDFF[10] ),
    .Y(_10257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _18858_ (.A1(\design_top.uart0.UART_RFIFO[2] ),
    .A2(_10106_),
    .B1(_00833_),
    .Y(_10258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _18859_ (.A1(_10256_),
    .A2(_10236_),
    .B1(_10257_),
    .B2(_10238_),
    .C1(_10258_),
    .X(_01122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _18860_ (.A1(_10706_),
    .A2(\design_top.core0.PC[2] ),
    .B1(_10171_),
    .Y(_10259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18861_ (.A1_N(_10175_),
    .A2_N(_10259_),
    .B1(_10175_),
    .B2(_10259_),
    .X(_01130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18862_ (.A(\design_top.core0.REG1[6][31] ),
    .Y(_02671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18863_ (.A(\design_top.core0.NXPC[3] ),
    .Y(_01132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18864_ (.A1_N(_03163_),
    .A2_N(_09964_),
    .B1(_03163_),
    .B2(_09964_),
    .X(_01133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18865_ (.A1_N(_10046_),
    .A2_N(_10050_),
    .B1(_10046_),
    .B2(_10050_),
    .X(_01134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18866_ (.A(\design_top.core0.REG1[4][31] ),
    .Y(_02669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18867_ (.A(_10084_),
    .B(_00816_),
    .X(_01135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18868_ (.A(_10086_),
    .B(_01135_),
    .X(_01136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18869_ (.A(_10087_),
    .X(_10260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18870_ (.A(_10260_),
    .X(_10261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18871_ (.A(_10261_),
    .B(_01136_),
    .X(_01137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18872_ (.A(\design_top.core0.REG1[5][31] ),
    .Y(_02670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _18873_ (.A(_01154_),
    .B(_00827_),
    .C(_00828_),
    .X(_01155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18874_ (.A(\design_top.RAMFF[3] ),
    .Y(_01158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18875_ (.A(\design_top.IOMUX[3][3] ),
    .Y(_10262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18876_ (.A(_10096_),
    .X(_10263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18877_ (.A(io_out[11]),
    .Y(_10264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18878_ (.A(_10100_),
    .X(_10265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18879_ (.A1(_10262_),
    .A2(_10263_),
    .B1(_10264_),
    .B2(_10265_),
    .X(_01159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18880_ (.A(\design_top.RAMFF[19] ),
    .Y(_01161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18881_ (.A(\design_top.IOMUX[3][19] ),
    .Y(_10266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18882_ (.A(\design_top.GPIOFF[3] ),
    .Y(_10267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18883_ (.A1(_10266_),
    .A2(_10263_),
    .B1(_10267_),
    .B2(_10265_),
    .X(_01162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18884_ (.A(\design_top.RAMFF[27] ),
    .Y(_01166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18885_ (.A(\design_top.IOMUX[3][27] ),
    .Y(_10268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18886_ (.A(\design_top.GPIOFF[11] ),
    .Y(_10269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18887_ (.A1(_10268_),
    .A2(_10263_),
    .B1(_10269_),
    .B2(_10265_),
    .X(_01167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18888_ (.A(\design_top.RAMFF[11] ),
    .Y(_01169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18889_ (.A(\design_top.IOMUX[3][11] ),
    .Y(_10270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18890_ (.A(\design_top.LEDFF[11] ),
    .Y(_10271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _18891_ (.A(\design_top.uart0.UART_RFIFO[3] ),
    .B(_10107_),
    .Y(_10272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _18892_ (.A1(_10270_),
    .A2(_10236_),
    .B1(_10271_),
    .B2(_10238_),
    .C1(_10272_),
    .X(_01170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18893_ (.A(\design_top.core0.REG1[2][31] ),
    .Y(_02666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _18894_ (.A1(_10702_),
    .A2(\design_top.core0.PC[3] ),
    .B1(_10170_),
    .X(_10273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18895_ (.A1_N(_10177_),
    .A2_N(_10273_),
    .B1(_10177_),
    .B2(_10273_),
    .X(_01834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18896_ (.A(_01834_),
    .Y(_01178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18897_ (.A(\design_top.core0.REG1[3][31] ),
    .Y(_02667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18898_ (.A(\design_top.core0.NXPC[4] ),
    .Y(_01180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18899_ (.A1_N(_03164_),
    .A2_N(_09965_),
    .B1(_03164_),
    .B2(_09965_),
    .X(_01182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18900_ (.A1_N(_08583_),
    .A2_N(_10051_),
    .B1(_08583_),
    .B2(_10051_),
    .X(_01183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18901_ (.A(\design_top.core0.REG1[1][31] ),
    .Y(_02665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18902_ (.A(_10045_),
    .X(_10274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18903_ (.A(_10274_),
    .B(_01186_),
    .X(_01187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18904_ (.A(_10261_),
    .B(_01187_),
    .X(_01188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18905_ (.A(_10084_),
    .B(_00973_),
    .X(_01193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18906_ (.A(_10090_),
    .X(_10275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18907_ (.A(_10092_),
    .X(_10276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _18908_ (.A(_01198_),
    .B(_10275_),
    .C(_10276_),
    .X(_01199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18909_ (.A(\design_top.RAMFF[4] ),
    .Y(_01202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18910_ (.A(\design_top.IOMUX[3][4] ),
    .Y(_10277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18911_ (.A(\design_top.LEDFF[4] ),
    .Y(_10278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18912_ (.A1(_10277_),
    .A2(_10263_),
    .B1(_10278_),
    .B2(_10265_),
    .X(_01203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18913_ (.A(\design_top.RAMFF[20] ),
    .Y(_01205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18914_ (.A(\design_top.IOMUX[3][20] ),
    .Y(_10279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18915_ (.A(\design_top.GPIOFF[4] ),
    .Y(_10280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18916_ (.A1(_10279_),
    .A2(_10263_),
    .B1(_10280_),
    .B2(_10265_),
    .X(_01206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18917_ (.A(\design_top.RAMFF[28] ),
    .Y(_01210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18918_ (.A(\design_top.IOMUX[3][28] ),
    .Y(_10281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18919_ (.A(_10095_),
    .X(_10282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18920_ (.A(\design_top.GPIOFF[12] ),
    .Y(_10283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18921_ (.A(_10099_),
    .X(_10284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18922_ (.A1(_10281_),
    .A2(_10282_),
    .B1(_10283_),
    .B2(_10284_),
    .X(_01211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18923_ (.A(\design_top.RAMFF[12] ),
    .Y(_01213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18924_ (.A(\design_top.IOMUX[3][12] ),
    .Y(_10285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18925_ (.A(\design_top.LEDFF[12] ),
    .Y(_10286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _18926_ (.A(\design_top.uart0.UART_RFIFO[4] ),
    .B(_10107_),
    .Y(_10287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _18927_ (.A1(_10285_),
    .A2(_10236_),
    .B1(_10286_),
    .B2(_10238_),
    .C1(_10287_),
    .X(_01214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18928_ (.A1_N(_10178_),
    .A2_N(_10169_),
    .B1(_10178_),
    .B2(_10169_),
    .X(_01838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18929_ (.A(_01838_),
    .Y(_01222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18930_ (.A(\design_top.core0.NXPC[5] ),
    .Y(_01224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _18931_ (.A(_08581_),
    .X(_10288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _18932_ (.A1(_03164_),
    .A2(_09965_),
    .B1(_01181_),
    .Y(_10289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18933_ (.A1_N(_10288_),
    .A2_N(_10289_),
    .B1(_10288_),
    .B2(_10289_),
    .X(_01225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18934_ (.A1(_03103_),
    .A2(_03097_),
    .B1(_08583_),
    .B2(_10051_),
    .X(_10290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18935_ (.A1_N(_10288_),
    .A2_N(_10290_),
    .B1(_10288_),
    .B2(_10290_),
    .X(_01226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18936_ (.A(_10274_),
    .B(_01228_),
    .X(_01229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18937_ (.A(_10261_),
    .B(_01229_),
    .X(_01230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18938_ (.A(_10084_),
    .B(_01043_),
    .X(_01235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _18939_ (.A(_01240_),
    .B(_10275_),
    .C(_10276_),
    .X(_01241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18940_ (.A(\design_top.RAMFF[5] ),
    .Y(_01244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18941_ (.A(\design_top.IOMUX[3][5] ),
    .Y(_10291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18942_ (.A(\design_top.LEDFF[5] ),
    .Y(_10292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18943_ (.A1(_10291_),
    .A2(_10282_),
    .B1(_10292_),
    .B2(_10284_),
    .X(_01245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18944_ (.A(\design_top.RAMFF[21] ),
    .Y(_01247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18945_ (.A(\design_top.IOMUX[3][21] ),
    .Y(_10293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18946_ (.A(\design_top.GPIOFF[5] ),
    .Y(_10294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18947_ (.A1(_10293_),
    .A2(_10282_),
    .B1(_10294_),
    .B2(_10284_),
    .X(_01248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18948_ (.A(\design_top.RAMFF[29] ),
    .Y(_01253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18949_ (.A(\design_top.IOMUX[3][29] ),
    .Y(_10295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18950_ (.A(\design_top.GPIOFF[13] ),
    .Y(_10296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18951_ (.A1(_10295_),
    .A2(_10282_),
    .B1(_10296_),
    .B2(_10284_),
    .X(_01254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18952_ (.A(\design_top.RAMFF[13] ),
    .Y(_01256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18953_ (.A(\design_top.IOMUX[3][13] ),
    .Y(_10297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18954_ (.A(\design_top.LEDFF[13] ),
    .Y(_10298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _18955_ (.A1(\design_top.uart0.UART_RFIFO[5] ),
    .A2(_10106_),
    .B1(_00833_),
    .Y(_10299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _18956_ (.A1(_10297_),
    .A2(_10096_),
    .B1(_10298_),
    .B2(_10100_),
    .C1(_10299_),
    .X(_01257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18957_ (.A1(_08447_),
    .A2(\design_top.core0.PC[4] ),
    .B1(_10178_),
    .B2(_10169_),
    .X(_10300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18958_ (.A1_N(_10168_),
    .A2_N(_10300_),
    .B1(_10168_),
    .B2(_10300_),
    .X(_01841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18959_ (.A(_01841_),
    .Y(_01265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18960_ (.A(\design_top.core0.NXPC[6] ),
    .Y(_01267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _18961_ (.A(_09966_),
    .B(_09967_),
    .X(_10301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18962_ (.A1_N(_01269_),
    .A2_N(_10301_),
    .B1(_01269_),
    .B2(_10301_),
    .X(_01270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18963_ (.A1(_00811_),
    .A2(_03094_),
    .B1(_10288_),
    .B2(_10290_),
    .X(_10302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18964_ (.A1_N(_08580_),
    .A2_N(_10302_),
    .B1(_08580_),
    .B2(_10302_),
    .X(_01271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18965_ (.A(_10274_),
    .B(_01274_),
    .X(_01275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18966_ (.A(_10261_),
    .B(_01275_),
    .X(_01276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18967_ (.A(_10084_),
    .B(_01098_),
    .X(_01281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _18968_ (.A(_01286_),
    .B(_10275_),
    .C(_10276_),
    .X(_01287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18969_ (.A(\design_top.RAMFF[6] ),
    .Y(_01290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18970_ (.A(\design_top.IOMUX[3][6] ),
    .Y(_10303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18971_ (.A(\design_top.LEDFF[6] ),
    .Y(_10304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18972_ (.A1(_10303_),
    .A2(_10282_),
    .B1(_10304_),
    .B2(_10284_),
    .X(_01291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18973_ (.A(\design_top.RAMFF[22] ),
    .Y(_01293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18974_ (.A(\design_top.IOMUX[3][22] ),
    .Y(_10305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18975_ (.A(\design_top.GPIOFF[6] ),
    .Y(_10306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18976_ (.A1(_10305_),
    .A2(_10103_),
    .B1(_10306_),
    .B2(_10105_),
    .X(_01294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18977_ (.A(\design_top.RAMFF[30] ),
    .Y(_01299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18978_ (.A(\design_top.IOMUX[3][30] ),
    .Y(_10307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18979_ (.A(\design_top.GPIOFF[14] ),
    .Y(_10308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18980_ (.A1(_10307_),
    .A2(_10103_),
    .B1(_10308_),
    .B2(_10105_),
    .X(_01300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18981_ (.A(\design_top.RAMFF[14] ),
    .Y(_01302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18982_ (.A(\design_top.IOMUX[3][14] ),
    .Y(_10309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18983_ (.A(\design_top.LEDFF[14] ),
    .Y(_10310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _18984_ (.A1(\design_top.uart0.UART_RFIFO[6] ),
    .A2(_10106_),
    .B1(_00833_),
    .Y(_10311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _18985_ (.A1(_10309_),
    .A2(_10096_),
    .B1(_10310_),
    .B2(_10100_),
    .C1(_10311_),
    .X(_01303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18986_ (.A1_N(_10181_),
    .A2_N(_10167_),
    .B1(_10181_),
    .B2(_10167_),
    .X(_01844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18987_ (.A(_01844_),
    .Y(_01311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18988_ (.A(\design_top.core0.NXPC[7] ),
    .Y(_01313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _18989_ (.A1(_01269_),
    .A2(_10301_),
    .B1(_01268_),
    .Y(_10312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _18990_ (.A1_N(_09952_),
    .A2_N(_10312_),
    .B1(_09952_),
    .B2(_10312_),
    .X(_01314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18991_ (.A1(_03087_),
    .A2(_03081_),
    .B1(_08580_),
    .B2(_10302_),
    .X(_10313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18992_ (.A(_10313_),
    .Y(_10314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _18993_ (.A1(_03166_),
    .A2(_10313_),
    .B1(_09952_),
    .B2(_10314_),
    .X(_01315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18994_ (.A(_10274_),
    .B(_00817_),
    .X(_01316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _18995_ (.A(_10261_),
    .B(_01316_),
    .X(_01317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _18996_ (.A(_01325_),
    .B(_10275_),
    .C(_10276_),
    .X(_01326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _18997_ (.A1(_08444_),
    .A2(\design_top.core0.PC[6] ),
    .B1(_10181_),
    .B2(_10167_),
    .X(_10315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _18998_ (.A1_N(_10166_),
    .A2_N(_10315_),
    .B1(_10166_),
    .B2(_10315_),
    .X(_01848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _18999_ (.A(_01848_),
    .Y(_01334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19000_ (.A(\design_top.core0.NXPC[8] ),
    .Y(_01336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19001_ (.A(_08592_),
    .X(_10316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19002_ (.A(_09969_),
    .Y(_10317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _19003_ (.A1(_10316_),
    .A2(_10317_),
    .B1(_03167_),
    .B2(_09969_),
    .X(_01338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19004_ (.A1_N(_10316_),
    .A2_N(_10055_),
    .B1(_10316_),
    .B2(_10055_),
    .X(_01339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19005_ (.A(_10260_),
    .X(_10318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19006_ (.A(_10318_),
    .B(_01343_),
    .X(_01344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19007_ (.A(_10274_),
    .B(_00974_),
    .X(_01346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19008_ (.A(_01349_),
    .B(_10275_),
    .C(_10276_),
    .X(_01350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19009_ (.A(_10184_),
    .X(_10319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _19010_ (.A1_N(_10319_),
    .A2_N(_10154_),
    .B1(_10319_),
    .B2(_10154_),
    .X(_01851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19011_ (.A(_01851_),
    .Y(_01358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19012_ (.A(\design_top.core0.NXPC[9] ),
    .Y(_01360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19013_ (.A(_08591_),
    .X(_10320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _19014_ (.A1(_03167_),
    .A2(_09969_),
    .B1(_01337_),
    .Y(_10321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19015_ (.A1_N(_10320_),
    .A2_N(_10321_),
    .B1(_10320_),
    .B2(_10321_),
    .X(_01361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19016_ (.A1(_03071_),
    .A2(_03065_),
    .B1(_10316_),
    .B2(_10055_),
    .X(_10322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19017_ (.A1_N(_10320_),
    .A2_N(_10322_),
    .B1(_10320_),
    .B2(_10322_),
    .X(_01362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19018_ (.A(_10318_),
    .B(_01365_),
    .X(_01366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19019_ (.A(_10045_),
    .X(_10323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19020_ (.A(_10323_),
    .B(_01044_),
    .X(_01368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19021_ (.A(_10090_),
    .X(_10324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19022_ (.A(_10092_),
    .X(_10325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19023_ (.A(_01371_),
    .B(_10324_),
    .C(_10325_),
    .X(_01372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _19024_ (.A1(_08441_),
    .A2(\design_top.core0.PC[8] ),
    .B1(_10319_),
    .B2(_10154_),
    .X(_10326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _19025_ (.A1_N(_10153_),
    .A2_N(_10326_),
    .B1(_10153_),
    .B2(_10326_),
    .X(_01855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19026_ (.A(_01855_),
    .Y(_01380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19027_ (.A(\design_top.core0.NXPC[10] ),
    .Y(_01382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31oi_2 _19028_ (.A1(_10320_),
    .A2(_10316_),
    .A3(_10317_),
    .B1(_09970_),
    .Y(_10327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19029_ (.A1_N(_03169_),
    .A2_N(_10327_),
    .B1(_03169_),
    .B2(_10327_),
    .X(_01384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19030_ (.A1(_00805_),
    .A2(_03062_),
    .B1(_08591_),
    .B2(_10322_),
    .X(_10328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19031_ (.A1_N(_08595_),
    .A2_N(_10328_),
    .B1(_08595_),
    .B2(_10328_),
    .X(_01385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19032_ (.A(_10318_),
    .B(_01389_),
    .X(_01390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19033_ (.A(_10323_),
    .B(_01099_),
    .X(_01392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19034_ (.A(_01395_),
    .B(_10324_),
    .C(_10325_),
    .X(_01396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19035_ (.A(_10152_),
    .Y(_10329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31oi_2 _19036_ (.A1(_10153_),
    .A2(_10154_),
    .A3(_10319_),
    .B1(_10186_),
    .Y(_10330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19037_ (.A1_N(_10329_),
    .A2_N(_10330_),
    .B1(_10329_),
    .B2(_10330_),
    .X(_01404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19038_ (.A(\design_top.core0.NXPC[11] ),
    .Y(_01406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _19039_ (.A1(_03169_),
    .A2(_10327_),
    .B1(_01383_),
    .Y(_10331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19040_ (.A1_N(_08589_),
    .A2_N(_10331_),
    .B1(_08589_),
    .B2(_10331_),
    .X(_01407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19041_ (.A1(_03055_),
    .A2(_03049_),
    .B1(_08595_),
    .B2(_10328_),
    .X(_10332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19042_ (.A(_10332_),
    .Y(_10333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19043_ (.A1(_03170_),
    .A2(_10332_),
    .B1(_08589_),
    .B2(_10333_),
    .X(_01408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19044_ (.A(_10318_),
    .B(_01410_),
    .X(_01411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19045_ (.A(_10323_),
    .B(_01149_),
    .X(_01413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19046_ (.A(_01416_),
    .B(_10324_),
    .C(_10325_),
    .X(_01417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19047_ (.A1(_02810_),
    .A2(_10151_),
    .B1(_10329_),
    .B2(_10330_),
    .X(_10334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19048_ (.A1_N(_10149_),
    .A2_N(_10334_),
    .B1(_10149_),
    .B2(_10334_),
    .X(_01425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19049_ (.A(\design_top.core0.NXPC[12] ),
    .Y(_01427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _19050_ (.A1(_09969_),
    .A2(_09958_),
    .B1(_09972_),
    .Y(_10335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19051_ (.A(_10335_),
    .Y(_10336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _19052_ (.A1(_08573_),
    .A2(_10335_),
    .B1(_03171_),
    .B2(_10336_),
    .X(_01429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19053_ (.A(_10059_),
    .X(_10337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19054_ (.A1_N(_10337_),
    .A2_N(_10044_),
    .B1(_10337_),
    .B2(_10044_),
    .X(_01430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19055_ (.A(_10318_),
    .B(_01434_),
    .X(_01435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19056_ (.A(_10323_),
    .B(_01193_),
    .X(_01437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19057_ (.A(_01440_),
    .B(_10324_),
    .C(_10325_),
    .X(_01441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _19058_ (.A1(_10319_),
    .A2(_10155_),
    .B1(_10188_),
    .Y(_10338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19059_ (.A(_10338_),
    .Y(_10339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19060_ (.A1(_10160_),
    .A2(_10338_),
    .B1(_10159_),
    .B2(_10339_),
    .X(_01867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19061_ (.A(_01867_),
    .Y(_01449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19062_ (.A(\design_top.core0.NXPC[13] ),
    .Y(_01451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _19063_ (.A1(_03171_),
    .A2(_10336_),
    .B1(_01428_),
    .Y(_10340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19064_ (.A1_N(_08568_),
    .A2_N(_10340_),
    .B1(_08568_),
    .B2(_10340_),
    .X(_01452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19065_ (.A(_10043_),
    .X(_03033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19066_ (.A1(_03157_),
    .A2(_03033_),
    .B1(_10337_),
    .B2(_10044_),
    .X(_10341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19067_ (.A1_N(_10042_),
    .A2_N(_10341_),
    .B1(_10042_),
    .B2(_10341_),
    .X(_01453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19068_ (.A(_10087_),
    .X(_10342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19069_ (.A(_10342_),
    .B(_01456_),
    .X(_01457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19070_ (.A(_10323_),
    .B(_01235_),
    .X(_01459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19071_ (.A(_01462_),
    .B(_10324_),
    .C(_10325_),
    .X(_01463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19072_ (.A1(_02798_),
    .A2(_10158_),
    .B1(_10160_),
    .B2(_10338_),
    .X(_10343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19073_ (.A1_N(_10157_),
    .A2_N(_10343_),
    .B1(_10157_),
    .B2(_10343_),
    .X(_01471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19074_ (.A(_01472_),
    .B(_08787_),
    .Y(_01473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _19075_ (.A(\design_top.core0.RESMODE[0] ),
    .B(_10224_),
    .C(_03196_),
    .Y(_01474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19076_ (.A(\design_top.core0.NXPC[14] ),
    .Y(_01475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _19077_ (.A1(_03172_),
    .A2(_03171_),
    .A3(_10336_),
    .B1(_09973_),
    .X(_10344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19078_ (.A1_N(_01477_),
    .A2_N(_10344_),
    .B1(_01477_),
    .B2(_10344_),
    .X(_01478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _19079_ (.A1(_10042_),
    .A2(_10044_),
    .A3(_10337_),
    .B1(_10040_),
    .X(_10345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19080_ (.A1_N(_10035_),
    .A2_N(_10345_),
    .B1(_10035_),
    .B2(_10345_),
    .X(_01479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19081_ (.A(\design_top.DACK[0] ),
    .B(\design_top.DACK[1] ),
    .Y(_02858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19082_ (.A(_10342_),
    .B(_01483_),
    .X(_01484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19083_ (.A(_10045_),
    .B(_01281_),
    .X(_01486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19084_ (.A(_10089_),
    .X(_10346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19085_ (.A(_10091_),
    .X(_10347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19086_ (.A(_01489_),
    .B(_10346_),
    .C(_10347_),
    .X(_01490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31oi_2 _19087_ (.A1(_10156_),
    .A2(_10159_),
    .A3(_10339_),
    .B1(_10190_),
    .Y(_10348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19088_ (.A1_N(_10162_),
    .A2_N(_10348_),
    .B1(_10162_),
    .B2(_10348_),
    .X(_01498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19089_ (.A(\design_top.core0.NXPC[15] ),
    .Y(_01500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _19090_ (.A1(_01477_),
    .A2(_10344_),
    .B1(_01476_),
    .Y(_10349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19091_ (.A1_N(_08571_),
    .A2_N(_10349_),
    .B1(_08571_),
    .B2(_10349_),
    .X(_01501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19092_ (.A(_10734_),
    .X(_03016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19093_ (.A1(_03155_),
    .A2(_03016_),
    .B1(_10035_),
    .B2(_10345_),
    .X(_10350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19094_ (.A1_N(_10036_),
    .A2_N(_10350_),
    .B1(_10036_),
    .B2(_10350_),
    .X(_01502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19095_ (.A(_10342_),
    .B(_00818_),
    .X(_01503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19096_ (.A(_01506_),
    .B(_10346_),
    .C(_10347_),
    .X(_01507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19097_ (.A1(_02786_),
    .A2(_10161_),
    .B1(_10162_),
    .B2(_10348_),
    .X(_10351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19098_ (.A1_N(_10164_),
    .A2_N(_10351_),
    .B1(_10164_),
    .B2(_10351_),
    .X(_01514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19099_ (.A(\design_top.core0.NXPC[16] ),
    .Y(_01516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19100_ (.A(_09976_),
    .Y(_10352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _19101_ (.A1(_08547_),
    .A2(_10352_),
    .B1(_03174_),
    .B2(_09976_),
    .X(_01518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19102_ (.A1_N(_10061_),
    .A2_N(_10062_),
    .B1(_10061_),
    .B2(_10062_),
    .X(_01519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19103_ (.A(_10342_),
    .B(_00975_),
    .X(_01525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19104_ (.A(_01528_),
    .B(_10346_),
    .C(_10347_),
    .X(_01529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19105_ (.A(_10195_),
    .X(_10353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _19106_ (.A1_N(_10353_),
    .A2_N(_10136_),
    .B1(_10353_),
    .B2(_10136_),
    .X(_01883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19107_ (.A(_01883_),
    .Y(_01536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19108_ (.A(\design_top.core0.NXPC[17] ),
    .Y(_01538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _19109_ (.A1(_03174_),
    .A2(_09976_),
    .B1(_01517_),
    .Y(_10354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19110_ (.A1_N(_08540_),
    .A2_N(_10354_),
    .B1(_08540_),
    .B2(_10354_),
    .X(_01539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19111_ (.A(_10740_),
    .X(_02999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19112_ (.A1(_03153_),
    .A2(_02999_),
    .B1(_10061_),
    .B2(_10062_),
    .X(_10355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19113_ (.A1_N(_10063_),
    .A2_N(_10355_),
    .B1(_10063_),
    .B2(_10355_),
    .X(_01540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19114_ (.A(_10342_),
    .B(_01045_),
    .X(_01545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19115_ (.A(_01548_),
    .B(_10346_),
    .C(_10347_),
    .X(_01549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _19116_ (.A1(_08467_),
    .A2(\design_top.core0.PC[16] ),
    .B1(_10353_),
    .B2(_10136_),
    .X(_10356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _19117_ (.A1_N(_10135_),
    .A2_N(_10356_),
    .B1(_10135_),
    .B2(_10356_),
    .X(_01887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19118_ (.A(_01887_),
    .Y(_01556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19119_ (.A(\design_top.core0.NXPC[18] ),
    .Y(_01558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31oi_2 _19120_ (.A1(_08540_),
    .A2(_08547_),
    .A3(_10352_),
    .B1(_09977_),
    .Y(_10357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19121_ (.A1_N(_01560_),
    .A2_N(_10357_),
    .B1(_01560_),
    .B2(_10357_),
    .X(_01561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _19122_ (.A1(_10062_),
    .A2(_10063_),
    .A3(_10061_),
    .B1(_10031_),
    .X(_10358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19123_ (.A1_N(_10023_),
    .A2_N(_10358_),
    .B1(_10023_),
    .B2(_10358_),
    .X(_01562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19124_ (.A(_10087_),
    .X(_10359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19125_ (.A(_10359_),
    .B(_01100_),
    .X(_01568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19126_ (.A(_01571_),
    .B(_10346_),
    .C(_10347_),
    .X(_01572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19127_ (.A(_10134_),
    .Y(_10360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31oi_2 _19128_ (.A1(_10135_),
    .A2(_10136_),
    .A3(_10353_),
    .B1(_10197_),
    .Y(_10361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19129_ (.A1_N(_10360_),
    .A2_N(_10361_),
    .B1(_10360_),
    .B2(_10361_),
    .X(_01579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19130_ (.A(\design_top.core0.NXPC[19] ),
    .Y(_01581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _19131_ (.A1(_01560_),
    .A2(_10357_),
    .B1(_01559_),
    .Y(_10362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19132_ (.A1_N(_08542_),
    .A2_N(_10362_),
    .B1(_08542_),
    .B2(_10362_),
    .X(_01582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19133_ (.A(_10021_),
    .X(_02982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19134_ (.A1(_03151_),
    .A2(_02982_),
    .B1(_10023_),
    .B2(_10358_),
    .X(_10363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19135_ (.A1_N(_10026_),
    .A2_N(_10363_),
    .B1(_10026_),
    .B2(_10363_),
    .X(_01583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19136_ (.A(_10359_),
    .B(_01150_),
    .X(_01587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19137_ (.A(_10089_),
    .X(_10364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19138_ (.A(_10091_),
    .X(_10365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19139_ (.A(_01590_),
    .B(_10364_),
    .C(_10365_),
    .X(_01591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19140_ (.A1(_02762_),
    .A2(_10133_),
    .B1(_10360_),
    .B2(_10361_),
    .X(_10366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19141_ (.A1_N(_10131_),
    .A2_N(_10366_),
    .B1(_10131_),
    .B2(_10366_),
    .X(_01598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19142_ (.A(\design_top.core0.NXPC[20] ),
    .Y(_01600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _19143_ (.A1(_09976_),
    .A2(_09956_),
    .B1(_09979_),
    .Y(_10367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19144_ (.A(_10367_),
    .Y(_10368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _19145_ (.A1(_08535_),
    .A2(_10367_),
    .B1(_03177_),
    .B2(_10368_),
    .X(_01602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19146_ (.A1_N(_10018_),
    .A2_N(_10066_),
    .B1(_10018_),
    .B2(_10066_),
    .X(_01603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19147_ (.A(_10359_),
    .B(_01194_),
    .X(_01609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19148_ (.A(_01612_),
    .B(_10364_),
    .C(_10365_),
    .X(_01613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _19149_ (.A1(_10353_),
    .A2(_10137_),
    .B1(_10199_),
    .Y(_10369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19150_ (.A(_10369_),
    .Y(_10370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19151_ (.A1(_10142_),
    .A2(_10369_),
    .B1(_10141_),
    .B2(_10370_),
    .X(_01899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19152_ (.A(_01899_),
    .Y(_01620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19153_ (.A(\design_top.core0.NXPC[21] ),
    .Y(_01622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _19154_ (.A1(_03177_),
    .A2(_10368_),
    .B1(_01601_),
    .Y(_10371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19155_ (.A1_N(_08532_),
    .A2_N(_10371_),
    .B1(_08532_),
    .B2(_10371_),
    .X(_01623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19156_ (.A(_10624_),
    .X(_02965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19157_ (.A1(_03149_),
    .A2(_02965_),
    .B1(_10018_),
    .B2(_10066_),
    .X(_10372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19158_ (.A1_N(_10019_),
    .A2_N(_10372_),
    .B1(_10019_),
    .B2(_10372_),
    .X(_01624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19159_ (.A(_10359_),
    .B(_01236_),
    .X(_01629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19160_ (.A(_01632_),
    .B(_10364_),
    .C(_10365_),
    .X(_01633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19161_ (.A1(_02750_),
    .A2(_10140_),
    .B1(_10142_),
    .B2(_10369_),
    .X(_10373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19162_ (.A1_N(_10139_),
    .A2_N(_10373_),
    .B1(_10139_),
    .B2(_10373_),
    .X(_01640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19163_ (.A(\design_top.core0.NXPC[22] ),
    .Y(_01642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _19164_ (.A1(_03178_),
    .A2(_03177_),
    .A3(_10368_),
    .B1(_09980_),
    .X(_10374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19165_ (.A1_N(_03179_),
    .A2_N(_10374_),
    .B1(_03179_),
    .B2(_10374_),
    .X(_01644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _19166_ (.A1(_10018_),
    .A2(_10019_),
    .A3(_10066_),
    .B1(_10017_),
    .X(_10375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19167_ (.A1_N(_10008_),
    .A2_N(_10375_),
    .B1(_10008_),
    .B2(_10375_),
    .X(_01645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19168_ (.A(_10359_),
    .B(_01282_),
    .X(_01651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19169_ (.A(_01654_),
    .B(_10364_),
    .C(_10365_),
    .X(_01655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31oi_2 _19170_ (.A1(_10138_),
    .A2(_10141_),
    .A3(_10370_),
    .B1(_10201_),
    .Y(_10376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19171_ (.A1_N(_10144_),
    .A2_N(_10376_),
    .B1(_10144_),
    .B2(_10376_),
    .X(_01662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19172_ (.A(\design_top.core0.NXPC[23] ),
    .Y(_01664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _19173_ (.A1(_03179_),
    .A2(_10374_),
    .B1(_01643_),
    .Y(_10377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19174_ (.A1_N(_08530_),
    .A2_N(_10377_),
    .B1(_08530_),
    .B2(_10377_),
    .X(_01665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19175_ (.A(_10006_),
    .X(_02948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19176_ (.A1(_03147_),
    .A2(_02948_),
    .B1(_10008_),
    .B2(_10375_),
    .X(_10378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19177_ (.A1_N(_10012_),
    .A2_N(_10378_),
    .B1(_10012_),
    .B2(_10378_),
    .X(_01666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19178_ (.A(_10087_),
    .X(_10379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19179_ (.A(_10379_),
    .B(_01322_),
    .X(_01669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19180_ (.A(_01672_),
    .B(_10364_),
    .C(_10365_),
    .X(_01673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19181_ (.A1(_02738_),
    .A2(_10143_),
    .B1(_10144_),
    .B2(_10376_),
    .X(_10380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19182_ (.A1_N(_10146_),
    .A2_N(_10380_),
    .B1(_10146_),
    .B2(_10380_),
    .X(_01680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19183_ (.A(\design_top.core0.NXPC[24] ),
    .Y(_01682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19184_ (.A1_N(_03181_),
    .A2_N(_09983_),
    .B1(_03181_),
    .B2(_09983_),
    .X(_01684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19185_ (.A1_N(_10068_),
    .A2_N(_10069_),
    .B1(_10068_),
    .B2(_10069_),
    .X(_01685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19186_ (.A(_10379_),
    .B(_01346_),
    .X(_01691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19187_ (.A(_10089_),
    .X(_10381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19188_ (.A(_10091_),
    .X(_10382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19189_ (.A(_01694_),
    .B(_10381_),
    .C(_10382_),
    .X(_01695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19190_ (.A1(_10207_),
    .A2(_10129_),
    .B1(_10206_),
    .B2(_10128_),
    .X(_01915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19191_ (.A(_01915_),
    .Y(_01702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19192_ (.A(\design_top.core0.NXPC[25] ),
    .Y(_01704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _19193_ (.A1(_03181_),
    .A2(_09983_),
    .B1(_01683_),
    .Y(_10383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19194_ (.A1_N(_08552_),
    .A2_N(_10383_),
    .B1(_08552_),
    .B2(_10383_),
    .X(_01705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19195_ (.A(_10613_),
    .X(_02931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19196_ (.A1(_03145_),
    .A2(_02931_),
    .B1(_10068_),
    .B2(_10069_),
    .X(_10384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19197_ (.A1_N(_10070_),
    .A2_N(_10384_),
    .B1(_10070_),
    .B2(_10384_),
    .X(_01706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19198_ (.A(_09939_),
    .B(_02849_),
    .Y(_02863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19199_ (.A(_10379_),
    .B(_01368_),
    .X(_01711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19200_ (.A(_01714_),
    .B(_10381_),
    .C(_10382_),
    .X(_01715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _19201_ (.A1(_08460_),
    .A2(\design_top.core0.PC[24] ),
    .B1(_10206_),
    .B2(_10128_),
    .X(_10385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _19202_ (.A1_N(_10126_),
    .A2_N(_10385_),
    .B1(_10126_),
    .B2(_10385_),
    .X(_01919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19203_ (.A(_01919_),
    .Y(_01722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19204_ (.A(\design_top.core0.NXPC[26] ),
    .Y(_01724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _19205_ (.A1(_03182_),
    .A2(_03181_),
    .A3(_09983_),
    .B1(_09985_),
    .X(_10386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19206_ (.A1_N(_03183_),
    .A2_N(_10386_),
    .B1(_03183_),
    .B2(_10386_),
    .X(_01726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _19207_ (.A1(_10069_),
    .A2(_10070_),
    .A3(_10068_),
    .B1(_10005_),
    .X(_10387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19208_ (.A1_N(_09997_),
    .A2_N(_10387_),
    .B1(_09997_),
    .B2(_10387_),
    .X(_01727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19209_ (.A(_10379_),
    .B(_01392_),
    .X(_01733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19210_ (.A(_01736_),
    .B(_10381_),
    .C(_10382_),
    .X(_01737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _19211_ (.A1(_10127_),
    .A2(_10129_),
    .A3(_10207_),
    .B1(_10124_),
    .X(_10388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19212_ (.A1_N(_10121_),
    .A2_N(_10388_),
    .B1(_10121_),
    .B2(_10388_),
    .X(_01744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19213_ (.A(\design_top.core0.NXPC[27] ),
    .Y(_01746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _19214_ (.A1(_03183_),
    .A2(_10386_),
    .B1(_01725_),
    .Y(_10389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19215_ (.A1_N(_08550_),
    .A2_N(_10389_),
    .B1(_08550_),
    .B2(_10389_),
    .X(_01747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19216_ (.A1(_03143_),
    .A2(_02914_),
    .B1(_09997_),
    .B2(_10387_),
    .X(_10390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19217_ (.A1_N(_10000_),
    .A2_N(_10390_),
    .B1(_10000_),
    .B2(_10390_),
    .X(_01748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19218_ (.A(_10379_),
    .B(_01413_),
    .X(_01752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19219_ (.A(_01755_),
    .B(_10381_),
    .C(_10382_),
    .X(_01756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19220_ (.A1(_02714_),
    .A2(_10118_),
    .B1(_10121_),
    .B2(_10388_),
    .X(_10391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19221_ (.A1_N(_10120_),
    .A2_N(_10391_),
    .B1(_10120_),
    .B2(_10391_),
    .X(_01763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19222_ (.A(\design_top.core0.NXPC[28] ),
    .Y(_01765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19223_ (.A1_N(_03185_),
    .A2_N(_09987_),
    .B1(_03185_),
    .B2(_09987_),
    .X(_01767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19224_ (.A1_N(_10073_),
    .A2_N(_09993_),
    .B1(_10073_),
    .B2(_09993_),
    .X(_01768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19225_ (.A(_10260_),
    .B(_01437_),
    .X(_01774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19226_ (.A(_01777_),
    .B(_10381_),
    .C(_10382_),
    .X(_01778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _19227_ (.A1(_10605_),
    .A2(\design_top.core0.PC[28] ),
    .B1(_10116_),
    .X(_10392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _19228_ (.A1_N(_10209_),
    .A2_N(_10392_),
    .B1(_10209_),
    .B2(_10392_),
    .X(_01931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19229_ (.A(_01931_),
    .Y(_01785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19230_ (.A(\design_top.core0.NXPC[29] ),
    .Y(_01787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _19231_ (.A(_01766_),
    .B(_09988_),
    .Y(_10393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a32o_2 _19232_ (.A1(_01766_),
    .A2(_09988_),
    .A3(_03186_),
    .B1(_08560_),
    .B2(_10393_),
    .X(_01788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19233_ (.A1(_03141_),
    .A2(_02897_),
    .B1(_10073_),
    .B2(_09993_),
    .X(_10394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19234_ (.A1_N(_09995_),
    .A2_N(_10394_),
    .B1(_09995_),
    .B2(_10394_),
    .X(_01789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19235_ (.A(_10260_),
    .B(_01459_),
    .X(_01794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19236_ (.A(_01797_),
    .B(_10090_),
    .C(_10092_),
    .X(_01798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _19237_ (.A1(_10600_),
    .A2(\design_top.core0.PC[29] ),
    .B1(_10115_),
    .X(_10395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _19238_ (.A1_N(_10210_),
    .A2_N(_10395_),
    .B1(_10210_),
    .B2(_10395_),
    .X(_01935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19239_ (.A(_01935_),
    .Y(_01805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19240_ (.A(\design_top.core0.NXPC[30] ),
    .Y(_01807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19241_ (.A1_N(_03187_),
    .A2_N(_09989_),
    .B1(_03187_),
    .B2(_09989_),
    .X(_01808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19242_ (.A1_N(_09991_),
    .A2_N(_10076_),
    .B1(_09991_),
    .B2(_10076_),
    .X(_01809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19243_ (.A(_10260_),
    .B(_01486_),
    .X(_01815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19244_ (.A(_01818_),
    .B(_10090_),
    .C(_10092_),
    .X(_01819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19245_ (.A1_N(_10114_),
    .A2_N(_10211_),
    .B1(_10114_),
    .B2(_10211_),
    .X(_01826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19246_ (.A(io_out[18]),
    .Y(_01830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19247_ (.A(_01130_),
    .Y(_01831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _19248_ (.A(io_out[19]),
    .B(io_out[18]),
    .Y(_10396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19249_ (.A1(io_out[19]),
    .A2(io_out[18]),
    .B1(_10396_),
    .X(_01833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19250_ (.A(_10396_),
    .Y(_10397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _19251_ (.A1_N(_08525_),
    .A2_N(_10397_),
    .B1(_08525_),
    .B2(_10397_),
    .X(_01836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _19252_ (.A(\design_top.IADDR[4] ),
    .B(_10397_),
    .C(\design_top.IADDR[5] ),
    .X(_10398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _19253_ (.A1(_08525_),
    .A2(_10397_),
    .B1(\design_top.IADDR[5] ),
    .Y(_10399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19254_ (.A(_10398_),
    .B(_10399_),
    .Y(_01840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _19255_ (.A(\design_top.IADDR[6] ),
    .B(_10398_),
    .Y(_10400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19256_ (.A1(\design_top.IADDR[6] ),
    .A2(_10398_),
    .B1(_10400_),
    .X(_01843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19257_ (.A(_10400_),
    .Y(_10401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _19258_ (.A(\design_top.IADDR[7] ),
    .B(_10401_),
    .Y(_10402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19259_ (.A1(\design_top.IADDR[7] ),
    .A2(_10401_),
    .B1(_10402_),
    .X(_01846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19260_ (.A(_10402_),
    .Y(_10403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _19261_ (.A(\design_top.IADDR[8] ),
    .B(_10403_),
    .Y(_10404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19262_ (.A1(\design_top.IADDR[8] ),
    .A2(_10403_),
    .B1(_10404_),
    .X(_01850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19263_ (.A(_10724_),
    .X(_10405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19264_ (.A(_10405_),
    .Y(_10406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19265_ (.A1(_10405_),
    .A2(_10729_),
    .B1(_10406_),
    .B2(_10728_),
    .X(_01852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19266_ (.A(_10404_),
    .Y(_10407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _19267_ (.A(\design_top.IADDR[9] ),
    .B(_10407_),
    .Y(_10408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19268_ (.A1(\design_top.IADDR[9] ),
    .A2(_10407_),
    .B1(_10408_),
    .X(_01854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19269_ (.A1(_02822_),
    .A2(_03065_),
    .B1(_10405_),
    .B2(_10729_),
    .X(_10409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19270_ (.A(_10409_),
    .Y(_10410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19271_ (.A1(_10726_),
    .A2(_10409_),
    .B1(_10725_),
    .B2(_10410_),
    .X(_01856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19272_ (.A(\design_top.IADDR[10] ),
    .Y(_10411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19273_ (.A(_10411_),
    .B(_10408_),
    .Y(_10412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _19274_ (.A1(_10411_),
    .A2(_10408_),
    .B1(_10412_),
    .Y(_01858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19275_ (.A(_01404_),
    .Y(_01859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _19276_ (.A1(_10726_),
    .A2(_10729_),
    .A3(_10405_),
    .B1(_10687_),
    .X(_10413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19277_ (.A(_10413_),
    .Y(_10414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19278_ (.A1(_10684_),
    .A2(_10413_),
    .B1(_10683_),
    .B2(_10414_),
    .X(_01860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _19279_ (.A(_10408_),
    .B(_10411_),
    .C_N(\design_top.IADDR[11] ),
    .X(_10415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19280_ (.A1(\design_top.IADDR[11] ),
    .A2(_10412_),
    .B1(_10415_),
    .X(_01862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19281_ (.A(_01425_),
    .Y(_01863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19282_ (.A1(_02810_),
    .A2(_03049_),
    .B1(_10684_),
    .B2(_10413_),
    .X(_10416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19283_ (.A(_10416_),
    .Y(_10417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19284_ (.A1(_10679_),
    .A2(_10416_),
    .B1(_10678_),
    .B2(_10417_),
    .X(_01864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19285_ (.A(_10415_),
    .Y(_10418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _19286_ (.A(\design_top.IADDR[12] ),
    .B(_10418_),
    .Y(_10419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19287_ (.A1(\design_top.IADDR[12] ),
    .A2(_10418_),
    .B1(_10419_),
    .X(_01866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _19288_ (.A1(_10405_),
    .A2(_10730_),
    .B1(_10690_),
    .Y(_10420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19289_ (.A(_10420_),
    .Y(_10421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19290_ (.A1(_10674_),
    .A2(_10421_),
    .B1(_10673_),
    .B2(_10420_),
    .X(_01868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19291_ (.A(_10419_),
    .Y(_10422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _19292_ (.A(\design_top.IADDR[13] ),
    .B(_10422_),
    .Y(_10423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19293_ (.A1(\design_top.IADDR[13] ),
    .A2(_10422_),
    .B1(_10423_),
    .X(_01870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19294_ (.A(_01471_),
    .Y(_01871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19295_ (.A1(_02798_),
    .A2(_03033_),
    .B1(_10674_),
    .B2(_10421_),
    .X(_10424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19296_ (.A(_10424_),
    .Y(_10425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19297_ (.A1(_10669_),
    .A2(_10424_),
    .B1(_10668_),
    .B2(_10425_),
    .X(_01872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19298_ (.A(_10423_),
    .Y(_10426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _19299_ (.A(\design_top.IADDR[14] ),
    .B(_10426_),
    .Y(_10427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19300_ (.A1(\design_top.IADDR[14] ),
    .A2(_10426_),
    .B1(_10427_),
    .X(_01874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19301_ (.A(_01498_),
    .Y(_01875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _19302_ (.A1(_10669_),
    .A2(_10674_),
    .A3(_10421_),
    .B1(_10733_),
    .X(_10428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19303_ (.A(_10428_),
    .Y(_10429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19304_ (.A1(_10666_),
    .A2(_10428_),
    .B1(_10665_),
    .B2(_10429_),
    .X(_01876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19305_ (.A(_10427_),
    .Y(_10430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _19306_ (.A(\design_top.IADDR[15] ),
    .B(_10430_),
    .Y(_10431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19307_ (.A1(\design_top.IADDR[15] ),
    .A2(_10430_),
    .B1(_10431_),
    .X(_01878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19308_ (.A(_01514_),
    .Y(_01879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19309_ (.A1(_02786_),
    .A2(_03016_),
    .B1(_10666_),
    .B2(_10428_),
    .X(_10432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19310_ (.A(_10432_),
    .Y(_10433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19311_ (.A1(_10660_),
    .A2(_10432_),
    .B1(_10659_),
    .B2(_10433_),
    .X(_01880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19312_ (.A(_10431_),
    .Y(_10434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _19313_ (.A(\design_top.IADDR[16] ),
    .B(_10434_),
    .Y(_10435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19314_ (.A1(\design_top.IADDR[16] ),
    .A2(_10434_),
    .B1(_10435_),
    .X(_01882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19315_ (.A(_10739_),
    .X(_10436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19316_ (.A(_10436_),
    .Y(_10437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19317_ (.A1(_10436_),
    .A2(_10742_),
    .B1(_10437_),
    .B2(_10741_),
    .X(_01884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19318_ (.A(_10435_),
    .Y(_10438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _19319_ (.A(\design_top.IADDR[17] ),
    .B(_10438_),
    .Y(_10439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19320_ (.A1(\design_top.IADDR[17] ),
    .A2(_10438_),
    .B1(_10439_),
    .X(_01886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19321_ (.A1(_02774_),
    .A2(_02999_),
    .B1(_10436_),
    .B2(_10742_),
    .X(_10440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19322_ (.A(_10440_),
    .Y(_10441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19323_ (.A1(_10745_),
    .A2(_10440_),
    .B1(_10744_),
    .B2(_10441_),
    .X(_01888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19324_ (.A(\design_top.IADDR[18] ),
    .Y(_10442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19325_ (.A(_10442_),
    .B(_10439_),
    .Y(_10443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _19326_ (.A1(_10442_),
    .A2(_10439_),
    .B1(_10443_),
    .Y(_01890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19327_ (.A(_01579_),
    .Y(_01891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _19328_ (.A1(_10742_),
    .A2(_10745_),
    .A3(_10436_),
    .B1(_10652_),
    .X(_10444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19329_ (.A(_10444_),
    .Y(_10445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19330_ (.A1(_10646_),
    .A2(_10444_),
    .B1(_10645_),
    .B2(_10445_),
    .X(_01892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _19331_ (.A(_10439_),
    .B(_10442_),
    .C_N(\design_top.IADDR[19] ),
    .X(_10446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19332_ (.A1(\design_top.IADDR[19] ),
    .A2(_10443_),
    .B1(_10446_),
    .X(_01894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19333_ (.A(_01598_),
    .Y(_01895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19334_ (.A1(_02762_),
    .A2(_02982_),
    .B1(_10646_),
    .B2(_10444_),
    .X(_10447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19335_ (.A(_10447_),
    .Y(_10448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19336_ (.A1(_10649_),
    .A2(_10447_),
    .B1(_10648_),
    .B2(_10448_),
    .X(_01896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19337_ (.A(_10446_),
    .Y(_10449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _19338_ (.A(\design_top.IADDR[20] ),
    .B(_10449_),
    .Y(_10450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19339_ (.A1(\design_top.IADDR[20] ),
    .A2(_10449_),
    .B1(_10450_),
    .X(_01898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _19340_ (.A1(_10436_),
    .A2(_10746_),
    .B1(_10656_),
    .Y(_10451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19341_ (.A(_10451_),
    .Y(_10452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19342_ (.A1(_10627_),
    .A2(_10452_),
    .B1(_10626_),
    .B2(_10451_),
    .X(_01900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19343_ (.A(_10450_),
    .Y(_10453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _19344_ (.A(\design_top.IADDR[21] ),
    .B(_10453_),
    .Y(_10454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19345_ (.A1(\design_top.IADDR[21] ),
    .A2(_10453_),
    .B1(_10454_),
    .X(_01902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19346_ (.A(_01640_),
    .Y(_01903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19347_ (.A1(_02750_),
    .A2(_02965_),
    .B1(_10627_),
    .B2(_10452_),
    .X(_10455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19348_ (.A(_10455_),
    .Y(_10456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19349_ (.A1(_10631_),
    .A2(_10455_),
    .B1(_10630_),
    .B2(_10456_),
    .X(_01904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19350_ (.A(_10454_),
    .Y(_10457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _19351_ (.A(\design_top.IADDR[22] ),
    .B(_10457_),
    .Y(_10458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19352_ (.A1(\design_top.IADDR[22] ),
    .A2(_10457_),
    .B1(_10458_),
    .X(_01906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19353_ (.A(_01662_),
    .Y(_01907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _19354_ (.A1(_10627_),
    .A2(_10631_),
    .A3(_10452_),
    .B1(_10749_),
    .X(_10459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19355_ (.A(_10459_),
    .Y(_10460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19356_ (.A1(_10637_),
    .A2(_10459_),
    .B1(_10636_),
    .B2(_10460_),
    .X(_01908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19357_ (.A(_10458_),
    .Y(_10461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _19358_ (.A(\design_top.IADDR[23] ),
    .B(_10461_),
    .Y(_10462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19359_ (.A1(\design_top.IADDR[23] ),
    .A2(_10461_),
    .B1(_10462_),
    .X(_01910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19360_ (.A(_01680_),
    .Y(_01911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19361_ (.A1(_02738_),
    .A2(_02948_),
    .B1(_10637_),
    .B2(_10459_),
    .X(_10463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19362_ (.A(_10463_),
    .Y(_10464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19363_ (.A1(_10641_),
    .A2(_10463_),
    .B1(_10640_),
    .B2(_10464_),
    .X(_01912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19364_ (.A(\design_top.IADDR[24] ),
    .Y(_10465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19365_ (.A(_10465_),
    .B(_10462_),
    .Y(_10466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _19366_ (.A1(_10465_),
    .A2(_10462_),
    .B1(_10466_),
    .Y(_01914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19367_ (.A(_10753_),
    .Y(_10467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19368_ (.A1(_10753_),
    .A2(_10615_),
    .B1(_10467_),
    .B2(_10614_),
    .X(_01916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _19369_ (.A(_10462_),
    .B(_10465_),
    .C_N(\design_top.IADDR[25] ),
    .X(_10468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19370_ (.A1(\design_top.IADDR[25] ),
    .A2(_10466_),
    .B1(_10468_),
    .X(_01918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19371_ (.A1(_02726_),
    .A2(_02931_),
    .B1(_10753_),
    .B2(_10615_),
    .X(_10469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19372_ (.A(_10469_),
    .Y(_10470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19373_ (.A1(_10612_),
    .A2(_10469_),
    .B1(_10611_),
    .B2(_10470_),
    .X(_01920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19374_ (.A(\design_top.IADDR[26] ),
    .Y(_10471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19375_ (.A(_10471_),
    .B(_10468_),
    .Y(_10472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _19376_ (.A1(_10471_),
    .A2(_10468_),
    .B1(_10472_),
    .Y(_01922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19377_ (.A(_01744_),
    .Y(_01923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _19378_ (.A1(_10612_),
    .A2(_10615_),
    .A3(_10753_),
    .B1(_10755_),
    .X(_10473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _19379_ (.A1_N(_10622_),
    .A2_N(_10473_),
    .B1(_10622_),
    .B2(_10473_),
    .Y(_01924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _19380_ (.A(_10468_),
    .B(_10471_),
    .C_N(\design_top.IADDR[27] ),
    .X(_10474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19381_ (.A1(\design_top.IADDR[27] ),
    .A2(_10472_),
    .B1(_10474_),
    .X(_01926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19382_ (.A(_01763_),
    .Y(_01927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19383_ (.A1(_02714_),
    .A2(_02914_),
    .B1(_10622_),
    .B2(_10473_),
    .X(_10475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _19384_ (.A1_N(_10618_),
    .A2_N(_10475_),
    .B1(_10618_),
    .B2(_10475_),
    .Y(_01928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19385_ (.A(_10474_),
    .Y(_10476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _19386_ (.A(\design_top.IADDR[28] ),
    .B(_10476_),
    .Y(_10477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19387_ (.A1(\design_top.IADDR[28] ),
    .A2(_10476_),
    .B1(_10477_),
    .X(_01930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19388_ (.A(_10759_),
    .Y(_10478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19389_ (.A1(_10759_),
    .A2(_10608_),
    .B1(_10478_),
    .B2(_10607_),
    .X(_01932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19390_ (.A(_10477_),
    .Y(_10479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _19391_ (.A(\design_top.IADDR[29] ),
    .B(_10479_),
    .Y(_10480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19392_ (.A1(\design_top.IADDR[29] ),
    .A2(_10479_),
    .B1(_10480_),
    .X(_01934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19393_ (.A1(_02702_),
    .A2(_02897_),
    .B1(_10759_),
    .B2(_10608_),
    .X(_10481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19394_ (.A(_10481_),
    .Y(_10482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19395_ (.A1(_10603_),
    .A2(_10481_),
    .B1(_10602_),
    .B2(_10482_),
    .X(_01936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19396_ (.A(_10480_),
    .Y(_10483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _19397_ (.A(\design_top.IADDR[30] ),
    .B(_10483_),
    .Y(_10484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19398_ (.A1(\design_top.IADDR[30] ),
    .A2(_10483_),
    .B1(_10484_),
    .X(_01938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19399_ (.A(_01826_),
    .Y(_01939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _19400_ (.A1_N(_10599_),
    .A2_N(_10762_),
    .B1(_10599_),
    .B2(_10762_),
    .Y(_01940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19401_ (.A(\design_top.IADDR[31] ),
    .Y(_10485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a32o_2 _19402_ (.A1(\design_top.IADDR[30] ),
    .A2(_10483_),
    .A3(_10485_),
    .B1(\design_top.IADDR[31] ),
    .B2(_10484_),
    .X(_01942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19403_ (.A(_00858_),
    .Y(_01943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _19404_ (.A(_08617_),
    .B(\design_top.uart0.UART_XSTATE[3] ),
    .C(_08618_),
    .D(_08612_),
    .X(_01945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19405_ (.A(\design_top.TIMER[0] ),
    .Y(_01950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19406_ (.A1(\design_top.TIMER[1] ),
    .A2(\design_top.TIMER[0] ),
    .B1_N(_10847_),
    .X(_01951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19407_ (.A1(\design_top.TIMER[2] ),
    .A2(_10847_),
    .B1_N(_10848_),
    .X(_01952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19408_ (.A1(\design_top.TIMER[3] ),
    .A2(_10848_),
    .B1_N(_10849_),
    .X(_01953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19409_ (.A1(\design_top.TIMER[4] ),
    .A2(_10849_),
    .B1_N(_10850_),
    .X(_01954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19410_ (.A1(\design_top.TIMER[5] ),
    .A2(_10850_),
    .B1_N(_10851_),
    .X(_01955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19411_ (.A1(\design_top.TIMER[6] ),
    .A2(_10851_),
    .B1_N(_10852_),
    .X(_01956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19412_ (.A1(\design_top.TIMER[7] ),
    .A2(_10852_),
    .B1_N(_10853_),
    .X(_01957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19413_ (.A1(\design_top.TIMER[8] ),
    .A2(_10853_),
    .B1_N(_10854_),
    .X(_01958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19414_ (.A1(\design_top.TIMER[9] ),
    .A2(_10854_),
    .B1_N(_10855_),
    .X(_01959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19415_ (.A1(\design_top.TIMER[10] ),
    .A2(_10855_),
    .B1_N(_10856_),
    .X(_01960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19416_ (.A1(\design_top.TIMER[11] ),
    .A2(_10856_),
    .B1_N(_10857_),
    .X(_01961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19417_ (.A1(\design_top.TIMER[12] ),
    .A2(_10857_),
    .B1_N(_10858_),
    .X(_01962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19418_ (.A1(\design_top.TIMER[13] ),
    .A2(_10858_),
    .B1_N(_10859_),
    .X(_01963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19419_ (.A1(\design_top.TIMER[14] ),
    .A2(_10859_),
    .B1_N(_10860_),
    .X(_01964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19420_ (.A1(\design_top.TIMER[15] ),
    .A2(_10860_),
    .B1_N(_10861_),
    .X(_01965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19421_ (.A(\design_top.TIMER[16] ),
    .B(_10861_),
    .X(_10486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19422_ (.A1(\design_top.TIMER[16] ),
    .A2(_10861_),
    .B1_N(_10486_),
    .X(_01966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19423_ (.A(\design_top.TIMER[17] ),
    .B(_10486_),
    .X(_10487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19424_ (.A1(\design_top.TIMER[17] ),
    .A2(_10486_),
    .B1_N(_10487_),
    .X(_01967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19425_ (.A(\design_top.TIMER[18] ),
    .B(_10487_),
    .X(_10488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19426_ (.A1(\design_top.TIMER[18] ),
    .A2(_10487_),
    .B1_N(_10488_),
    .X(_01968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19427_ (.A1(\design_top.TIMER[19] ),
    .A2(_10488_),
    .B1_N(_10862_),
    .X(_01969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19428_ (.A(\design_top.TIMER[20] ),
    .B(_10862_),
    .X(_10489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19429_ (.A1(\design_top.TIMER[20] ),
    .A2(_10862_),
    .B1_N(_10489_),
    .X(_01970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19430_ (.A1(\design_top.TIMER[21] ),
    .A2(_10489_),
    .B1_N(_10863_),
    .X(_01971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19431_ (.A(\design_top.TIMER[22] ),
    .B(_10863_),
    .X(_10490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19432_ (.A1(\design_top.TIMER[22] ),
    .A2(_10863_),
    .B1_N(_10490_),
    .X(_01972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19433_ (.A1(\design_top.TIMER[23] ),
    .A2(_10490_),
    .B1_N(_10864_),
    .X(_01973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19434_ (.A(\design_top.TIMER[24] ),
    .B(_10864_),
    .Y(_10491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _19435_ (.A1(\design_top.TIMER[24] ),
    .A2(_10864_),
    .B1(_10491_),
    .X(_01974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19436_ (.A(\design_top.TIMER[25] ),
    .Y(_10492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _19437_ (.A1(_10492_),
    .A2(_10491_),
    .B1(_10865_),
    .Y(_01975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19438_ (.A1(\design_top.TIMER[26] ),
    .A2(_10865_),
    .B1_N(_10866_),
    .X(_01976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19439_ (.A1(\design_top.TIMER[27] ),
    .A2(_10866_),
    .B1_N(_10867_),
    .X(_01977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19440_ (.A(\design_top.TIMER[28] ),
    .B(_10867_),
    .X(_10493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19441_ (.A1(\design_top.TIMER[28] ),
    .A2(_10867_),
    .B1_N(_10493_),
    .X(_01978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19442_ (.A(\design_top.TIMER[29] ),
    .B(_10493_),
    .X(_10494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _19443_ (.A1(\design_top.TIMER[29] ),
    .A2(_10493_),
    .B1_N(_10494_),
    .X(_01979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19444_ (.A1_N(\design_top.TIMER[30] ),
    .A2_N(_10494_),
    .B1(\design_top.TIMER[30] ),
    .B2(_10494_),
    .X(_01980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19445_ (.A1(\design_top.TIMER[30] ),
    .A2(_10494_),
    .B1(\design_top.TIMER[31] ),
    .X(_10495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19446_ (.A(_03197_),
    .B(_10495_),
    .X(_01981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19447_ (.A1(\design_top.core0.XJALR ),
    .A2(\design_top.core0.XJAL ),
    .B1(_02661_),
    .X(_02870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19448_ (.A(_08599_),
    .B(_02849_),
    .Y(_02848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _19449_ (.A(_08502_),
    .B(_09914_),
    .C(_09913_),
    .X(_03159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _19450_ (.A(_08502_),
    .B(\design_top.core0.FCT3[0] ),
    .C(\design_top.core0.FCT3[2] ),
    .X(_03161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19451_ (.A(_09913_),
    .B(_02854_),
    .Y(_02852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19452_ (.A(_08599_),
    .B(_02854_),
    .Y(_02853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _19453_ (.A1(_10082_),
    .A2(_09954_),
    .B1(_00938_),
    .Y(_00940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _19454_ (.A(_08564_),
    .B(_08598_),
    .C_N(_00940_),
    .X(_03189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19455_ (.A(_10628_),
    .X(_02956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _19456_ (.A(_10743_),
    .X(_02990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _19457_ (.A1(_03077_),
    .A2(_00809_),
    .B1(_03086_),
    .B2(_03081_),
    .X(_10496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _19458_ (.A1(_03093_),
    .A2(_00811_),
    .B1(_03102_),
    .B2(_03097_),
    .X(_10497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _19459_ (.A1(_03110_),
    .A2(_10717_),
    .B1(_03119_),
    .B2(_10770_),
    .X(_10498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _19460_ (.A1(_09947_),
    .A2(_10691_),
    .B1(_09950_),
    .B2(_10696_),
    .X(_10499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19461_ (.A1(_03110_),
    .A2(_10717_),
    .B1(_03102_),
    .B2(_03097_),
    .X(_10500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19462_ (.A1(_03134_),
    .A2(_10822_),
    .B1(_03127_),
    .B2(_10713_),
    .X(_10501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4bb_2 _19463_ (.A(_10498_),
    .B(_10499_),
    .C_N(_10500_),
    .D_N(_10501_),
    .X(_10502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19464_ (.A(_09941_),
    .B(_02641_),
    .Y(_10503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _19465_ (.A1(_03134_),
    .A2(_10822_),
    .B1(_10503_),
    .Y(_10504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _19466_ (.A1(_03119_),
    .A2(_10770_),
    .B1(_03077_),
    .B2(_00809_),
    .C1(_10504_),
    .X(_10505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4b_2 _19467_ (.A(_10496_),
    .B(_10497_),
    .C(_10502_),
    .D_N(_10505_),
    .X(_10506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _19468_ (.A1(_02956_),
    .A2(_02961_),
    .B1(_10624_),
    .B2(_02970_),
    .X(_10507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _19469_ (.A1(_02995_),
    .A2(_02990_),
    .B1(_02999_),
    .B2(_03004_),
    .X(_10508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19470_ (.A1(_02956_),
    .A2(_02961_),
    .B1(_10740_),
    .B2(_03004_),
    .X(_10509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221ai_2 _19471_ (.A1(_10624_),
    .A2(_02970_),
    .B1(_02995_),
    .B2(_02990_),
    .C1(_10509_),
    .Y(_10510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19472_ (.A(_02978_),
    .Y(_10511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19473_ (.A(_02978_),
    .B(_02973_),
    .X(_10512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _19474_ (.A1(_10021_),
    .A2(_02987_),
    .B1_N(_10512_),
    .Y(_10513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _19475_ (.A1(_10511_),
    .A2(_08541_),
    .B1(_10021_),
    .B2(_02987_),
    .C1(_10513_),
    .X(_10514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19476_ (.A(_02944_),
    .Y(_10515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22oi_2 _19477_ (.A1(_10010_),
    .A2(_10515_),
    .B1(_10006_),
    .B2(_02953_),
    .Y(_10516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _19478_ (.A1(_10010_),
    .A2(_10515_),
    .B1(_10006_),
    .B2(_02953_),
    .C1(_10516_),
    .X(_10517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _19479_ (.A(_10514_),
    .B(_10517_),
    .Y(_10518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _19480_ (.A(_10507_),
    .B(_10508_),
    .C(_10510_),
    .D(_10518_),
    .X(_10519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _19481_ (.A1(_02922_),
    .A2(_02927_),
    .B1(_02931_),
    .B2(_02936_),
    .X(_10520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _19482_ (.A1(_10598_),
    .A2(_02884_),
    .B1(_02888_),
    .B2(_02893_),
    .Y(_10521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19483_ (.A(_02884_),
    .Y(_10522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22oi_2 _19484_ (.A1(_02888_),
    .A2(_02893_),
    .B1(_02897_),
    .B2(_02902_),
    .Y(_10523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221ai_2 _19485_ (.A1(_02931_),
    .A2(_02936_),
    .B1(_10597_),
    .B2(_10522_),
    .C1(_10523_),
    .Y(_10524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19486_ (.A(_02684_),
    .B(_02875_),
    .Y(_10525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _19487_ (.A1(_10083_),
    .A2(_02875_),
    .B1(_10525_),
    .X(_10526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _19488_ (.A1(_02905_),
    .A2(_02910_),
    .B1(_10604_),
    .B2(_02902_),
    .Y(_10527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _19489_ (.A1(_02905_),
    .A2(_02910_),
    .B1(_10756_),
    .B2(_02919_),
    .X(_10528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19490_ (.A1(_02914_),
    .A2(_02919_),
    .B1(_02922_),
    .B2(_02927_),
    .X(_10529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4b_2 _19491_ (.A(_10526_),
    .B(_10527_),
    .C(_10528_),
    .D_N(_10529_),
    .X(_10530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _19492_ (.A(_10520_),
    .B(_10521_),
    .C(_10524_),
    .D(_10530_),
    .X(_10531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _19493_ (.A1(_03012_),
    .A2(_10032_),
    .B1(_03021_),
    .B2(_10734_),
    .X(_10532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _19494_ (.A1(_10216_),
    .A2(_10682_),
    .B1(_08590_),
    .B2(_10215_),
    .X(_10533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _19495_ (.A1(_03029_),
    .A2(_03024_),
    .B1(_03038_),
    .B2(_10043_),
    .X(_10534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19496_ (.A1(_03029_),
    .A2(_03024_),
    .B1(_03021_),
    .B2(_03016_),
    .X(_10535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4b_2 _19497_ (.A(_10532_),
    .B(_10533_),
    .C(_10534_),
    .D_N(_10535_),
    .X(_10536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19498_ (.A1(_10676_),
    .A2(_10218_),
    .B1(_10216_),
    .B2(_10682_),
    .X(_10537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19499_ (.A1(_03070_),
    .A2(_03065_),
    .B1(_00803_),
    .B2(_03045_),
    .X(_10538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _19500_ (.A1(_03012_),
    .A2(_03007_),
    .B1(_03038_),
    .B2(_10043_),
    .C1(_10538_),
    .X(_10539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19501_ (.A1(_10214_),
    .A2(_10685_),
    .B1(_08590_),
    .B2(_10215_),
    .X(_10540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and4b_2 _19502_ (.A_N(_10536_),
    .B(_10537_),
    .C(_10539_),
    .D(_10540_),
    .X(_10541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4b_2 _19503_ (.A(_10506_),
    .B(_10519_),
    .C(_10531_),
    .D_N(_10541_),
    .X(_10542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19504_ (.A(_02875_),
    .Y(_10543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211ai_2 _19505_ (.A1(_02939_),
    .A2(_02944_),
    .B1(_02948_),
    .C1(_02953_),
    .Y(_10544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _19506_ (.A1(_02995_),
    .A2(_02990_),
    .B1(_10508_),
    .C1(_10514_),
    .X(_10545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a32o_2 _19507_ (.A1(_02982_),
    .A2(_02987_),
    .A3(_10512_),
    .B1(_02978_),
    .B2(_02973_),
    .X(_10546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19508_ (.A1(_02965_),
    .A2(_02970_),
    .B1(_10545_),
    .B2(_10546_),
    .X(_10547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221ai_2 _19509_ (.A1(_02956_),
    .A2(_02961_),
    .B1(_10507_),
    .B2(_10547_),
    .C1(_10517_),
    .Y(_10548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _19510_ (.A1(_10533_),
    .A2(_10540_),
    .B1(_10537_),
    .Y(_10549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _19511_ (.A1(_00803_),
    .A2(_03045_),
    .B1(_03038_),
    .B2(_03033_),
    .C1(_10549_),
    .X(_10550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19512_ (.A1(_10534_),
    .A2(_10550_),
    .B1(_10535_),
    .X(_10551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19513_ (.A1(_03012_),
    .A2(_03007_),
    .B1(_10532_),
    .B2(_10551_),
    .X(_10552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19514_ (.A1(_03119_),
    .A2(_10770_),
    .B1(_10503_),
    .B2(_10501_),
    .X(_10553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19515_ (.A1(_10498_),
    .A2(_10553_),
    .B1(_10500_),
    .X(_10554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ba_2 _19516_ (.A1(_10497_),
    .A2(_10554_),
    .B1_N(_10499_),
    .X(_10555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _19517_ (.A1(_03077_),
    .A2(_00809_),
    .B1(_10496_),
    .B2(_10555_),
    .C1(_10541_),
    .X(_10556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21bai_2 _19518_ (.A1(_10552_),
    .A2(_10556_),
    .B1_N(_10519_),
    .Y(_10557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2111a_2 _19519_ (.A1(_10010_),
    .A2(_10515_),
    .B1(_10544_),
    .C1(_10548_),
    .D1(_10557_),
    .X(_10558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _19520_ (.A1(_10520_),
    .A2(_10529_),
    .B1(_10528_),
    .Y(_10559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _19521_ (.A1(_10527_),
    .A2(_10559_),
    .B1(_10523_),
    .X(_10560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _19522_ (.A1(_10597_),
    .A2(_10522_),
    .B1(_10521_),
    .B2(_10560_),
    .Y(_10561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _19523_ (.A1(_10083_),
    .A2(_02875_),
    .B1(_10561_),
    .Y(_10562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221ai_2 _19524_ (.A1(_10078_),
    .A2(_10543_),
    .B1(_10531_),
    .B2(_10558_),
    .C1(_10562_),
    .Y(_10563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _19525_ (.A(_10542_),
    .B(_10563_),
    .X(_03160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2b_2 _19526_ (.A(_09991_),
    .B_N(_10081_),
    .X(_10564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _19527_ (.A(_09993_),
    .B(_09995_),
    .C(_10564_),
    .X(_10565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _19528_ (.A1(_03139_),
    .A2(_02879_),
    .A3(_10080_),
    .B1(_10083_),
    .B2(_03138_),
    .X(_10566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221ai_2 _19529_ (.A1(_10075_),
    .A2(_10564_),
    .B1(_10073_),
    .B2(_10565_),
    .C1(_10566_),
    .Y(_03158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _19530_ (.A1(_10078_),
    .A2(_10543_),
    .B1(_10525_),
    .B2(_10563_),
    .C1(_10542_),
    .X(_03137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19531_ (.A1(_03039_),
    .A2(_03033_),
    .B1(_08573_),
    .B2(_10337_),
    .X(_10567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19532_ (.A1(_03030_),
    .A2(_03024_),
    .B1(_08568_),
    .B2(_10567_),
    .X(_10568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19533_ (.A1(_03022_),
    .A2(_03016_),
    .B1(_08566_),
    .B2(_10568_),
    .X(_10569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19534_ (.A1(_03013_),
    .A2(_03007_),
    .B1(_08571_),
    .B2(_10569_),
    .X(_10570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19535_ (.A(_02876_),
    .Y(_10571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _19536_ (.A(_08555_),
    .Y(_10572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _19537_ (.A1(_02937_),
    .A2(_10613_),
    .A3(_08552_),
    .B1(_02928_),
    .B2(_02922_),
    .X(_10573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19538_ (.A1(_02920_),
    .A2(_10756_),
    .B1(_10572_),
    .B2(_10573_),
    .X(_10574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19539_ (.A1(_02911_),
    .A2(_02905_),
    .B1(_08550_),
    .B2(_10574_),
    .X(_10575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19540_ (.A1(_02903_),
    .A2(_10604_),
    .B1(_08561_),
    .B2(_10575_),
    .X(_10576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19541_ (.A1(_02894_),
    .A2(_02888_),
    .B1(_08560_),
    .B2(_10576_),
    .X(_10577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19542_ (.A1(_02885_),
    .A2(_02879_),
    .B1(_08557_),
    .B2(_10577_),
    .X(_10578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _19543_ (.A1(_03005_),
    .A2(_02999_),
    .A3(_08540_),
    .B1(_02996_),
    .B2(_02990_),
    .X(_10579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19544_ (.A1(_02988_),
    .A2(_02982_),
    .B1(_08545_),
    .B2(_10579_),
    .X(_10580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19545_ (.A1(_02979_),
    .A2(_02973_),
    .B1(_08542_),
    .B2(_10580_),
    .X(_10581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _19546_ (.A1(_02971_),
    .A2(_02965_),
    .A3(_08532_),
    .B1(_02962_),
    .B2(_02956_),
    .X(_10582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19547_ (.A1(_02954_),
    .A2(_02948_),
    .B1(_08537_),
    .B2(_10582_),
    .X(_10583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19548_ (.A(_08530_),
    .B(_10583_),
    .X(_10584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _19549_ (.A1(_02945_),
    .A2(_02939_),
    .B1(_08538_),
    .B2(_10581_),
    .C1(_10584_),
    .X(_10585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _19550_ (.A1(_08558_),
    .A2(_10578_),
    .B1(_08563_),
    .B2(_10585_),
    .X(_10586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221ai_2 _19551_ (.A1(_08564_),
    .A2(_10570_),
    .B1(_10078_),
    .B2(_10571_),
    .C1(_10586_),
    .Y(_03136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19552_ (.A(_09937_),
    .B(_02849_),
    .Y(_02851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19553_ (.A(_10085_),
    .B(_09962_),
    .Y(_03121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19554_ (.A(_10088_),
    .B(_10693_),
    .Y(_03104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19555_ (.A(_03071_),
    .B(_10685_),
    .Y(_03072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19556_ (.A(_03039_),
    .B(_10672_),
    .Y(_03040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19557_ (.A(_03005_),
    .B(_08546_),
    .Y(_03006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19558_ (.A(_02971_),
    .B(_08533_),
    .Y(_02972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19559_ (.A(_02937_),
    .B(_08553_),
    .Y(_02938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19560_ (.A(_02885_),
    .B(_10597_),
    .Y(_02886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _19561_ (.A(_10083_),
    .B(_10571_),
    .X(_02878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _19562_ (.A(_08486_),
    .B(_10595_),
    .Y(_02869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2b_2 _19563_ (.A_N(\design_top.uart0.UART_RXDFF[1] ),
    .B(_09845_),
    .Y(_02625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _19564_ (.A1_N(_10954_),
    .A2_N(_10785_),
    .B1(\design_top.MEM[0][15] ),
    .B2(_10800_),
    .X(_07431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19565_ (.LO(io_oeb[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19566_ (.LO(io_oeb[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19567_ (.LO(io_oeb[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19568_ (.LO(io_oeb[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19569_ (.LO(io_oeb[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19570_ (.LO(io_oeb[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19571_ (.LO(io_oeb[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19572_ (.LO(io_oeb[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19573_ (.LO(io_oeb[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19574_ (.LO(io_oeb[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19575_ (.LO(io_oeb[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19576_ (.LO(io_oeb[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19577_ (.LO(io_oeb[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19578_ (.LO(io_oeb[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19579_ (.LO(io_oeb[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19580_ (.LO(io_oeb[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19581_ (.LO(io_oeb[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19582_ (.LO(io_oeb[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19583_ (.LO(io_oeb[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19584_ (.LO(io_oeb[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19585_ (.LO(io_oeb[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19586_ (.LO(io_oeb[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19587_ (.LO(io_oeb[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19588_ (.LO(io_oeb[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19589_ (.LO(io_oeb[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19590_ (.LO(io_oeb[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19591_ (.LO(io_oeb[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19592_ (.LO(io_oeb[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19593_ (.LO(io_oeb[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19594_ (.LO(io_oeb[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19595_ (.LO(io_oeb[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19596_ (.LO(io_oeb[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19597_ (.LO(io_oeb[32]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19598_ (.LO(io_oeb[33]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19599_ (.LO(io_oeb[34]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19600_ (.LO(io_oeb[35]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19601_ (.LO(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19602_ (.LO(io_oeb[37]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19603_ (.LO(io_out[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19604_ (.LO(io_out[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19605_ (.LO(io_out[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19606_ (.LO(io_out[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19607_ (.LO(io_out[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19608_ (.LO(io_out[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19609_ (.LO(io_out[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19610_ (.LO(io_out[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19611_ (.LO(io_out[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19612_ (.LO(io_out[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19613_ (.LO(io_out[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19614_ (.LO(io_out[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19615_ (.LO(io_out[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19616_ (.LO(io_out[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19617_ (.LO(io_out[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19618_ (.LO(io_out[32]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19619_ (.LO(io_out[33]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19620_ (.LO(io_out[34]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19621_ (.LO(io_out[35]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19622_ (.LO(io_out[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19623_ (.LO(io_out[37]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19624_ (.LO(la_data_out[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19625_ (.LO(la_data_out[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19626_ (.LO(la_data_out[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19627_ (.LO(la_data_out[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19628_ (.LO(la_data_out[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19629_ (.LO(la_data_out[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19630_ (.LO(la_data_out[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19631_ (.LO(la_data_out[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19632_ (.LO(la_data_out[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19633_ (.LO(la_data_out[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19634_ (.LO(la_data_out[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19635_ (.LO(la_data_out[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19636_ (.LO(la_data_out[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19637_ (.LO(la_data_out[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19638_ (.LO(la_data_out[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19639_ (.LO(la_data_out[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19640_ (.LO(la_data_out[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19641_ (.LO(la_data_out[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19642_ (.LO(la_data_out[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19643_ (.LO(la_data_out[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19644_ (.LO(la_data_out[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19645_ (.LO(la_data_out[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19646_ (.LO(la_data_out[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19647_ (.LO(la_data_out[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19648_ (.LO(la_data_out[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19649_ (.LO(la_data_out[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19650_ (.LO(la_data_out[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19651_ (.LO(la_data_out[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19652_ (.LO(la_data_out[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19653_ (.LO(la_data_out[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19654_ (.LO(la_data_out[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19655_ (.LO(la_data_out[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19656_ (.LO(la_data_out[32]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19657_ (.LO(la_data_out[33]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19658_ (.LO(la_data_out[34]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19659_ (.LO(la_data_out[35]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19660_ (.LO(la_data_out[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19661_ (.LO(la_data_out[37]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19662_ (.LO(la_data_out[38]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19663_ (.LO(la_data_out[39]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19664_ (.LO(la_data_out[40]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19665_ (.LO(la_data_out[41]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19666_ (.LO(la_data_out[42]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19667_ (.LO(la_data_out[43]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19668_ (.LO(la_data_out[44]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19669_ (.LO(la_data_out[45]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19670_ (.LO(la_data_out[46]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19671_ (.LO(la_data_out[47]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19672_ (.LO(la_data_out[48]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19673_ (.LO(la_data_out[49]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19674_ (.LO(la_data_out[50]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19675_ (.LO(la_data_out[51]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19676_ (.LO(la_data_out[52]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19677_ (.LO(la_data_out[53]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19678_ (.LO(la_data_out[54]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19679_ (.LO(la_data_out[55]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19680_ (.LO(la_data_out[56]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19681_ (.LO(la_data_out[57]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19682_ (.LO(la_data_out[58]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19683_ (.LO(la_data_out[59]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19684_ (.LO(la_data_out[60]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19685_ (.LO(la_data_out[61]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19686_ (.LO(la_data_out[62]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19687_ (.LO(la_data_out[63]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19688_ (.LO(la_data_out[64]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19689_ (.LO(la_data_out[65]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19690_ (.LO(la_data_out[66]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19691_ (.LO(la_data_out[67]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19692_ (.LO(la_data_out[68]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19693_ (.LO(la_data_out[69]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19694_ (.LO(la_data_out[70]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19695_ (.LO(la_data_out[71]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19696_ (.LO(la_data_out[72]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19697_ (.LO(la_data_out[73]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19698_ (.LO(la_data_out[74]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19699_ (.LO(la_data_out[75]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19700_ (.LO(la_data_out[76]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19701_ (.LO(la_data_out[77]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19702_ (.LO(la_data_out[78]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19703_ (.LO(la_data_out[79]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19704_ (.LO(la_data_out[80]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19705_ (.LO(la_data_out[81]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19706_ (.LO(la_data_out[82]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19707_ (.LO(la_data_out[83]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19708_ (.LO(la_data_out[84]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19709_ (.LO(la_data_out[85]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19710_ (.LO(la_data_out[86]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19711_ (.LO(la_data_out[87]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19712_ (.LO(la_data_out[88]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19713_ (.LO(la_data_out[89]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19714_ (.LO(la_data_out[90]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19715_ (.LO(la_data_out[91]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19716_ (.LO(la_data_out[92]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19717_ (.LO(la_data_out[93]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19718_ (.LO(la_data_out[94]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19719_ (.LO(la_data_out[95]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19720_ (.LO(la_data_out[96]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19721_ (.LO(la_data_out[97]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19722_ (.LO(la_data_out[98]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19723_ (.LO(la_data_out[99]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19724_ (.LO(la_data_out[100]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19725_ (.LO(la_data_out[101]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19726_ (.LO(la_data_out[102]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19727_ (.LO(la_data_out[103]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19728_ (.LO(la_data_out[104]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19729_ (.LO(la_data_out[105]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19730_ (.LO(la_data_out[106]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19731_ (.LO(la_data_out[107]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19732_ (.LO(la_data_out[108]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19733_ (.LO(la_data_out[109]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19734_ (.LO(la_data_out[110]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19735_ (.LO(la_data_out[111]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19736_ (.LO(la_data_out[112]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19737_ (.LO(la_data_out[113]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19738_ (.LO(la_data_out[114]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19739_ (.LO(la_data_out[115]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19740_ (.LO(la_data_out[116]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19741_ (.LO(la_data_out[117]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19742_ (.LO(la_data_out[118]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19743_ (.LO(la_data_out[119]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19744_ (.LO(la_data_out[120]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19745_ (.LO(la_data_out[121]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19746_ (.LO(la_data_out[122]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19747_ (.LO(la_data_out[123]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19748_ (.LO(la_data_out[124]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19749_ (.LO(la_data_out[125]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19750_ (.LO(la_data_out[126]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19751_ (.LO(la_data_out[127]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19752_ (.LO(user_irq[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19753_ (.LO(user_irq[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19754_ (.LO(user_irq[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19755_ (.LO(wbs_ack_o),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19756_ (.LO(wbs_dat_o[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19757_ (.LO(wbs_dat_o[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19758_ (.LO(wbs_dat_o[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19759_ (.LO(wbs_dat_o[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19760_ (.LO(wbs_dat_o[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19761_ (.LO(wbs_dat_o[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19762_ (.LO(wbs_dat_o[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19763_ (.LO(wbs_dat_o[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19764_ (.LO(wbs_dat_o[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19765_ (.LO(wbs_dat_o[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19766_ (.LO(wbs_dat_o[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19767_ (.LO(wbs_dat_o[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19768_ (.LO(wbs_dat_o[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19769_ (.LO(wbs_dat_o[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19770_ (.LO(wbs_dat_o[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19771_ (.LO(wbs_dat_o[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19772_ (.LO(wbs_dat_o[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19773_ (.LO(wbs_dat_o[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19774_ (.LO(wbs_dat_o[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19775_ (.LO(wbs_dat_o[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19776_ (.LO(wbs_dat_o[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19777_ (.LO(wbs_dat_o[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19778_ (.LO(wbs_dat_o[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19779_ (.LO(wbs_dat_o[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19780_ (.LO(wbs_dat_o[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19781_ (.LO(wbs_dat_o[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19782_ (.LO(wbs_dat_o[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19783_ (.LO(wbs_dat_o[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19784_ (.LO(wbs_dat_o[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19785_ (.LO(wbs_dat_o[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19786_ (.LO(wbs_dat_o[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _19787_ (.LO(wbs_dat_o[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _19788_ (.A(io_out[15]),
    .X(\design_top.GPIOFF[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _19789_ (.A(io_out[8]),
    .X(\design_top.LEDFF[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _19790_ (.A(io_out[9]),
    .X(\design_top.LEDFF[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _19791_ (.A(io_out[10]),
    .X(\design_top.LEDFF[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _19792_ (.A(io_out[11]),
    .X(\design_top.LEDFF[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _19793_ (.A(io_out[14]),
    .X(\design_top.XTIMER ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19794_ (.A0(_03161_),
    .A1(_02854_),
    .S(io_out[12]),
    .X(_11368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19795_ (.A0(_02847_),
    .A1(_00783_),
    .S(_02852_),
    .X(_11369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19796_ (.A0(\design_top.ROMFF[0] ),
    .A1(\design_top.ROMFF2[0] ),
    .S(\design_top.HLT2 ),
    .X(io_out[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19797_ (.A0(\design_top.ROMFF[1] ),
    .A1(\design_top.ROMFF2[1] ),
    .S(\design_top.HLT2 ),
    .X(io_out[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19798_ (.A0(\design_top.ROMFF[2] ),
    .A1(\design_top.ROMFF2[2] ),
    .S(\design_top.HLT2 ),
    .X(io_out[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19799_ (.A0(\design_top.ROMFF[3] ),
    .A1(\design_top.ROMFF2[3] ),
    .S(\design_top.HLT2 ),
    .X(io_out[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19800_ (.A0(_03134_),
    .A1(_00756_),
    .S(_02847_),
    .X(_00757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19801_ (.A0(_00757_),
    .A1(_00755_),
    .S(_02852_),
    .X(\design_top.DATAO[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19802_ (.A0(_03127_),
    .A1(_00759_),
    .S(_02847_),
    .X(_00760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19803_ (.A0(_00760_),
    .A1(_00758_),
    .S(_02852_),
    .X(\design_top.DATAO[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19804_ (.A0(_03119_),
    .A1(_00762_),
    .S(_02847_),
    .X(_00763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19805_ (.A0(_00763_),
    .A1(_00761_),
    .S(_02852_),
    .X(\design_top.DATAO[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19806_ (.A0(_03110_),
    .A1(_00765_),
    .S(_02847_),
    .X(_00766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19807_ (.A0(_00766_),
    .A1(_00764_),
    .S(_02852_),
    .X(\design_top.DATAO[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19808_ (.A0(_03102_),
    .A1(_00768_),
    .S(_02847_),
    .X(_00769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19809_ (.A0(_00769_),
    .A1(_00767_),
    .S(_02852_),
    .X(\design_top.DATAO[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19810_ (.A0(_03093_),
    .A1(_00771_),
    .S(_02847_),
    .X(_00772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19811_ (.A0(_00772_),
    .A1(_00770_),
    .S(_02852_),
    .X(\design_top.DATAO[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19812_ (.A0(_03086_),
    .A1(_00774_),
    .S(_02847_),
    .X(_00775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19813_ (.A0(_00775_),
    .A1(_00773_),
    .S(_02852_),
    .X(\design_top.DATAO[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19814_ (.A0(_03077_),
    .A1(_00777_),
    .S(_02847_),
    .X(_00778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19815_ (.A0(_00778_),
    .A1(_00776_),
    .S(_02852_),
    .X(\design_top.DATAO[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19816_ (.A0(_03070_),
    .A1(_00865_),
    .S(_02847_),
    .X(_00866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19817_ (.A0(_00866_),
    .A1(_00864_),
    .S(_02852_),
    .X(\design_top.DATAO[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19818_ (.A0(_03061_),
    .A1(_00868_),
    .S(_02847_),
    .X(_00869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19819_ (.A0(_00869_),
    .A1(_00867_),
    .S(_02852_),
    .X(\design_top.DATAO[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19820_ (.A0(_03054_),
    .A1(_00871_),
    .S(_02847_),
    .X(_00872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19821_ (.A0(_00872_),
    .A1(_00870_),
    .S(_02852_),
    .X(\design_top.DATAO[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19822_ (.A0(_03045_),
    .A1(_00874_),
    .S(_02847_),
    .X(_00875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19823_ (.A0(_00875_),
    .A1(_00873_),
    .S(_02852_),
    .X(\design_top.DATAO[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19824_ (.A0(_03038_),
    .A1(_00877_),
    .S(_02847_),
    .X(_00878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19825_ (.A0(_00878_),
    .A1(_00876_),
    .S(_02852_),
    .X(\design_top.DATAO[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19826_ (.A0(_03029_),
    .A1(_00880_),
    .S(_02847_),
    .X(_00881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19827_ (.A0(_00881_),
    .A1(_00879_),
    .S(_02852_),
    .X(\design_top.DATAO[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19828_ (.A0(_03021_),
    .A1(_00883_),
    .S(_02847_),
    .X(_00884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19829_ (.A0(_00884_),
    .A1(_00882_),
    .S(_02852_),
    .X(\design_top.DATAO[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19830_ (.A0(_03012_),
    .A1(_00886_),
    .S(_02847_),
    .X(_00887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19831_ (.A0(_00887_),
    .A1(_00885_),
    .S(_02852_),
    .X(\design_top.DATAO[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19832_ (.A0(_03004_),
    .A1(_00889_),
    .S(_02847_),
    .X(_00890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19833_ (.A0(_00890_),
    .A1(_00888_),
    .S(_02852_),
    .X(\design_top.DATAO[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19834_ (.A0(_02995_),
    .A1(_00892_),
    .S(_02847_),
    .X(_00893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19835_ (.A0(_00893_),
    .A1(_00891_),
    .S(_02852_),
    .X(\design_top.DATAO[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19836_ (.A0(_02987_),
    .A1(_00895_),
    .S(_02847_),
    .X(_00896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19837_ (.A0(_00896_),
    .A1(_00894_),
    .S(_02852_),
    .X(\design_top.DATAO[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19838_ (.A0(_02978_),
    .A1(_00898_),
    .S(_02847_),
    .X(_00899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19839_ (.A0(_00899_),
    .A1(_00897_),
    .S(_02852_),
    .X(\design_top.DATAO[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19840_ (.A0(_02970_),
    .A1(_00901_),
    .S(_02847_),
    .X(_00902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19841_ (.A0(_00902_),
    .A1(_00900_),
    .S(_02852_),
    .X(\design_top.DATAO[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19842_ (.A0(_02961_),
    .A1(_00904_),
    .S(_02847_),
    .X(_00905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19843_ (.A0(_00905_),
    .A1(_00903_),
    .S(_02852_),
    .X(\design_top.DATAO[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19844_ (.A0(_02953_),
    .A1(_00907_),
    .S(_02847_),
    .X(_00908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19845_ (.A0(_00908_),
    .A1(_00906_),
    .S(_02852_),
    .X(\design_top.DATAO[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19846_ (.A0(_02944_),
    .A1(_00910_),
    .S(_02847_),
    .X(_00911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19847_ (.A0(_00911_),
    .A1(_00909_),
    .S(_02852_),
    .X(\design_top.DATAO[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19848_ (.A0(_02936_),
    .A1(_00913_),
    .S(_02847_),
    .X(_00914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19849_ (.A0(_00914_),
    .A1(_00912_),
    .S(_02852_),
    .X(\design_top.DATAO[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19850_ (.A0(_02927_),
    .A1(_00916_),
    .S(_02847_),
    .X(_00917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19851_ (.A0(_00917_),
    .A1(_00915_),
    .S(_02852_),
    .X(\design_top.DATAO[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19852_ (.A0(_02919_),
    .A1(_00919_),
    .S(_02847_),
    .X(_00920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19853_ (.A0(_00920_),
    .A1(_00918_),
    .S(_02852_),
    .X(\design_top.DATAO[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19854_ (.A0(_02910_),
    .A1(_00922_),
    .S(_02847_),
    .X(_00923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19855_ (.A0(_00923_),
    .A1(_00921_),
    .S(_02852_),
    .X(\design_top.DATAO[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19856_ (.A0(_02902_),
    .A1(_00925_),
    .S(_02847_),
    .X(_00926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19857_ (.A0(_00926_),
    .A1(_00924_),
    .S(_02852_),
    .X(\design_top.DATAO[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19858_ (.A0(_02893_),
    .A1(_00928_),
    .S(_02847_),
    .X(_00929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19859_ (.A0(_00929_),
    .A1(_00927_),
    .S(_02852_),
    .X(\design_top.DATAO[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19860_ (.A0(_02884_),
    .A1(_00931_),
    .S(_02847_),
    .X(_00932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19861_ (.A0(_00932_),
    .A1(_00930_),
    .S(_02852_),
    .X(\design_top.DATAO[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19862_ (.A0(_02875_),
    .A1(_03268_),
    .S(_02847_),
    .X(_03269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19863_ (.A0(_03269_),
    .A1(_03267_),
    .S(_02852_),
    .X(\design_top.DATAO[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19864_ (.A0(\design_top.ROMFF[7] ),
    .A1(\design_top.ROMFF2[7] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19865_ (.A0(\design_top.ROMFF[8] ),
    .A1(\design_top.ROMFF2[8] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19866_ (.A0(\design_top.ROMFF[9] ),
    .A1(\design_top.ROMFF2[9] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19867_ (.A0(\design_top.ROMFF[10] ),
    .A1(\design_top.ROMFF2[10] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19868_ (.A0(\design_top.ROMFF[12] ),
    .A1(\design_top.ROMFF2[12] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19869_ (.A0(\design_top.ROMFF[13] ),
    .A1(\design_top.ROMFF2[13] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19870_ (.A0(\design_top.ROMFF[14] ),
    .A1(\design_top.ROMFF2[14] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19871_ (.A0(\design_top.ROMFF[15] ),
    .A1(\design_top.ROMFF2[15] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19872_ (.A0(\design_top.ROMFF[16] ),
    .A1(\design_top.ROMFF2[16] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19873_ (.A0(\design_top.ROMFF[17] ),
    .A1(\design_top.ROMFF2[17] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19874_ (.A0(\design_top.ROMFF[18] ),
    .A1(\design_top.ROMFF2[18] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19875_ (.A0(\design_top.ROMFF[20] ),
    .A1(\design_top.ROMFF2[20] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19876_ (.A0(\design_top.ROMFF[21] ),
    .A1(\design_top.ROMFF2[21] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19877_ (.A0(\design_top.ROMFF[22] ),
    .A1(\design_top.ROMFF2[22] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19878_ (.A0(\design_top.ROMFF[23] ),
    .A1(\design_top.ROMFF2[23] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19879_ (.A0(\design_top.ROMFF[30] ),
    .A1(\design_top.ROMFF2[30] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19880_ (.A0(\design_top.ROMFF[31] ),
    .A1(\design_top.ROMFF2[31] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19881_ (.A0(_01946_),
    .A1(_01947_),
    .S(\design_top.uart0.UART_XSTATE[2] ),
    .X(_01948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19882_ (.A0(_01945_),
    .A1(_01948_),
    .S(\design_top.uart0.UART_XSTATE[3] ),
    .X(io_out[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19883_ (.A0(_01949_),
    .A1(_02625_),
    .S(_02662_),
    .X(_02626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19884_ (.A0(_02623_),
    .A1(_00985_),
    .S(_02663_),
    .X(_02624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19885_ (.A0(_01075_),
    .A1(_02850_),
    .S(_02869_),
    .X(_01829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19886_ (.A0(_01007_),
    .A1(_02855_),
    .S(_02869_),
    .X(_01828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19887_ (.A0(_01819_),
    .A1(_03187_),
    .S(_02853_),
    .X(_01820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19888_ (.A0(_01820_),
    .A1(_02886_),
    .S(_03159_),
    .X(_01821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19889_ (.A0(_00841_),
    .A1(_01301_),
    .S(_02849_),
    .X(_01822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19890_ (.A0(_01823_),
    .A1(_02690_),
    .S(_00854_),
    .X(_01824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19891_ (.A0(_01824_),
    .A1(_01807_),
    .S(_02870_),
    .X(_01825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19892_ (.A0(_01825_),
    .A1(_01826_),
    .S(_00857_),
    .X(_01827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19893_ (.A0(_01487_),
    .A1(_02684_),
    .S(_03103_),
    .X(_01816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19894_ (.A0(_01815_),
    .A1(_01816_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_01817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19895_ (.A0(_02879_),
    .A1(_02888_),
    .S(_03135_),
    .X(_01810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19896_ (.A0(_01810_),
    .A1(_01769_),
    .S(_03128_),
    .X(_01811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19897_ (.A0(_01811_),
    .A1(_01729_),
    .S(_03120_),
    .X(_01812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19898_ (.A0(_01812_),
    .A1(_01648_),
    .S(_03111_),
    .X(_01813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19899_ (.A0(_01813_),
    .A1(_01483_),
    .S(_03103_),
    .X(_01814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19900_ (.A0(_01798_),
    .A1(_03186_),
    .S(_02853_),
    .X(_01799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19901_ (.A0(_01799_),
    .A1(_02895_),
    .S(_03159_),
    .X(_01800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19902_ (.A0(_00841_),
    .A1(_01255_),
    .S(_02849_),
    .X(_01801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19903_ (.A0(_01802_),
    .A1(_02696_),
    .S(_00854_),
    .X(_01803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19904_ (.A0(_01803_),
    .A1(_01787_),
    .S(_02870_),
    .X(_01804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19905_ (.A0(_01804_),
    .A1(_01805_),
    .S(_00857_),
    .X(_01806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19906_ (.A0(_01460_),
    .A1(_02684_),
    .S(_03103_),
    .X(_01795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19907_ (.A0(_01794_),
    .A1(_01795_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_01796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19908_ (.A0(_00786_),
    .A1(_00788_),
    .S(_03128_),
    .X(_01790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19909_ (.A0(_01790_),
    .A1(_01707_),
    .S(_03120_),
    .X(_01791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19910_ (.A0(_01791_),
    .A1(_01626_),
    .S(_03111_),
    .X(_01792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19911_ (.A0(_01792_),
    .A1(_01456_),
    .S(_03103_),
    .X(_01793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19912_ (.A0(_01778_),
    .A1(_03185_),
    .S(_02853_),
    .X(_01779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19913_ (.A0(_01779_),
    .A1(_02904_),
    .S(_03159_),
    .X(_01780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19914_ (.A0(_00841_),
    .A1(_01212_),
    .S(_02849_),
    .X(_01781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19915_ (.A0(_01782_),
    .A1(_02702_),
    .S(_00854_),
    .X(_01783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19916_ (.A0(_01783_),
    .A1(_01765_),
    .S(_02870_),
    .X(_01784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19917_ (.A0(_01784_),
    .A1(_01785_),
    .S(_00857_),
    .X(_01786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19918_ (.A0(_01438_),
    .A1(_02684_),
    .S(_03103_),
    .X(_01775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19919_ (.A0(_01774_),
    .A1(_01775_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_01776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19920_ (.A0(_01769_),
    .A1(_01728_),
    .S(_03128_),
    .X(_01770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19921_ (.A0(_01770_),
    .A1(_01687_),
    .S(_03120_),
    .X(_01771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19922_ (.A0(_01771_),
    .A1(_01606_),
    .S(_03111_),
    .X(_01772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19923_ (.A0(_01772_),
    .A1(_01434_),
    .S(_03103_),
    .X(_01773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19924_ (.A0(_02897_),
    .A1(_02905_),
    .S(_03135_),
    .X(_01769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19925_ (.A0(_01756_),
    .A1(_03184_),
    .S(_02853_),
    .X(_01757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19926_ (.A0(_01757_),
    .A1(_02912_),
    .S(_03159_),
    .X(_01758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19927_ (.A0(_00841_),
    .A1(_01168_),
    .S(_02849_),
    .X(_01759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19928_ (.A0(_01760_),
    .A1(_02708_),
    .S(_00854_),
    .X(_01761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19929_ (.A0(_01761_),
    .A1(_01746_),
    .S(_02870_),
    .X(_01762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19930_ (.A0(_01762_),
    .A1(_01763_),
    .S(_00857_),
    .X(_01764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19931_ (.A0(_01414_),
    .A1(_02684_),
    .S(_03103_),
    .X(_01753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19932_ (.A0(_01752_),
    .A1(_01753_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_01754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19933_ (.A0(_00790_),
    .A1(_00794_),
    .S(_03120_),
    .X(_01749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19934_ (.A0(_01749_),
    .A1(_01584_),
    .S(_03111_),
    .X(_01750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19935_ (.A0(_01750_),
    .A1(_01410_),
    .S(_03103_),
    .X(_01751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19936_ (.A0(_01737_),
    .A1(_03183_),
    .S(_02853_),
    .X(_01738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19937_ (.A0(_01738_),
    .A1(_02921_),
    .S(_03159_),
    .X(_01739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19938_ (.A0(_00841_),
    .A1(_01120_),
    .S(_02849_),
    .X(_01740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19939_ (.A0(_01741_),
    .A1(_02714_),
    .S(_00854_),
    .X(_01742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19940_ (.A0(_01742_),
    .A1(_01724_),
    .S(_02870_),
    .X(_01743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19941_ (.A0(_01743_),
    .A1(_01744_),
    .S(_00857_),
    .X(_01745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19942_ (.A0(_01393_),
    .A1(_02684_),
    .S(_03103_),
    .X(_01734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19943_ (.A0(_01733_),
    .A1(_01734_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_01735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19944_ (.A0(_01729_),
    .A1(_01647_),
    .S(_03120_),
    .X(_01730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19945_ (.A0(_01730_),
    .A1(_01565_),
    .S(_03111_),
    .X(_01731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19946_ (.A0(_01731_),
    .A1(_01389_),
    .S(_03103_),
    .X(_01732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19947_ (.A0(_01728_),
    .A1(_01686_),
    .S(_03128_),
    .X(_01729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19948_ (.A0(_02914_),
    .A1(_02922_),
    .S(_03135_),
    .X(_01728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19949_ (.A0(_01715_),
    .A1(_03182_),
    .S(_02853_),
    .X(_01716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19950_ (.A0(_01716_),
    .A1(_02929_),
    .S(_03159_),
    .X(_01717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19951_ (.A0(_00841_),
    .A1(_01065_),
    .S(_02849_),
    .X(_01718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19952_ (.A0(_01719_),
    .A1(_02720_),
    .S(_00854_),
    .X(_01720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19953_ (.A0(_01720_),
    .A1(_01704_),
    .S(_02870_),
    .X(_01721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19954_ (.A0(_01721_),
    .A1(_01722_),
    .S(_00857_),
    .X(_01723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19955_ (.A0(_01369_),
    .A1(_02684_),
    .S(_03103_),
    .X(_01712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19956_ (.A0(_01711_),
    .A1(_01712_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_01713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19957_ (.A0(_01707_),
    .A1(_01625_),
    .S(_03120_),
    .X(_01708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19958_ (.A0(_01708_),
    .A1(_01542_),
    .S(_03111_),
    .X(_01709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19959_ (.A0(_01709_),
    .A1(_01365_),
    .S(_03103_),
    .X(_01710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19960_ (.A0(_00789_),
    .A1(_00792_),
    .S(_03128_),
    .X(_01707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19961_ (.A0(_01695_),
    .A1(_03181_),
    .S(_02853_),
    .X(_01696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19962_ (.A0(_01696_),
    .A1(_02938_),
    .S(_03159_),
    .X(_01697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19963_ (.A0(_00841_),
    .A1(_00997_),
    .S(_02849_),
    .X(_01698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19964_ (.A0(_01699_),
    .A1(_02726_),
    .S(_00854_),
    .X(_01700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19965_ (.A0(_01700_),
    .A1(_01682_),
    .S(_02870_),
    .X(_01701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19966_ (.A0(_01701_),
    .A1(_01702_),
    .S(_00857_),
    .X(_01703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19967_ (.A0(_01347_),
    .A1(_02684_),
    .S(_03103_),
    .X(_01692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19968_ (.A0(_01691_),
    .A1(_01692_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_01693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19969_ (.A0(_01687_),
    .A1(_01605_),
    .S(_03120_),
    .X(_01688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19970_ (.A0(_01688_),
    .A1(_01522_),
    .S(_03111_),
    .X(_01689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19971_ (.A0(_01689_),
    .A1(_01343_),
    .S(_03103_),
    .X(_01690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19972_ (.A0(_01686_),
    .A1(_01646_),
    .S(_03128_),
    .X(_01687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19973_ (.A0(_02931_),
    .A1(_02939_),
    .S(_03135_),
    .X(_01686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19974_ (.A0(_01673_),
    .A1(_03180_),
    .S(_02853_),
    .X(_01674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19975_ (.A0(_01674_),
    .A1(_02946_),
    .S(_03159_),
    .X(_01675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19976_ (.A0(_00841_),
    .A1(_00845_),
    .S(_02849_),
    .X(_01676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19977_ (.A0(_01677_),
    .A1(_02732_),
    .S(_00854_),
    .X(_01678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19978_ (.A0(_01678_),
    .A1(_01664_),
    .S(_02870_),
    .X(_01679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19979_ (.A0(_01679_),
    .A1(_01680_),
    .S(_00857_),
    .X(_01681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19980_ (.A0(_01323_),
    .A1(_02684_),
    .S(_03103_),
    .X(_01670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19981_ (.A0(_01669_),
    .A1(_01670_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_01671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19982_ (.A0(_00798_),
    .A1(_00808_),
    .S(_03111_),
    .X(_01667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19983_ (.A0(_01667_),
    .A1(_01316_),
    .S(_03103_),
    .X(_01668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19984_ (.A0(_01655_),
    .A1(_03179_),
    .S(_02853_),
    .X(_01656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19985_ (.A0(_01656_),
    .A1(_02955_),
    .S(_03159_),
    .X(_01657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19986_ (.A0(_00841_),
    .A1(_01296_),
    .S(_02849_),
    .X(_01658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19987_ (.A0(_01659_),
    .A1(_02738_),
    .S(_00854_),
    .X(_01660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19988_ (.A0(_01660_),
    .A1(_01642_),
    .S(_02870_),
    .X(_01661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19989_ (.A0(_01661_),
    .A1(_01662_),
    .S(_00857_),
    .X(_01663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19990_ (.A0(_01284_),
    .A1(_02684_),
    .S(_03103_),
    .X(_01652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19991_ (.A0(_01651_),
    .A1(_01652_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_01653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19992_ (.A0(_01648_),
    .A1(_01482_),
    .S(_03111_),
    .X(_01649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19993_ (.A0(_01649_),
    .A1(_01275_),
    .S(_03103_),
    .X(_01650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19994_ (.A0(_01647_),
    .A1(_01564_),
    .S(_03120_),
    .X(_01648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19995_ (.A0(_01646_),
    .A1(_01604_),
    .S(_03128_),
    .X(_01647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19996_ (.A0(_02948_),
    .A1(_02956_),
    .S(_03135_),
    .X(_01646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19997_ (.A0(_01633_),
    .A1(_03178_),
    .S(_02853_),
    .X(_01634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19998_ (.A0(_01634_),
    .A1(_02963_),
    .S(_03159_),
    .X(_01635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _19999_ (.A0(_00841_),
    .A1(_01250_),
    .S(_02849_),
    .X(_01636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20000_ (.A0(_01637_),
    .A1(_02744_),
    .S(_00854_),
    .X(_01638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20001_ (.A0(_01638_),
    .A1(_01622_),
    .S(_02870_),
    .X(_01639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20002_ (.A0(_01639_),
    .A1(_01640_),
    .S(_00857_),
    .X(_01641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20003_ (.A0(_01238_),
    .A1(_02684_),
    .S(_03103_),
    .X(_01630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20004_ (.A0(_01629_),
    .A1(_01630_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_01631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20005_ (.A0(_01626_),
    .A1(_01455_),
    .S(_03111_),
    .X(_01627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20006_ (.A0(_01627_),
    .A1(_01229_),
    .S(_03103_),
    .X(_01628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20007_ (.A0(_01625_),
    .A1(_01541_),
    .S(_03120_),
    .X(_01626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20008_ (.A0(_00793_),
    .A1(_00795_),
    .S(_03128_),
    .X(_01625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20009_ (.A0(_01613_),
    .A1(_03177_),
    .S(_02853_),
    .X(_01614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20010_ (.A0(_01614_),
    .A1(_02972_),
    .S(_03159_),
    .X(_01615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20011_ (.A0(_00841_),
    .A1(_01207_),
    .S(_02849_),
    .X(_01616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20012_ (.A0(_01617_),
    .A1(_02750_),
    .S(_00854_),
    .X(_01618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20013_ (.A0(_01618_),
    .A1(_01600_),
    .S(_02870_),
    .X(_01619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20014_ (.A0(_01619_),
    .A1(_01620_),
    .S(_00857_),
    .X(_01621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20015_ (.A0(_01196_),
    .A1(_02684_),
    .S(_03103_),
    .X(_01610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20016_ (.A0(_01609_),
    .A1(_01610_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_01611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20017_ (.A0(_01606_),
    .A1(_01433_),
    .S(_03111_),
    .X(_01607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20018_ (.A0(_01607_),
    .A1(_01187_),
    .S(_03103_),
    .X(_01608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20019_ (.A0(_01605_),
    .A1(_01521_),
    .S(_03120_),
    .X(_01606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20020_ (.A0(_01604_),
    .A1(_01563_),
    .S(_03128_),
    .X(_01605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20021_ (.A0(_02965_),
    .A1(_02973_),
    .S(_03135_),
    .X(_01604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20022_ (.A0(_01591_),
    .A1(_03176_),
    .S(_02853_),
    .X(_01592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20023_ (.A0(_01592_),
    .A1(_02980_),
    .S(_03159_),
    .X(_01593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20024_ (.A0(_00841_),
    .A1(_01163_),
    .S(_02849_),
    .X(_01594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20025_ (.A0(_01595_),
    .A1(_02756_),
    .S(_00854_),
    .X(_01596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20026_ (.A0(_01596_),
    .A1(_01581_),
    .S(_02870_),
    .X(_01597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20027_ (.A0(_01597_),
    .A1(_01598_),
    .S(_00857_),
    .X(_01599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20028_ (.A0(_01152_),
    .A1(_02684_),
    .S(_03103_),
    .X(_01588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20029_ (.A0(_01587_),
    .A1(_01588_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_01589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20030_ (.A0(_01584_),
    .A1(_01409_),
    .S(_03111_),
    .X(_01585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20031_ (.A0(_01585_),
    .A1(_01136_),
    .S(_03103_),
    .X(_01586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20032_ (.A0(_00797_),
    .A1(_00802_),
    .S(_03120_),
    .X(_01584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20033_ (.A0(_01572_),
    .A1(_01560_),
    .S(_02853_),
    .X(_01573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20034_ (.A0(_01573_),
    .A1(_02989_),
    .S(_03159_),
    .X(_01574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20035_ (.A0(_00841_),
    .A1(_01115_),
    .S(_02849_),
    .X(_01575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20036_ (.A0(_01576_),
    .A1(_02762_),
    .S(_00854_),
    .X(_01577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20037_ (.A0(_01577_),
    .A1(_01558_),
    .S(_02870_),
    .X(_01578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20038_ (.A0(_01578_),
    .A1(_01579_),
    .S(_00857_),
    .X(_01580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20039_ (.A0(_01103_),
    .A1(_02684_),
    .S(_03103_),
    .X(_01569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20040_ (.A0(_01568_),
    .A1(_01569_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_01570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20041_ (.A0(_01565_),
    .A1(_01388_),
    .S(_03111_),
    .X(_01566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20042_ (.A0(_01566_),
    .A1(_01085_),
    .S(_03103_),
    .X(_01567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20043_ (.A0(_01564_),
    .A1(_01481_),
    .S(_03120_),
    .X(_01565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20044_ (.A0(_01563_),
    .A1(_01520_),
    .S(_03128_),
    .X(_01564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20045_ (.A0(_02982_),
    .A1(_02990_),
    .S(_03135_),
    .X(_01563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20046_ (.A0(_01549_),
    .A1(_03175_),
    .S(_02853_),
    .X(_01550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20047_ (.A0(_01550_),
    .A1(_02997_),
    .S(_03159_),
    .X(_01551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20048_ (.A0(_00841_),
    .A1(_01059_),
    .S(_02849_),
    .X(_01552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20049_ (.A0(_01553_),
    .A1(_02768_),
    .S(_00854_),
    .X(_01554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20050_ (.A0(_01554_),
    .A1(_01538_),
    .S(_02870_),
    .X(_01555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20051_ (.A0(_01555_),
    .A1(_01556_),
    .S(_00857_),
    .X(_01557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20052_ (.A0(_01048_),
    .A1(_02684_),
    .S(_03103_),
    .X(_01546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20053_ (.A0(_01545_),
    .A1(_01546_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_01547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20054_ (.A0(_01542_),
    .A1(_01364_),
    .S(_03111_),
    .X(_01543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20055_ (.A0(_01543_),
    .A1(_01015_),
    .S(_03103_),
    .X(_01544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20056_ (.A0(_01541_),
    .A1(_01454_),
    .S(_03120_),
    .X(_01542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20057_ (.A0(_00796_),
    .A1(_00800_),
    .S(_03128_),
    .X(_01541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20058_ (.A0(_01529_),
    .A1(_03174_),
    .S(_02853_),
    .X(_01530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20059_ (.A0(_01530_),
    .A1(_03006_),
    .S(_03159_),
    .X(_01531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20060_ (.A0(_00841_),
    .A1(_00990_),
    .S(_02849_),
    .X(_01532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20061_ (.A0(_01533_),
    .A1(_02774_),
    .S(_00854_),
    .X(_01534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20062_ (.A0(_01534_),
    .A1(_01516_),
    .S(_02870_),
    .X(_01535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20063_ (.A0(_01535_),
    .A1(_01536_),
    .S(_00857_),
    .X(_01537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20064_ (.A0(_00975_),
    .A1(_02684_),
    .S(_03103_),
    .X(_01526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20065_ (.A0(_01525_),
    .A1(_01526_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_01527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20066_ (.A0(_01522_),
    .A1(_01342_),
    .S(_03111_),
    .X(_01523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20067_ (.A0(_01523_),
    .A1(_00944_),
    .S(_03103_),
    .X(_01524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20068_ (.A0(_01521_),
    .A1(_01432_),
    .S(_03120_),
    .X(_01522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20069_ (.A0(_01520_),
    .A1(_01480_),
    .S(_03128_),
    .X(_01521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20070_ (.A0(_02999_),
    .A1(_03007_),
    .S(_03135_),
    .X(_01520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20071_ (.A0(_01507_),
    .A1(_03173_),
    .S(_02853_),
    .X(_01508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20072_ (.A0(_01508_),
    .A1(_03014_),
    .S(_03159_),
    .X(_01509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20073_ (.A0(_00840_),
    .A1(_00839_),
    .S(_02849_),
    .X(_01510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20074_ (.A0(_01511_),
    .A1(_02780_),
    .S(_00854_),
    .X(_01512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20075_ (.A0(_01512_),
    .A1(_01500_),
    .S(_02870_),
    .X(_01513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20076_ (.A0(_01513_),
    .A1(_01514_),
    .S(_00857_),
    .X(_01515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20077_ (.A0(_01319_),
    .A1(_01321_),
    .S(_03111_),
    .X(_01504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20078_ (.A0(_01490_),
    .A1(_01477_),
    .S(_02853_),
    .X(_01491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20079_ (.A0(_01491_),
    .A1(_03023_),
    .S(_03159_),
    .X(_01492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20080_ (.A0(_01301_),
    .A1(_01304_),
    .S(_02850_),
    .X(_01493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20081_ (.A0(_01493_),
    .A1(_01304_),
    .S(_02849_),
    .X(_01494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20082_ (.A0(_01495_),
    .A1(_02786_),
    .S(_00854_),
    .X(_01496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20083_ (.A0(_01496_),
    .A1(_01475_),
    .S(_02870_),
    .X(_01497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20084_ (.A0(_01497_),
    .A1(_01498_),
    .S(_00857_),
    .X(_01499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20085_ (.A0(_01283_),
    .A1(_02684_),
    .S(_03111_),
    .X(_01487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20086_ (.A0(_01278_),
    .A1(_01280_),
    .S(_03111_),
    .X(_01485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20087_ (.A0(_01482_),
    .A1(_01274_),
    .S(_03111_),
    .X(_01483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20088_ (.A0(_01481_),
    .A1(_01387_),
    .S(_03120_),
    .X(_01482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20089_ (.A0(_01480_),
    .A1(_01431_),
    .S(_03128_),
    .X(_01481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20090_ (.A0(_03016_),
    .A1(_03024_),
    .S(_03135_),
    .X(_01480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20091_ (.A0(_01463_),
    .A1(_03172_),
    .S(_02853_),
    .X(_01464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20092_ (.A0(_01464_),
    .A1(_03031_),
    .S(_03159_),
    .X(_01465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20093_ (.A0(_01255_),
    .A1(_01258_),
    .S(_02850_),
    .X(_01466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20094_ (.A0(_01466_),
    .A1(_01258_),
    .S(_02849_),
    .X(_01467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20095_ (.A0(_01468_),
    .A1(_02792_),
    .S(_00854_),
    .X(_01469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20096_ (.A0(_01469_),
    .A1(_01451_),
    .S(_02870_),
    .X(_01470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20097_ (.A0(_01470_),
    .A1(_01471_),
    .S(_00857_),
    .X(_01472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20098_ (.A0(_01237_),
    .A1(_02684_),
    .S(_03111_),
    .X(_01460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20099_ (.A0(_01232_),
    .A1(_01234_),
    .S(_03111_),
    .X(_01458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20100_ (.A0(_01455_),
    .A1(_01228_),
    .S(_03111_),
    .X(_01456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20101_ (.A0(_01454_),
    .A1(_01363_),
    .S(_03120_),
    .X(_01455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20102_ (.A0(_00801_),
    .A1(_00804_),
    .S(_03128_),
    .X(_01454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20103_ (.A0(_01441_),
    .A1(_03171_),
    .S(_02853_),
    .X(_01442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20104_ (.A0(_01442_),
    .A1(_03040_),
    .S(_03159_),
    .X(_01443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20105_ (.A0(_01212_),
    .A1(_01215_),
    .S(_02850_),
    .X(_01444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20106_ (.A0(_01444_),
    .A1(_01215_),
    .S(_02849_),
    .X(_01445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20107_ (.A0(_01446_),
    .A1(_02798_),
    .S(_00854_),
    .X(_01447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20108_ (.A0(_01447_),
    .A1(_01427_),
    .S(_02870_),
    .X(_01448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20109_ (.A0(_01448_),
    .A1(_01449_),
    .S(_00857_),
    .X(_01450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20110_ (.A0(_01195_),
    .A1(_02684_),
    .S(_03111_),
    .X(_01438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20111_ (.A0(_01190_),
    .A1(_01192_),
    .S(_03111_),
    .X(_01436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20112_ (.A0(_01433_),
    .A1(_01186_),
    .S(_03111_),
    .X(_01434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20113_ (.A0(_01432_),
    .A1(_01341_),
    .S(_03120_),
    .X(_01433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20114_ (.A0(_01431_),
    .A1(_01386_),
    .S(_03128_),
    .X(_01432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20115_ (.A0(_03033_),
    .A1(_00803_),
    .S(_03135_),
    .X(_01431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20116_ (.A0(_01417_),
    .A1(_03170_),
    .S(_02853_),
    .X(_01418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20117_ (.A0(_01418_),
    .A1(_03047_),
    .S(_03159_),
    .X(_01419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20118_ (.A0(_01168_),
    .A1(_01171_),
    .S(_02850_),
    .X(_01420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20119_ (.A0(_01420_),
    .A1(_01171_),
    .S(_02849_),
    .X(_01421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20120_ (.A0(_01422_),
    .A1(_02804_),
    .S(_00854_),
    .X(_01423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20121_ (.A0(_01423_),
    .A1(_01406_),
    .S(_02870_),
    .X(_01424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20122_ (.A0(_01424_),
    .A1(_01425_),
    .S(_00857_),
    .X(_01426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20123_ (.A0(_01151_),
    .A1(_02684_),
    .S(_03111_),
    .X(_01414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20124_ (.A0(_01143_),
    .A1(_01147_),
    .S(_03111_),
    .X(_01412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20125_ (.A0(_01409_),
    .A1(_01135_),
    .S(_03111_),
    .X(_01410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20126_ (.A0(_00807_),
    .A1(_00813_),
    .S(_03120_),
    .X(_01409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20127_ (.A0(_01396_),
    .A1(_03169_),
    .S(_02853_),
    .X(_01397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20128_ (.A0(_01397_),
    .A1(_03056_),
    .S(_03159_),
    .X(_01398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20129_ (.A0(_01120_),
    .A1(_01123_),
    .S(_02850_),
    .X(_01399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20130_ (.A0(_01399_),
    .A1(_01123_),
    .S(_02849_),
    .X(_01400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20131_ (.A0(_01401_),
    .A1(_02810_),
    .S(_00854_),
    .X(_01402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20132_ (.A0(_01402_),
    .A1(_01382_),
    .S(_02870_),
    .X(_01403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20133_ (.A0(_01403_),
    .A1(_01404_),
    .S(_00857_),
    .X(_01405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20134_ (.A0(_01102_),
    .A1(_02684_),
    .S(_03111_),
    .X(_01393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20135_ (.A0(_01092_),
    .A1(_01096_),
    .S(_03111_),
    .X(_01391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20136_ (.A0(_01388_),
    .A1(_01084_),
    .S(_03111_),
    .X(_01389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20137_ (.A0(_01387_),
    .A1(_01273_),
    .S(_03120_),
    .X(_01388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20138_ (.A0(_01386_),
    .A1(_01340_),
    .S(_03128_),
    .X(_01387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20139_ (.A0(_03049_),
    .A1(_00805_),
    .S(_03135_),
    .X(_01386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20140_ (.A0(_01372_),
    .A1(_03168_),
    .S(_02853_),
    .X(_01373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20141_ (.A0(_01373_),
    .A1(_03063_),
    .S(_03159_),
    .X(_01374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20142_ (.A0(_01065_),
    .A1(_01068_),
    .S(_02850_),
    .X(_01375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20143_ (.A0(_01375_),
    .A1(_01068_),
    .S(_02849_),
    .X(_01376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20144_ (.A0(_01377_),
    .A1(_02816_),
    .S(_00854_),
    .X(_01378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20145_ (.A0(_01378_),
    .A1(_01360_),
    .S(_02870_),
    .X(_01379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20146_ (.A0(_01379_),
    .A1(_01380_),
    .S(_00857_),
    .X(_01381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20147_ (.A0(_01047_),
    .A1(_02684_),
    .S(_03111_),
    .X(_01369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20148_ (.A0(_01030_),
    .A1(_01038_),
    .S(_03111_),
    .X(_01367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20149_ (.A0(_01364_),
    .A1(_01014_),
    .S(_03111_),
    .X(_01365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20150_ (.A0(_01363_),
    .A1(_01227_),
    .S(_03120_),
    .X(_01364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20151_ (.A0(_00806_),
    .A1(_00810_),
    .S(_03128_),
    .X(_01363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20152_ (.A0(_01350_),
    .A1(_03167_),
    .S(_02853_),
    .X(_01351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20153_ (.A0(_01351_),
    .A1(_03072_),
    .S(_03159_),
    .X(_01352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20154_ (.A0(_00997_),
    .A1(_01000_),
    .S(_02850_),
    .X(_01353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20155_ (.A0(_01353_),
    .A1(_01000_),
    .S(_02849_),
    .X(_01354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20156_ (.A0(_01355_),
    .A1(_02822_),
    .S(_00854_),
    .X(_01356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20157_ (.A0(_01356_),
    .A1(_01336_),
    .S(_02870_),
    .X(_01357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20158_ (.A0(_01357_),
    .A1(_01358_),
    .S(_00857_),
    .X(_01359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20159_ (.A0(_00974_),
    .A1(_02684_),
    .S(_03111_),
    .X(_01347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20160_ (.A0(_00959_),
    .A1(_00967_),
    .S(_03111_),
    .X(_01345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20161_ (.A0(_01342_),
    .A1(_00943_),
    .S(_03111_),
    .X(_01343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20162_ (.A0(_01341_),
    .A1(_01185_),
    .S(_03120_),
    .X(_01342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20163_ (.A0(_01340_),
    .A1(_01272_),
    .S(_03128_),
    .X(_01341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20164_ (.A0(_03065_),
    .A1(_00809_),
    .S(_03135_),
    .X(_01340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20165_ (.A0(_01326_),
    .A1(_03166_),
    .S(_02853_),
    .X(_01327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20166_ (.A0(_01327_),
    .A1(_03079_),
    .S(_03159_),
    .X(_01328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20167_ (.A0(_00845_),
    .A1(_00848_),
    .S(_02850_),
    .X(_01329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20168_ (.A0(_01329_),
    .A1(_00848_),
    .S(_02849_),
    .X(_01330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20169_ (.A0(_01331_),
    .A1(_02828_),
    .S(_00854_),
    .X(_01332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20170_ (.A0(_01332_),
    .A1(_01313_),
    .S(_02870_),
    .X(_01333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20171_ (.A0(_01333_),
    .A1(_01334_),
    .S(_00857_),
    .X(_01335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20172_ (.A0(_01321_),
    .A1(_02684_),
    .S(_03111_),
    .X(_01323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20173_ (.A0(_01321_),
    .A1(_00822_),
    .S(_03111_),
    .X(_01322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20174_ (.A0(_01146_),
    .A1(_01148_),
    .S(_03120_),
    .X(_01321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20175_ (.A0(_01139_),
    .A1(_01141_),
    .S(_03120_),
    .X(_01318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20176_ (.A0(_01318_),
    .A1(_01319_),
    .S(_03111_),
    .X(_01320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20177_ (.A0(_01142_),
    .A1(_01145_),
    .S(_03120_),
    .X(_01319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20178_ (.A0(_01287_),
    .A1(_01269_),
    .S(_02853_),
    .X(_01288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20179_ (.A0(_01288_),
    .A1(_03088_),
    .S(_03159_),
    .X(_01289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20180_ (.A0(_01292_),
    .A1(_01304_),
    .S(_00754_),
    .X(_01305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20181_ (.A0(_01305_),
    .A1(_01296_),
    .S(_03273_),
    .X(_01306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20182_ (.A0(_01306_),
    .A1(_01301_),
    .S(_02866_),
    .X(_01307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20183_ (.A0(_01296_),
    .A1(_01292_),
    .S(_02850_),
    .X(_01297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20184_ (.A0(_01297_),
    .A1(_01292_),
    .S(_02849_),
    .X(_01298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20185_ (.A0(_01308_),
    .A1(_02834_),
    .S(_00854_),
    .X(_01309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20186_ (.A0(_01309_),
    .A1(_01267_),
    .S(_02870_),
    .X(_01310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20187_ (.A0(_01310_),
    .A1(_01311_),
    .S(_00857_),
    .X(_01312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20188_ (.A0(_01302_),
    .A1(_01303_),
    .S(\design_top.XADDR[31] ),
    .X(_01304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20189_ (.A0(_01299_),
    .A1(_01300_),
    .S(\design_top.XADDR[31] ),
    .X(_01301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20190_ (.A0(_00994_),
    .A1(_01294_),
    .S(\design_top.XADDR[3] ),
    .X(_01295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20191_ (.A0(_01293_),
    .A1(_01295_),
    .S(\design_top.XADDR[31] ),
    .X(_01296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20192_ (.A0(_01290_),
    .A1(_01291_),
    .S(\design_top.XADDR[31] ),
    .X(_01292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20193_ (.A0(_01280_),
    .A1(_01283_),
    .S(_03111_),
    .X(_01284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20194_ (.A0(_01101_),
    .A1(_02684_),
    .S(_03120_),
    .X(_01283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20195_ (.A0(_01280_),
    .A1(_01281_),
    .S(_03111_),
    .X(_01282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20196_ (.A0(_01095_),
    .A1(_01097_),
    .S(_03120_),
    .X(_01280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20197_ (.A0(_01088_),
    .A1(_01090_),
    .S(_03120_),
    .X(_01277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20198_ (.A0(_01277_),
    .A1(_01278_),
    .S(_03111_),
    .X(_01279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20199_ (.A0(_01091_),
    .A1(_01094_),
    .S(_03120_),
    .X(_01278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20200_ (.A0(_01273_),
    .A1(_01083_),
    .S(_03120_),
    .X(_01274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20201_ (.A0(_01272_),
    .A1(_01184_),
    .S(_03128_),
    .X(_01273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20202_ (.A0(_03081_),
    .A1(_00811_),
    .S(_03135_),
    .X(_01272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20203_ (.A0(_01241_),
    .A1(_03165_),
    .S(_02853_),
    .X(_01242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20204_ (.A0(_01242_),
    .A1(_03095_),
    .S(_03159_),
    .X(_01243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20205_ (.A0(_01246_),
    .A1(_01258_),
    .S(_00754_),
    .X(_01259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20206_ (.A0(_01259_),
    .A1(_01250_),
    .S(_03273_),
    .X(_01260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20207_ (.A0(_01260_),
    .A1(_01255_),
    .S(_02866_),
    .X(_01261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20208_ (.A0(_01250_),
    .A1(_01246_),
    .S(_02850_),
    .X(_01251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20209_ (.A0(_01251_),
    .A1(_01246_),
    .S(_02849_),
    .X(_01252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20210_ (.A0(_01262_),
    .A1(_02840_),
    .S(_00854_),
    .X(_01263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20211_ (.A0(_01263_),
    .A1(_01224_),
    .S(_02870_),
    .X(_01264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20212_ (.A0(_01264_),
    .A1(_01265_),
    .S(_00857_),
    .X(_01266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20213_ (.A0(_01256_),
    .A1(_01257_),
    .S(\design_top.XADDR[31] ),
    .X(_01258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20214_ (.A0(_01253_),
    .A1(_01254_),
    .S(\design_top.XADDR[31] ),
    .X(_01255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20215_ (.A0(_00994_),
    .A1(_01248_),
    .S(\design_top.XADDR[3] ),
    .X(_01249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20216_ (.A0(_01247_),
    .A1(_01249_),
    .S(\design_top.XADDR[31] ),
    .X(_01250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20217_ (.A0(_01244_),
    .A1(_01245_),
    .S(\design_top.XADDR[31] ),
    .X(_01246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20218_ (.A0(_01234_),
    .A1(_01237_),
    .S(_03111_),
    .X(_01238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20219_ (.A0(_01046_),
    .A1(_02684_),
    .S(_03120_),
    .X(_01237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20220_ (.A0(_01234_),
    .A1(_01235_),
    .S(_03111_),
    .X(_01236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20221_ (.A0(_01037_),
    .A1(_01041_),
    .S(_03120_),
    .X(_01234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20222_ (.A0(_01022_),
    .A1(_01026_),
    .S(_03120_),
    .X(_01231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20223_ (.A0(_01231_),
    .A1(_01232_),
    .S(_03111_),
    .X(_01233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20224_ (.A0(_01029_),
    .A1(_01034_),
    .S(_03120_),
    .X(_01232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20225_ (.A0(_01227_),
    .A1(_01013_),
    .S(_03120_),
    .X(_01228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20226_ (.A0(_00812_),
    .A1(_00814_),
    .S(_03128_),
    .X(_01227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20227_ (.A0(_01199_),
    .A1(_03164_),
    .S(_02853_),
    .X(_01200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20228_ (.A0(_01200_),
    .A1(_03104_),
    .S(_03159_),
    .X(_01201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20229_ (.A0(_01204_),
    .A1(_01215_),
    .S(_00754_),
    .X(_01216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20230_ (.A0(_01216_),
    .A1(_01207_),
    .S(_03273_),
    .X(_01217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20231_ (.A0(_01217_),
    .A1(_01212_),
    .S(_02866_),
    .X(_01218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20232_ (.A0(_01207_),
    .A1(_01204_),
    .S(_02850_),
    .X(_01208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20233_ (.A0(_01208_),
    .A1(_01204_),
    .S(_02849_),
    .X(_01209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20234_ (.A0(_01219_),
    .A1(_02846_),
    .S(_00854_),
    .X(_01220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20235_ (.A0(_01220_),
    .A1(_01180_),
    .S(_02870_),
    .X(_01221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20236_ (.A0(_01221_),
    .A1(_01222_),
    .S(_00857_),
    .X(_01223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20237_ (.A0(_01213_),
    .A1(_01214_),
    .S(\design_top.XADDR[31] ),
    .X(_01215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20238_ (.A0(_01210_),
    .A1(_01211_),
    .S(\design_top.XADDR[31] ),
    .X(_01212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20239_ (.A0(_01205_),
    .A1(_01206_),
    .S(\design_top.XADDR[31] ),
    .X(_01207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20240_ (.A0(_01202_),
    .A1(_01203_),
    .S(\design_top.XADDR[31] ),
    .X(_01204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20241_ (.A0(_01192_),
    .A1(_01195_),
    .S(_03111_),
    .X(_01196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20242_ (.A0(_00973_),
    .A1(_02684_),
    .S(_03120_),
    .X(_01195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20243_ (.A0(_01192_),
    .A1(_01193_),
    .S(_03111_),
    .X(_01194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20244_ (.A0(_00966_),
    .A1(_00970_),
    .S(_03120_),
    .X(_01192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20245_ (.A0(_00951_),
    .A1(_00955_),
    .S(_03120_),
    .X(_01189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20246_ (.A0(_01189_),
    .A1(_01190_),
    .S(_03111_),
    .X(_01191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20247_ (.A0(_00958_),
    .A1(_00963_),
    .S(_03120_),
    .X(_01190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20248_ (.A0(_01185_),
    .A1(_00942_),
    .S(_03120_),
    .X(_01186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20249_ (.A0(_01184_),
    .A1(_01082_),
    .S(_03128_),
    .X(_01185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20250_ (.A0(_03097_),
    .A1(_03105_),
    .S(_03135_),
    .X(_01184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20251_ (.A0(_01155_),
    .A1(_03163_),
    .S(_02853_),
    .X(_01156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20252_ (.A0(_01156_),
    .A1(_03112_),
    .S(_03159_),
    .X(_01157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20253_ (.A0(_01160_),
    .A1(_01171_),
    .S(_00754_),
    .X(_01172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20254_ (.A0(_01172_),
    .A1(_01163_),
    .S(_03273_),
    .X(_01173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20255_ (.A0(_01173_),
    .A1(_01168_),
    .S(_02866_),
    .X(_01174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20256_ (.A0(_01163_),
    .A1(_01160_),
    .S(_02850_),
    .X(_01164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20257_ (.A0(_01164_),
    .A1(_01160_),
    .S(_02849_),
    .X(_01165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20258_ (.A0(_01175_),
    .A1(_02652_),
    .S(_00854_),
    .X(_01176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20259_ (.A0(_01176_),
    .A1(_01132_),
    .S(_02870_),
    .X(_01177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20260_ (.A0(_01177_),
    .A1(_01178_),
    .S(_00857_),
    .X(_01179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20261_ (.A0(_01169_),
    .A1(_01170_),
    .S(\design_top.XADDR[31] ),
    .X(_01171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20262_ (.A0(_01166_),
    .A1(_01167_),
    .S(\design_top.XADDR[31] ),
    .X(_01168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20263_ (.A0(_01161_),
    .A1(_01162_),
    .S(\design_top.XADDR[31] ),
    .X(_01163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20264_ (.A0(_01158_),
    .A1(_01159_),
    .S(\design_top.XADDR[31] ),
    .X(_01160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20265_ (.A0(_01147_),
    .A1(_01151_),
    .S(_03111_),
    .X(_01152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20266_ (.A0(_01148_),
    .A1(_02684_),
    .S(_03120_),
    .X(_01151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20267_ (.A0(_01147_),
    .A1(_01149_),
    .S(_03111_),
    .X(_01150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20268_ (.A0(_01148_),
    .A1(_00821_),
    .S(_03120_),
    .X(_01149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20269_ (.A0(_01040_),
    .A1(_01042_),
    .S(_03128_),
    .X(_01148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20270_ (.A0(_01145_),
    .A1(_01146_),
    .S(_03120_),
    .X(_01147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20271_ (.A0(_01036_),
    .A1(_01039_),
    .S(_03128_),
    .X(_01146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20272_ (.A0(_01033_),
    .A1(_01035_),
    .S(_03128_),
    .X(_01145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20273_ (.A0(_01018_),
    .A1(_01020_),
    .S(_03128_),
    .X(_01138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20274_ (.A0(_01138_),
    .A1(_01139_),
    .S(_03120_),
    .X(_01140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20275_ (.A0(_01140_),
    .A1(_01143_),
    .S(_03111_),
    .X(_01144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20276_ (.A0(_01141_),
    .A1(_01142_),
    .S(_03120_),
    .X(_01143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20277_ (.A0(_01028_),
    .A1(_01032_),
    .S(_03128_),
    .X(_01142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20278_ (.A0(_01025_),
    .A1(_01027_),
    .S(_03128_),
    .X(_01141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20279_ (.A0(_01021_),
    .A1(_01024_),
    .S(_03128_),
    .X(_01139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20280_ (.A0(_01106_),
    .A1(_01079_),
    .S(_02853_),
    .X(_01107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20281_ (.A0(_01107_),
    .A1(_03121_),
    .S(_03159_),
    .X(_01108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20282_ (.A0(_01111_),
    .A1(_01123_),
    .S(_00754_),
    .X(_01124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20283_ (.A0(_01124_),
    .A1(_01115_),
    .S(_03273_),
    .X(_01125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20284_ (.A0(_01125_),
    .A1(_01120_),
    .S(_02866_),
    .X(_01126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20285_ (.A0(_01115_),
    .A1(_01111_),
    .S(_02850_),
    .X(_01116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20286_ (.A0(_01116_),
    .A1(_01111_),
    .S(_02849_),
    .X(_01117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20287_ (.A0(_01127_),
    .A1(_02627_),
    .S(_00854_),
    .X(_01128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20288_ (.A0(_01128_),
    .A1(_01077_),
    .S(_02870_),
    .X(_01129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20289_ (.A0(_01129_),
    .A1(_01130_),
    .S(_00857_),
    .X(_01131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20290_ (.A0(_01121_),
    .A1(_01122_),
    .S(\design_top.XADDR[31] ),
    .X(_01123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20291_ (.A0(_01118_),
    .A1(_01119_),
    .S(\design_top.XADDR[31] ),
    .X(_01120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20292_ (.A0(_00994_),
    .A1(_01113_),
    .S(\design_top.XADDR[3] ),
    .X(_01114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20293_ (.A0(_01112_),
    .A1(_01114_),
    .S(\design_top.XADDR[31] ),
    .X(_01115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20294_ (.A0(_01109_),
    .A1(_01110_),
    .S(\design_top.XADDR[31] ),
    .X(_01111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20295_ (.A0(_01096_),
    .A1(_01102_),
    .S(_03111_),
    .X(_01103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20296_ (.A0(_01097_),
    .A1(_01101_),
    .S(_03120_),
    .X(_01102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20297_ (.A0(_00972_),
    .A1(_02684_),
    .S(_03128_),
    .X(_01101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20298_ (.A0(_01096_),
    .A1(_01099_),
    .S(_03111_),
    .X(_01100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20299_ (.A0(_01097_),
    .A1(_01098_),
    .S(_03120_),
    .X(_01099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20300_ (.A0(_00969_),
    .A1(_00971_),
    .S(_03128_),
    .X(_01097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20301_ (.A0(_01094_),
    .A1(_01095_),
    .S(_03120_),
    .X(_01096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20302_ (.A0(_00965_),
    .A1(_00968_),
    .S(_03128_),
    .X(_01095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20303_ (.A0(_00962_),
    .A1(_00964_),
    .S(_03128_),
    .X(_01094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20304_ (.A0(_00947_),
    .A1(_00949_),
    .S(_03128_),
    .X(_01087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20305_ (.A0(_01087_),
    .A1(_01088_),
    .S(_03120_),
    .X(_01089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20306_ (.A0(_01089_),
    .A1(_01092_),
    .S(_03111_),
    .X(_01093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20307_ (.A0(_01090_),
    .A1(_01091_),
    .S(_03120_),
    .X(_01092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20308_ (.A0(_00957_),
    .A1(_00961_),
    .S(_03128_),
    .X(_01091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20309_ (.A0(_00954_),
    .A1(_00956_),
    .S(_03128_),
    .X(_01090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20310_ (.A0(_00950_),
    .A1(_00953_),
    .S(_03128_),
    .X(_01088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20311_ (.A0(_01082_),
    .A1(_00941_),
    .S(_03128_),
    .X(_01083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20312_ (.A0(_03114_),
    .A1(_03122_),
    .S(_03135_),
    .X(_01082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20313_ (.A0(_01051_),
    .A1(_03129_),
    .S(_02853_),
    .X(_01052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20314_ (.A0(_01052_),
    .A1(_01010_),
    .S(_03159_),
    .X(_01053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20315_ (.A0(_01056_),
    .A1(_01068_),
    .S(_00754_),
    .X(_01069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20316_ (.A0(_01069_),
    .A1(_01059_),
    .S(_03273_),
    .X(_01070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20317_ (.A0(_01070_),
    .A1(_01065_),
    .S(_02866_),
    .X(_01071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20318_ (.A0(_01059_),
    .A1(_01056_),
    .S(_02850_),
    .X(_01060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20319_ (.A0(_01060_),
    .A1(_01056_),
    .S(_02849_),
    .X(_01061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20320_ (.A0(_01072_),
    .A1(_02642_),
    .S(_00854_),
    .X(_01073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20321_ (.A0(_01073_),
    .A1(_01009_),
    .S(_02870_),
    .X(_01074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20322_ (.A0(_01074_),
    .A1(_01075_),
    .S(_00857_),
    .X(_01076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20323_ (.A0(_01066_),
    .A1(_01067_),
    .S(\design_top.XADDR[31] ),
    .X(_01068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20324_ (.A0(_00994_),
    .A1(_01063_),
    .S(\design_top.XADDR[3] ),
    .X(_01064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20325_ (.A0(_01062_),
    .A1(_01064_),
    .S(\design_top.XADDR[31] ),
    .X(_01065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20326_ (.A0(_01057_),
    .A1(_01058_),
    .S(\design_top.XADDR[31] ),
    .X(_01059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20327_ (.A0(_01054_),
    .A1(_01055_),
    .S(\design_top.XADDR[31] ),
    .X(_01056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20328_ (.A0(_01038_),
    .A1(_01047_),
    .S(_03111_),
    .X(_01048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20329_ (.A0(_01041_),
    .A1(_01046_),
    .S(_03120_),
    .X(_01047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20330_ (.A0(_01042_),
    .A1(_02684_),
    .S(_03128_),
    .X(_01046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20331_ (.A0(_01038_),
    .A1(_01044_),
    .S(_03111_),
    .X(_01045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20332_ (.A0(_01041_),
    .A1(_01043_),
    .S(_03120_),
    .X(_01044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20333_ (.A0(_01042_),
    .A1(_00820_),
    .S(_03128_),
    .X(_01043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20334_ (.A0(_02888_),
    .A1(_02879_),
    .S(_03135_),
    .X(_01042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20335_ (.A0(_01039_),
    .A1(_01040_),
    .S(_03128_),
    .X(_01041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20336_ (.A0(_02905_),
    .A1(_02897_),
    .S(_03135_),
    .X(_01040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20337_ (.A0(_02922_),
    .A1(_02914_),
    .S(_03135_),
    .X(_01039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20338_ (.A0(_01034_),
    .A1(_01037_),
    .S(_03120_),
    .X(_01038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20339_ (.A0(_01035_),
    .A1(_01036_),
    .S(_03128_),
    .X(_01037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20340_ (.A0(_02939_),
    .A1(_02931_),
    .S(_03135_),
    .X(_01036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20341_ (.A0(_02956_),
    .A1(_02948_),
    .S(_03135_),
    .X(_01035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20342_ (.A0(_01032_),
    .A1(_01033_),
    .S(_03128_),
    .X(_01034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20343_ (.A0(_02973_),
    .A1(_02965_),
    .S(_03135_),
    .X(_01033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20344_ (.A0(_02990_),
    .A1(_02982_),
    .S(_03135_),
    .X(_01032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20345_ (.A0(_03122_),
    .A1(_03114_),
    .S(_03135_),
    .X(_01017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20346_ (.A0(_01017_),
    .A1(_01018_),
    .S(_03128_),
    .X(_01019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20347_ (.A0(_01019_),
    .A1(_01022_),
    .S(_03120_),
    .X(_01023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20348_ (.A0(_01023_),
    .A1(_01030_),
    .S(_03111_),
    .X(_01031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20349_ (.A0(_01026_),
    .A1(_01029_),
    .S(_03120_),
    .X(_01030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20350_ (.A0(_01027_),
    .A1(_01028_),
    .S(_03128_),
    .X(_01029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20351_ (.A0(_03007_),
    .A1(_02999_),
    .S(_03135_),
    .X(_01028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20352_ (.A0(_03024_),
    .A1(_03016_),
    .S(_03135_),
    .X(_01027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20353_ (.A0(_01024_),
    .A1(_01025_),
    .S(_03128_),
    .X(_01026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20354_ (.A0(_00803_),
    .A1(_03033_),
    .S(_03135_),
    .X(_01025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20355_ (.A0(_00805_),
    .A1(_03049_),
    .S(_03135_),
    .X(_01024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20356_ (.A0(_01020_),
    .A1(_01021_),
    .S(_03128_),
    .X(_01022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20357_ (.A0(_00809_),
    .A1(_03065_),
    .S(_03135_),
    .X(_01021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20358_ (.A0(_00811_),
    .A1(_03081_),
    .S(_03135_),
    .X(_01020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20359_ (.A0(_03105_),
    .A1(_03097_),
    .S(_03135_),
    .X(_01018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20360_ (.A0(_00977_),
    .A1(_00945_),
    .S(_02847_),
    .X(_00978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20361_ (.A0(_00978_),
    .A1(_00940_),
    .S(_02852_),
    .X(_00979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20362_ (.A0(_00979_),
    .A1(_03136_),
    .S(_00827_),
    .X(_00980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20363_ (.A0(_00980_),
    .A1(_03158_),
    .S(_00828_),
    .X(_00981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20364_ (.A0(_00981_),
    .A1(_00940_),
    .S(_02853_),
    .X(_00982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20365_ (.A0(_00982_),
    .A1(_00939_),
    .S(_03159_),
    .X(_00983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20366_ (.A0(_00987_),
    .A1(_01000_),
    .S(_00754_),
    .X(_01001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20367_ (.A0(_01001_),
    .A1(_00990_),
    .S(_03273_),
    .X(_01002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20368_ (.A0(_01002_),
    .A1(_00997_),
    .S(_02866_),
    .X(_01003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20369_ (.A0(_00990_),
    .A1(_00987_),
    .S(_02850_),
    .X(_00991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20370_ (.A0(_00991_),
    .A1(_00987_),
    .S(_02849_),
    .X(_00992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20371_ (.A0(_01004_),
    .A1(_02643_),
    .S(_00854_),
    .X(_01005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20372_ (.A0(_01005_),
    .A1(_00937_),
    .S(_02870_),
    .X(_01006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20373_ (.A0(_01006_),
    .A1(_01007_),
    .S(_00857_),
    .X(_01008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20374_ (.A0(_00998_),
    .A1(_00999_),
    .S(\design_top.XADDR[31] ),
    .X(_01000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20375_ (.A0(_00994_),
    .A1(_00995_),
    .S(\design_top.XADDR[3] ),
    .X(_00996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20376_ (.A0(_00993_),
    .A1(_00996_),
    .S(\design_top.XADDR[31] ),
    .X(_00997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20377_ (.A0(_00988_),
    .A1(_00989_),
    .S(\design_top.XADDR[31] ),
    .X(_00990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20378_ (.A0(_00984_),
    .A1(_00986_),
    .S(\design_top.XADDR[31] ),
    .X(_00987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20379_ (.A0(_03162_),
    .A1(_03122_),
    .S(_03135_),
    .X(_00946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20380_ (.A0(_00946_),
    .A1(_00947_),
    .S(_03128_),
    .X(_00948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20381_ (.A0(_00948_),
    .A1(_00951_),
    .S(_03120_),
    .X(_00952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20382_ (.A0(_00952_),
    .A1(_00959_),
    .S(_03111_),
    .X(_00960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20383_ (.A0(_00960_),
    .A1(_00975_),
    .S(_03103_),
    .X(_00976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20384_ (.A0(_00967_),
    .A1(_00974_),
    .S(_03111_),
    .X(_00975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20385_ (.A0(_00970_),
    .A1(_00973_),
    .S(_03120_),
    .X(_00974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20386_ (.A0(_00971_),
    .A1(_00972_),
    .S(_03128_),
    .X(_00973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20387_ (.A0(_02879_),
    .A1(_02684_),
    .S(_03135_),
    .X(_00972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20388_ (.A0(_02897_),
    .A1(_02888_),
    .S(_03135_),
    .X(_00971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20389_ (.A0(_00968_),
    .A1(_00969_),
    .S(_03128_),
    .X(_00970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20390_ (.A0(_02914_),
    .A1(_02905_),
    .S(_03135_),
    .X(_00969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20391_ (.A0(_02931_),
    .A1(_02922_),
    .S(_03135_),
    .X(_00968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20392_ (.A0(_00963_),
    .A1(_00966_),
    .S(_03120_),
    .X(_00967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20393_ (.A0(_00964_),
    .A1(_00965_),
    .S(_03128_),
    .X(_00966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20394_ (.A0(_02948_),
    .A1(_02939_),
    .S(_03135_),
    .X(_00965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20395_ (.A0(_02965_),
    .A1(_02956_),
    .S(_03135_),
    .X(_00964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20396_ (.A0(_00961_),
    .A1(_00962_),
    .S(_03128_),
    .X(_00963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20397_ (.A0(_02982_),
    .A1(_02973_),
    .S(_03135_),
    .X(_00962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20398_ (.A0(_02999_),
    .A1(_02990_),
    .S(_03135_),
    .X(_00961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20399_ (.A0(_00955_),
    .A1(_00958_),
    .S(_03120_),
    .X(_00959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20400_ (.A0(_00956_),
    .A1(_00957_),
    .S(_03128_),
    .X(_00958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20401_ (.A0(_03016_),
    .A1(_03007_),
    .S(_03135_),
    .X(_00957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20402_ (.A0(_03033_),
    .A1(_03024_),
    .S(_03135_),
    .X(_00956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20403_ (.A0(_00953_),
    .A1(_00954_),
    .S(_03128_),
    .X(_00955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20404_ (.A0(_03049_),
    .A1(_00803_),
    .S(_03135_),
    .X(_00954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20405_ (.A0(_03065_),
    .A1(_00805_),
    .S(_03135_),
    .X(_00953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20406_ (.A0(_00949_),
    .A1(_00950_),
    .S(_03128_),
    .X(_00951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20407_ (.A0(_03081_),
    .A1(_00809_),
    .S(_03135_),
    .X(_00950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20408_ (.A0(_03097_),
    .A1(_00811_),
    .S(_03135_),
    .X(_00949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20409_ (.A0(_03114_),
    .A1(_03105_),
    .S(_03135_),
    .X(_00947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20410_ (.A0(\design_top.core0.XIDATA[10] ),
    .A1(\design_top.core0.RESMODE[3] ),
    .S(\design_top.core0.XRES ),
    .X(_00863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20411_ (.A0(\design_top.core0.XIDATA[9] ),
    .A1(\design_top.core0.RESMODE[2] ),
    .S(\design_top.core0.XRES ),
    .X(_00862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20412_ (.A0(\design_top.core0.XIDATA[8] ),
    .A1(\design_top.core0.RESMODE[1] ),
    .S(\design_top.core0.XRES ),
    .X(_00861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20413_ (.A0(\design_top.core0.XIDATA[7] ),
    .A1(\design_top.core0.RESMODE[0] ),
    .S(\design_top.core0.XRES ),
    .X(_00860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20414_ (.A0(_00829_),
    .A1(_03188_),
    .S(_02853_),
    .X(_00830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20415_ (.A0(_00830_),
    .A1(_02877_),
    .S(_03159_),
    .X(_00831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20416_ (.A0(_00841_),
    .A1(_00836_),
    .S(_02849_),
    .X(_00842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20417_ (.A0(_00853_),
    .A1(_00780_),
    .S(_00854_),
    .X(_00855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20418_ (.A0(_00855_),
    .A1(_00779_),
    .S(_02870_),
    .X(_00856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20419_ (.A0(_00856_),
    .A1(_00858_),
    .S(_00857_),
    .X(_00859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20420_ (.A0(_00848_),
    .A1(_00839_),
    .S(_00754_),
    .X(_00849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20421_ (.A0(_00849_),
    .A1(_00845_),
    .S(_03273_),
    .X(_00850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20422_ (.A0(_00850_),
    .A1(_00836_),
    .S(_02866_),
    .X(_00851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20423_ (.A0(_00846_),
    .A1(_00847_),
    .S(\design_top.XADDR[31] ),
    .X(_00848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20424_ (.A0(_00843_),
    .A1(_00844_),
    .S(\design_top.XADDR[31] ),
    .X(_00845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20425_ (.A0(_00836_),
    .A1(_00839_),
    .S(_02850_),
    .X(_00840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20426_ (.A0(_00837_),
    .A1(_00838_),
    .S(\design_top.XADDR[31] ),
    .X(_00839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20427_ (.A0(_00834_),
    .A1(_03198_),
    .S(_00833_),
    .X(_00835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20428_ (.A0(_00832_),
    .A1(_00835_),
    .S(\design_top.XADDR[31] ),
    .X(_00836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20429_ (.A0(_00824_),
    .A1(_02684_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_00825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20430_ (.A0(_02684_),
    .A1(_02879_),
    .S(_03135_),
    .X(_00785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20431_ (.A0(_00785_),
    .A1(_00786_),
    .S(_03128_),
    .X(_00787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20432_ (.A0(_00787_),
    .A1(_00790_),
    .S(_03120_),
    .X(_00791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20433_ (.A0(_00791_),
    .A1(_00798_),
    .S(_03111_),
    .X(_00799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20434_ (.A0(_00799_),
    .A1(_00818_),
    .S(_03103_),
    .X(_00819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20435_ (.A0(_00808_),
    .A1(_00817_),
    .S(_03111_),
    .X(_00818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20436_ (.A0(_00813_),
    .A1(_00816_),
    .S(_03120_),
    .X(_00817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20437_ (.A0(_00814_),
    .A1(_00815_),
    .S(_03128_),
    .X(_00816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20438_ (.A0(_03122_),
    .A1(_03162_),
    .S(_03135_),
    .X(_00815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20439_ (.A0(_03105_),
    .A1(_03114_),
    .S(_03135_),
    .X(_00814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20440_ (.A0(_00810_),
    .A1(_00812_),
    .S(_03128_),
    .X(_00813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20441_ (.A0(_00811_),
    .A1(_03097_),
    .S(_03135_),
    .X(_00812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20442_ (.A0(_00809_),
    .A1(_03081_),
    .S(_03135_),
    .X(_00810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20443_ (.A0(_00802_),
    .A1(_00807_),
    .S(_03120_),
    .X(_00808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20444_ (.A0(_00804_),
    .A1(_00806_),
    .S(_03128_),
    .X(_00807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20445_ (.A0(_00805_),
    .A1(_03065_),
    .S(_03135_),
    .X(_00806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20446_ (.A0(_00803_),
    .A1(_03049_),
    .S(_03135_),
    .X(_00804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20447_ (.A0(_00800_),
    .A1(_00801_),
    .S(_03128_),
    .X(_00802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20448_ (.A0(_03024_),
    .A1(_03033_),
    .S(_03135_),
    .X(_00801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20449_ (.A0(_03007_),
    .A1(_03016_),
    .S(_03135_),
    .X(_00800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20450_ (.A0(_00794_),
    .A1(_00797_),
    .S(_03120_),
    .X(_00798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20451_ (.A0(_00795_),
    .A1(_00796_),
    .S(_03128_),
    .X(_00797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20452_ (.A0(_02990_),
    .A1(_02999_),
    .S(_03135_),
    .X(_00796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20453_ (.A0(_02973_),
    .A1(_02982_),
    .S(_03135_),
    .X(_00795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20454_ (.A0(_00792_),
    .A1(_00793_),
    .S(_03128_),
    .X(_00794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20455_ (.A0(_02956_),
    .A1(_02965_),
    .S(_03135_),
    .X(_00793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20456_ (.A0(_02939_),
    .A1(_02948_),
    .S(_03135_),
    .X(_00792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20457_ (.A0(_00788_),
    .A1(_00789_),
    .S(_03128_),
    .X(_00790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20458_ (.A0(_02922_),
    .A1(_02931_),
    .S(_03135_),
    .X(_00789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20459_ (.A0(_02905_),
    .A1(_02914_),
    .S(_03135_),
    .X(_00788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20460_ (.A0(_02888_),
    .A1(_02897_),
    .S(_03135_),
    .X(_00786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20461_ (.A0(_00752_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_00753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20462_ (.A0(_00750_),
    .A1(_03936_),
    .S(_00008_),
    .X(_00751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20463_ (.A0(_00748_),
    .A1(\design_top.IDATA[18] ),
    .S(_00008_),
    .X(_00749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20464_ (.A0(_00746_),
    .A1(\design_top.IDATA[17] ),
    .S(_00008_),
    .X(_00747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20465_ (.A0(_00744_),
    .A1(\design_top.IDATA[16] ),
    .S(_00008_),
    .X(_00745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20466_ (.A0(_00742_),
    .A1(\design_top.IDATA[15] ),
    .S(_00008_),
    .X(_00743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20467_ (.A0(_00740_),
    .A1(\design_top.IDATA[14] ),
    .S(_00008_),
    .X(_00741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20468_ (.A0(_00738_),
    .A1(\design_top.IDATA[13] ),
    .S(_00008_),
    .X(_00739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20469_ (.A0(_00735_),
    .A1(\design_top.IDATA[12] ),
    .S(_00008_),
    .X(_00736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20470_ (.A0(_00736_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20471_ (.A0(\design_top.ROMFF[11] ),
    .A1(\design_top.ROMFF2[11] ),
    .S(\design_top.HLT2 ),
    .X(_00710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20472_ (.A0(\design_top.ROMFF[29] ),
    .A1(\design_top.ROMFF2[29] ),
    .S(\design_top.HLT2 ),
    .X(_00693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20473_ (.A0(\design_top.ROMFF[28] ),
    .A1(\design_top.ROMFF2[28] ),
    .S(\design_top.HLT2 ),
    .X(_03968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20474_ (.A0(\design_top.ROMFF[27] ),
    .A1(\design_top.ROMFF2[27] ),
    .S(\design_top.HLT2 ),
    .X(_03964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20475_ (.A0(\design_top.ROMFF[26] ),
    .A1(\design_top.ROMFF2[26] ),
    .S(\design_top.HLT2 ),
    .X(_03960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20476_ (.A0(\design_top.ROMFF[25] ),
    .A1(\design_top.ROMFF2[25] ),
    .S(\design_top.HLT2 ),
    .X(_03956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20477_ (.A0(\design_top.ROMFF[24] ),
    .A1(\design_top.ROMFF2[24] ),
    .S(\design_top.HLT2 ),
    .X(_03952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20478_ (.A0(\design_top.ROMFF[19] ),
    .A1(\design_top.ROMFF2[19] ),
    .S(\design_top.HLT2 ),
    .X(_03936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20479_ (.A0(\design_top.ROMFF[6] ),
    .A1(\design_top.ROMFF2[6] ),
    .S(\design_top.HLT2 ),
    .X(_03272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20480_ (.A0(\design_top.ROMFF[5] ),
    .A1(\design_top.ROMFF2[5] ),
    .S(\design_top.HLT2 ),
    .X(_03271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20481_ (.A0(\design_top.ROMFF[4] ),
    .A1(\design_top.ROMFF2[4] ),
    .S(\design_top.HLT2 ),
    .X(_03270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20482_ (.A0(_03200_),
    .A1(_02851_),
    .S(_02854_),
    .X(_03201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20483_ (.A0(_00940_),
    .A1(_03189_),
    .S(_02852_),
    .X(_03190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20484_ (.A0(_03190_),
    .A1(_03160_),
    .S(_03161_),
    .X(_03191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20485_ (.A0(_03191_),
    .A1(_03158_),
    .S(_03159_),
    .X(_03192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20486_ (.A0(_03192_),
    .A1(_03137_),
    .S(_02848_),
    .X(_03193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20487_ (.A0(_03193_),
    .A1(_03136_),
    .S(_02853_),
    .X(_03194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20488_ (.A0(_03038_),
    .A1(\design_top.core0.UIMM[12] ),
    .S(\design_top.core0.XMCC ),
    .X(_03157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20489_ (.A0(_03029_),
    .A1(\design_top.core0.UIMM[13] ),
    .S(\design_top.core0.XMCC ),
    .X(_03156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20490_ (.A0(_03021_),
    .A1(\design_top.core0.UIMM[14] ),
    .S(\design_top.core0.XMCC ),
    .X(_03155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20491_ (.A0(_03012_),
    .A1(\design_top.core0.UIMM[15] ),
    .S(\design_top.core0.XMCC ),
    .X(_03154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20492_ (.A0(_03004_),
    .A1(\design_top.core0.UIMM[16] ),
    .S(\design_top.core0.XMCC ),
    .X(_03153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20493_ (.A0(_02995_),
    .A1(\design_top.core0.UIMM[17] ),
    .S(\design_top.core0.XMCC ),
    .X(_03152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20494_ (.A0(_02987_),
    .A1(\design_top.core0.UIMM[18] ),
    .S(\design_top.core0.XMCC ),
    .X(_03151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20495_ (.A0(_02978_),
    .A1(\design_top.core0.UIMM[19] ),
    .S(\design_top.core0.XMCC ),
    .X(_03150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20496_ (.A0(_02970_),
    .A1(\design_top.core0.UIMM[20] ),
    .S(\design_top.core0.XMCC ),
    .X(_03149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20497_ (.A0(_02961_),
    .A1(\design_top.core0.UIMM[21] ),
    .S(\design_top.core0.XMCC ),
    .X(_03148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20498_ (.A0(_02953_),
    .A1(\design_top.core0.UIMM[22] ),
    .S(\design_top.core0.XMCC ),
    .X(_03147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20499_ (.A0(_02944_),
    .A1(\design_top.core0.UIMM[23] ),
    .S(\design_top.core0.XMCC ),
    .X(_03146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20500_ (.A0(_02936_),
    .A1(\design_top.core0.UIMM[24] ),
    .S(\design_top.core0.XMCC ),
    .X(_03145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20501_ (.A0(_02927_),
    .A1(\design_top.core0.UIMM[25] ),
    .S(\design_top.core0.XMCC ),
    .X(_03144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20502_ (.A0(_02919_),
    .A1(\design_top.core0.UIMM[26] ),
    .S(\design_top.core0.XMCC ),
    .X(_03143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20503_ (.A0(_02910_),
    .A1(\design_top.core0.UIMM[27] ),
    .S(\design_top.core0.XMCC ),
    .X(_03142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20504_ (.A0(_02902_),
    .A1(\design_top.core0.UIMM[28] ),
    .S(\design_top.core0.XMCC ),
    .X(_03141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20505_ (.A0(_02893_),
    .A1(\design_top.core0.UIMM[29] ),
    .S(\design_top.core0.XMCC ),
    .X(_03140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20506_ (.A0(_02884_),
    .A1(\design_top.core0.UIMM[30] ),
    .S(\design_top.core0.XMCC ),
    .X(_03139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20507_ (.A0(_02875_),
    .A1(\design_top.core0.UIMM[31] ),
    .S(\design_top.core0.XMCC ),
    .X(_03138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20508_ (.A0(_03134_),
    .A1(\design_top.core0.SIMM[0] ),
    .S(\design_top.core0.XMCC ),
    .X(_03135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20509_ (.A0(_03127_),
    .A1(\design_top.core0.SIMM[1] ),
    .S(\design_top.core0.XMCC ),
    .X(_03128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20510_ (.A0(_03119_),
    .A1(\design_top.core0.SIMM[2] ),
    .S(\design_top.core0.XMCC ),
    .X(_03120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20511_ (.A0(_03110_),
    .A1(\design_top.core0.SIMM[3] ),
    .S(\design_top.core0.XMCC ),
    .X(_03111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20512_ (.A0(_03102_),
    .A1(\design_top.core0.SIMM[4] ),
    .S(\design_top.core0.XMCC ),
    .X(_03103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20513_ (.A0(_03093_),
    .A1(\design_top.core0.SIMM[5] ),
    .S(\design_top.core0.XMCC ),
    .X(_03094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20514_ (.A0(_03086_),
    .A1(\design_top.core0.SIMM[6] ),
    .S(\design_top.core0.XMCC ),
    .X(_03087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20515_ (.A0(_03077_),
    .A1(\design_top.core0.SIMM[7] ),
    .S(\design_top.core0.XMCC ),
    .X(_03078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20516_ (.A0(_03070_),
    .A1(\design_top.core0.SIMM[8] ),
    .S(\design_top.core0.XMCC ),
    .X(_03071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20517_ (.A0(_03061_),
    .A1(\design_top.core0.SIMM[9] ),
    .S(\design_top.core0.XMCC ),
    .X(_03062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20518_ (.A0(_03054_),
    .A1(\design_top.core0.SIMM[10] ),
    .S(\design_top.core0.XMCC ),
    .X(_03055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20519_ (.A0(_03045_),
    .A1(\design_top.core0.SIMM[11] ),
    .S(\design_top.core0.XMCC ),
    .X(_03046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20520_ (.A0(_03038_),
    .A1(\design_top.core0.SIMM[12] ),
    .S(\design_top.core0.XMCC ),
    .X(_03039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20521_ (.A0(_03029_),
    .A1(\design_top.core0.SIMM[13] ),
    .S(\design_top.core0.XMCC ),
    .X(_03030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20522_ (.A0(_03021_),
    .A1(\design_top.core0.SIMM[14] ),
    .S(\design_top.core0.XMCC ),
    .X(_03022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20523_ (.A0(_03012_),
    .A1(\design_top.core0.SIMM[15] ),
    .S(\design_top.core0.XMCC ),
    .X(_03013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20524_ (.A0(_03004_),
    .A1(\design_top.core0.SIMM[16] ),
    .S(\design_top.core0.XMCC ),
    .X(_03005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20525_ (.A0(_02995_),
    .A1(\design_top.core0.SIMM[17] ),
    .S(\design_top.core0.XMCC ),
    .X(_02996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20526_ (.A0(_02987_),
    .A1(\design_top.core0.SIMM[18] ),
    .S(\design_top.core0.XMCC ),
    .X(_02988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20527_ (.A0(_02978_),
    .A1(\design_top.core0.SIMM[19] ),
    .S(\design_top.core0.XMCC ),
    .X(_02979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20528_ (.A0(_02970_),
    .A1(\design_top.core0.SIMM[20] ),
    .S(\design_top.core0.XMCC ),
    .X(_02971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20529_ (.A0(_02961_),
    .A1(\design_top.core0.SIMM[21] ),
    .S(\design_top.core0.XMCC ),
    .X(_02962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20530_ (.A0(_02953_),
    .A1(\design_top.core0.SIMM[22] ),
    .S(\design_top.core0.XMCC ),
    .X(_02954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20531_ (.A0(_02944_),
    .A1(\design_top.core0.SIMM[23] ),
    .S(\design_top.core0.XMCC ),
    .X(_02945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20532_ (.A0(_02936_),
    .A1(\design_top.core0.SIMM[24] ),
    .S(\design_top.core0.XMCC ),
    .X(_02937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20533_ (.A0(_02927_),
    .A1(\design_top.core0.SIMM[25] ),
    .S(\design_top.core0.XMCC ),
    .X(_02928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20534_ (.A0(_02919_),
    .A1(\design_top.core0.SIMM[26] ),
    .S(\design_top.core0.XMCC ),
    .X(_02920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20535_ (.A0(_02910_),
    .A1(\design_top.core0.SIMM[27] ),
    .S(\design_top.core0.XMCC ),
    .X(_02911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20536_ (.A0(_02902_),
    .A1(\design_top.core0.SIMM[28] ),
    .S(\design_top.core0.XMCC ),
    .X(_02903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20537_ (.A0(_02893_),
    .A1(\design_top.core0.SIMM[29] ),
    .S(\design_top.core0.XMCC ),
    .X(_02894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20538_ (.A0(_02884_),
    .A1(\design_top.core0.SIMM[30] ),
    .S(\design_top.core0.XMCC ),
    .X(_02885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20539_ (.A0(_02875_),
    .A1(\design_top.core0.SIMM[31] ),
    .S(\design_top.core0.XMCC ),
    .X(_02876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20540_ (.A0(_02867_),
    .A1(_02863_),
    .S(_02854_),
    .X(_02868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20541_ (.A0(_02864_),
    .A1(_02863_),
    .S(_02854_),
    .X(_02865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20542_ (.A0(_02856_),
    .A1(_02851_),
    .S(_02854_),
    .X(_02857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20543_ (.A0(_02655_),
    .A1(_02658_),
    .S(_00688_),
    .X(_02659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20544_ (.A0(_02656_),
    .A1(_02657_),
    .S(_00687_),
    .X(_02658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20545_ (.A0(_02653_),
    .A1(_02654_),
    .S(_00687_),
    .X(_02655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20546_ (.A0(_02646_),
    .A1(_02649_),
    .S(_00688_),
    .X(_02650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20547_ (.A0(_02647_),
    .A1(_02648_),
    .S(_00687_),
    .X(_02649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20548_ (.A0(_02644_),
    .A1(_02645_),
    .S(_00687_),
    .X(_02646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20549_ (.A0(_02637_),
    .A1(_02640_),
    .S(_00688_),
    .X(_02641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20550_ (.A0(_02638_),
    .A1(_02639_),
    .S(_00687_),
    .X(_02640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20551_ (.A0(_02635_),
    .A1(_02636_),
    .S(_00687_),
    .X(_02637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20552_ (.A0(_02630_),
    .A1(_02633_),
    .S(_00688_),
    .X(_02634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20553_ (.A0(_02631_),
    .A1(_02632_),
    .S(_00687_),
    .X(_02633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20554_ (.A0(_02628_),
    .A1(_02629_),
    .S(_00687_),
    .X(_02630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20555_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_03260_),
    .X(_00180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20556_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_03260_),
    .X(_00179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20557_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_03260_),
    .X(_00178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20558_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_03260_),
    .X(_00177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20559_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_03260_),
    .X(_00176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20560_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_03260_),
    .X(_00175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20561_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_03260_),
    .X(_00174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20562_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_03260_),
    .X(_00173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20563_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_03243_),
    .X(_00284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20564_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_03243_),
    .X(_00283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20565_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_03243_),
    .X(_00282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20566_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_03243_),
    .X(_00281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20567_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_03243_),
    .X(_00280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20568_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_03243_),
    .X(_00279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20569_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_03243_),
    .X(_00278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20570_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_03243_),
    .X(_00277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20571_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_03241_),
    .X(_00292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20572_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_03241_),
    .X(_00291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20573_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_03241_),
    .X(_00290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20574_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_03241_),
    .X(_00289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20575_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_03241_),
    .X(_00288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20576_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_03241_),
    .X(_00287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20577_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_03241_),
    .X(_00286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20578_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_03241_),
    .X(_00285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20579_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_03222_),
    .X(_00300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20580_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_03222_),
    .X(_00299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20581_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_03222_),
    .X(_00298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20582_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_03222_),
    .X(_00297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20583_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_03222_),
    .X(_00296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20584_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_03222_),
    .X(_00295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20585_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_03222_),
    .X(_00294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20586_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_03222_),
    .X(_00293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20587_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_03220_),
    .X(_00308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20588_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_03220_),
    .X(_00307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20589_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_03220_),
    .X(_00306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20590_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_03220_),
    .X(_00305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20591_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_03220_),
    .X(_00304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20592_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_03220_),
    .X(_00303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20593_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_03220_),
    .X(_00302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20594_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_03220_),
    .X(_00301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20595_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_03218_),
    .X(_00316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20596_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_03218_),
    .X(_00315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20597_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_03218_),
    .X(_00314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20598_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_03218_),
    .X(_00313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20599_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_03218_),
    .X(_00312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20600_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_03218_),
    .X(_00311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20601_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_03218_),
    .X(_00310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20602_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_03218_),
    .X(_00309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20603_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_03217_),
    .X(_00324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20604_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_03217_),
    .X(_00323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20605_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_03217_),
    .X(_00322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20606_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_03217_),
    .X(_00321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20607_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_03217_),
    .X(_00320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20608_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_03217_),
    .X(_00319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20609_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_03217_),
    .X(_00318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20610_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_03217_),
    .X(_00317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20611_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_03266_),
    .X(_00332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20612_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_03266_),
    .X(_00331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20613_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_03266_),
    .X(_00330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20614_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_03266_),
    .X(_00329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20615_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_03266_),
    .X(_00328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20616_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_03266_),
    .X(_00327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20617_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_03266_),
    .X(_00326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20618_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_03266_),
    .X(_00325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20619_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_03263_),
    .X(_00356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20620_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_03263_),
    .X(_00355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20621_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_03263_),
    .X(_00354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20622_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_03263_),
    .X(_00353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20623_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_03263_),
    .X(_00352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20624_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_03263_),
    .X(_00351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20625_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_03263_),
    .X(_00350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20626_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_03263_),
    .X(_00349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20627_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_03233_),
    .X(_00444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20628_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_03233_),
    .X(_00443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20629_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_03233_),
    .X(_00442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20630_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_03233_),
    .X(_00441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20631_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_03233_),
    .X(_00440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20632_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_03233_),
    .X(_00439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20633_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_03233_),
    .X(_00438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20634_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_03233_),
    .X(_00437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20635_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_03227_),
    .X(_00532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20636_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_03227_),
    .X(_00531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20637_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_03227_),
    .X(_00530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20638_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_03227_),
    .X(_00529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20639_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_03227_),
    .X(_00528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20640_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_03227_),
    .X(_00527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20641_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_03227_),
    .X(_00526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20642_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_03227_),
    .X(_00525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20643_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_03207_),
    .X(_00620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20644_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_03207_),
    .X(_00619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20645_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_03207_),
    .X(_00618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20646_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_03207_),
    .X(_00617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20647_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_03207_),
    .X(_00616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20648_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_03207_),
    .X(_00615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20649_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_03207_),
    .X(_00614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20650_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_03207_),
    .X(_00613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20651_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_03212_),
    .X(_00660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20652_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_03212_),
    .X(_00659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20653_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_03212_),
    .X(_00658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20654_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_03212_),
    .X(_00657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20655_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_03212_),
    .X(_00656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20656_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_03212_),
    .X(_00655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20657_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_03212_),
    .X(_00654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20658_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_03212_),
    .X(_00653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20659_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_03213_),
    .X(_00668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20660_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_03213_),
    .X(_00667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20661_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_03213_),
    .X(_00666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20662_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_03213_),
    .X(_00665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20663_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_03213_),
    .X(_00664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20664_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_03213_),
    .X(_00663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20665_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_03213_),
    .X(_00662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20666_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_03213_),
    .X(_00661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20667_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_03214_),
    .X(_00676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20668_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_03214_),
    .X(_00675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20669_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_03214_),
    .X(_00674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20670_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_03214_),
    .X(_00673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20671_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_03214_),
    .X(_00672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20672_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_03214_),
    .X(_00671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20673_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_03214_),
    .X(_00670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20674_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_03214_),
    .X(_00669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20675_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_03265_),
    .X(_00340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20676_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_03265_),
    .X(_00339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20677_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_03265_),
    .X(_00338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20678_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_03265_),
    .X(_00337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20679_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_03265_),
    .X(_00336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20680_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_03265_),
    .X(_00335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20681_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_03265_),
    .X(_00334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20682_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_03265_),
    .X(_00333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20683_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_03264_),
    .X(_00348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20684_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_03264_),
    .X(_00347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20685_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_03264_),
    .X(_00346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20686_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_03264_),
    .X(_00345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20687_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_03264_),
    .X(_00344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20688_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_03264_),
    .X(_00343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20689_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_03264_),
    .X(_00342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20690_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_03264_),
    .X(_00341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20691_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_03215_),
    .X(_00684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20692_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_03215_),
    .X(_00683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20693_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_03215_),
    .X(_00682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20694_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_03215_),
    .X(_00681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20695_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_03215_),
    .X(_00680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20696_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_03215_),
    .X(_00679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20697_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_03215_),
    .X(_00678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20698_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_03215_),
    .X(_00677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20699_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_03259_),
    .X(_00188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20700_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_03259_),
    .X(_00187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20701_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_03259_),
    .X(_00186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20702_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_03259_),
    .X(_00185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20703_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_03259_),
    .X(_00184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20704_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_03259_),
    .X(_00183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20705_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_03259_),
    .X(_00182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20706_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_03259_),
    .X(_00181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20707_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_03262_),
    .X(_00364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20708_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_03262_),
    .X(_00363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20709_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_03262_),
    .X(_00362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20710_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_03262_),
    .X(_00361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20711_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_03262_),
    .X(_00360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20712_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_03262_),
    .X(_00359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20713_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_03262_),
    .X(_00358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20714_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_03262_),
    .X(_00357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20715_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_03226_),
    .X(_00476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20716_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_03226_),
    .X(_00475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20717_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_03226_),
    .X(_00474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20718_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_03226_),
    .X(_00473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20719_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_03226_),
    .X(_00472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20720_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_03226_),
    .X(_00471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20721_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_03226_),
    .X(_00470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20722_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_03226_),
    .X(_00469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20723_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_03257_),
    .X(_00204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20724_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_03257_),
    .X(_00203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20725_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_03257_),
    .X(_00202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20726_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_03257_),
    .X(_00201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20727_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_03257_),
    .X(_00200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20728_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_03257_),
    .X(_00199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20729_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_03257_),
    .X(_00198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20730_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_03257_),
    .X(_00197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20731_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_03256_),
    .X(_00212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20732_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_03256_),
    .X(_00211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20733_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_03256_),
    .X(_00210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20734_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_03256_),
    .X(_00209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20735_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_03256_),
    .X(_00208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20736_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_03256_),
    .X(_00207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20737_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_03256_),
    .X(_00206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20738_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_03256_),
    .X(_00205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20739_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_03261_),
    .X(_00372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20740_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_03261_),
    .X(_00371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20741_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_03261_),
    .X(_00370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20742_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_03261_),
    .X(_00369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20743_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_03261_),
    .X(_00368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20744_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_03261_),
    .X(_00367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20745_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_03261_),
    .X(_00366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20746_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_03261_),
    .X(_00365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20747_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_03255_),
    .X(_00220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20748_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_03255_),
    .X(_00219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20749_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_03255_),
    .X(_00218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20750_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_03255_),
    .X(_00217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20751_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_03255_),
    .X(_00216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20752_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_03255_),
    .X(_00215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20753_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_03255_),
    .X(_00214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20754_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_03255_),
    .X(_00213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20755_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_03254_),
    .X(_00228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20756_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_03254_),
    .X(_00227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20757_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_03254_),
    .X(_00226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20758_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_03254_),
    .X(_00225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20759_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_03254_),
    .X(_00224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20760_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_03254_),
    .X(_00223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20761_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_03254_),
    .X(_00222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20762_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_03254_),
    .X(_00221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20763_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_03225_),
    .X(_00540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20764_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_03225_),
    .X(_00539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20765_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_03225_),
    .X(_00538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20766_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_03225_),
    .X(_00537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20767_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_03225_),
    .X(_00536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20768_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_03225_),
    .X(_00535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20769_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_03225_),
    .X(_00534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20770_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_03225_),
    .X(_00533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20771_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_03258_),
    .X(_00196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20772_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_03258_),
    .X(_00195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20773_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_03258_),
    .X(_00194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20774_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_03258_),
    .X(_00193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20775_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_03258_),
    .X(_00192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20776_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_03258_),
    .X(_00191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20777_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_03258_),
    .X(_00190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20778_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_03258_),
    .X(_00189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20779_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_03239_),
    .X(_00548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20780_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_03239_),
    .X(_00547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20781_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_03239_),
    .X(_00546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20782_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_03239_),
    .X(_00545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20783_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_03239_),
    .X(_00544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20784_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_03239_),
    .X(_00543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20785_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_03239_),
    .X(_00542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20786_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_03239_),
    .X(_00541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20787_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_03238_),
    .X(_00572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20788_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_03238_),
    .X(_00571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20789_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_03238_),
    .X(_00570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20790_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_03238_),
    .X(_00569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20791_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_03238_),
    .X(_00568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20792_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_03238_),
    .X(_00567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20793_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_03238_),
    .X(_00566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20794_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_03238_),
    .X(_00565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20795_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_03237_),
    .X(_00556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20796_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_03237_),
    .X(_00555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20797_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_03237_),
    .X(_00554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20798_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_03237_),
    .X(_00553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20799_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_03237_),
    .X(_00552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20800_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_03237_),
    .X(_00551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20801_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_03237_),
    .X(_00550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20802_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_03237_),
    .X(_00549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20803_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_03202_),
    .X(_00580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20804_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_03202_),
    .X(_00579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20805_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_03202_),
    .X(_00578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20806_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_03202_),
    .X(_00577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20807_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_03202_),
    .X(_00576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20808_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_03202_),
    .X(_00575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20809_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_03202_),
    .X(_00574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20810_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_03202_),
    .X(_00573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20811_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_03240_),
    .X(_00564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20812_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_03240_),
    .X(_00563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20813_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_03240_),
    .X(_00562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20814_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_03240_),
    .X(_00561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20815_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_03240_),
    .X(_00560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20816_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_03240_),
    .X(_00559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20817_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_03240_),
    .X(_00558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20818_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_03240_),
    .X(_00557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20819_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_03224_),
    .X(_00484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20820_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_03224_),
    .X(_00483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20821_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_03224_),
    .X(_00482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20822_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_03224_),
    .X(_00481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20823_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_03224_),
    .X(_00480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20824_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_03224_),
    .X(_00479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20825_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_03224_),
    .X(_00478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20826_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_03224_),
    .X(_00477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20827_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_03246_),
    .X(_00404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20828_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_03246_),
    .X(_00403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20829_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_03246_),
    .X(_00402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20830_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_03246_),
    .X(_00401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20831_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_03246_),
    .X(_00400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20832_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_03246_),
    .X(_00399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20833_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_03246_),
    .X(_00398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20834_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_03246_),
    .X(_00397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20835_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_03242_),
    .X(_00412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20836_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_03242_),
    .X(_00411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20837_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_03242_),
    .X(_00410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20838_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_03242_),
    .X(_00409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20839_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_03242_),
    .X(_00408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20840_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_03242_),
    .X(_00407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20841_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_03242_),
    .X(_00406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20842_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_03242_),
    .X(_00405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20843_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_03223_),
    .X(_00492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20844_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_03223_),
    .X(_00491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20845_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_03223_),
    .X(_00490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20846_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_03223_),
    .X(_00489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20847_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_03223_),
    .X(_00488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20848_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_03223_),
    .X(_00487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20849_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_03223_),
    .X(_00486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20850_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_03223_),
    .X(_00485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20851_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_03221_),
    .X(_00420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20852_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_03221_),
    .X(_00419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20853_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_03221_),
    .X(_00418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20854_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_03221_),
    .X(_00417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20855_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_03221_),
    .X(_00416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20856_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_03221_),
    .X(_00415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20857_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_03221_),
    .X(_00414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20858_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_03221_),
    .X(_00413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20859_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_03235_),
    .X(_00500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20860_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_03235_),
    .X(_00499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20861_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_03235_),
    .X(_00498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20862_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_03235_),
    .X(_00497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20863_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_03235_),
    .X(_00496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20864_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_03235_),
    .X(_00495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20865_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_03235_),
    .X(_00494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20866_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_03235_),
    .X(_00493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20867_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_03219_),
    .X(_00428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20868_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_03219_),
    .X(_00427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20869_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_03219_),
    .X(_00426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20870_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_03219_),
    .X(_00425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20871_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_03219_),
    .X(_00424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20872_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_03219_),
    .X(_00423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20873_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_03219_),
    .X(_00422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20874_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_03219_),
    .X(_00421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20875_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_03234_),
    .X(_00508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20876_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_03234_),
    .X(_00507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20877_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_03234_),
    .X(_00506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20878_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_03234_),
    .X(_00505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20879_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_03234_),
    .X(_00504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20880_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_03234_),
    .X(_00503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20881_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_03234_),
    .X(_00502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20882_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_03234_),
    .X(_00501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20883_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_03236_),
    .X(_00436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20884_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_03236_),
    .X(_00435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20885_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_03236_),
    .X(_00434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20886_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_03236_),
    .X(_00433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20887_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_03236_),
    .X(_00432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20888_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_03236_),
    .X(_00431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20889_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_03236_),
    .X(_00430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20890_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_03236_),
    .X(_00429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20891_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_03231_),
    .X(_00516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20892_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_03231_),
    .X(_00515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20893_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_03231_),
    .X(_00514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20894_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_03231_),
    .X(_00513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20895_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_03231_),
    .X(_00512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20896_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_03231_),
    .X(_00511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20897_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_03231_),
    .X(_00510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20898_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_03231_),
    .X(_00509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20899_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_03232_),
    .X(_00452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20900_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_03232_),
    .X(_00451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20901_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_03232_),
    .X(_00450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20902_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_03232_),
    .X(_00449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20903_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_03232_),
    .X(_00448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20904_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_03232_),
    .X(_00447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20905_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_03232_),
    .X(_00446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20906_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_03232_),
    .X(_00445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20907_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_03229_),
    .X(_00524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20908_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_03229_),
    .X(_00523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20909_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_03229_),
    .X(_00522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20910_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_03229_),
    .X(_00521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20911_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_03229_),
    .X(_00520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20912_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_03229_),
    .X(_00519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20913_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_03229_),
    .X(_00518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20914_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_03229_),
    .X(_00517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20915_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_03230_),
    .X(_00460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20916_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_03230_),
    .X(_00459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20917_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_03230_),
    .X(_00458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20918_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_03230_),
    .X(_00457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20919_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_03230_),
    .X(_00456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20920_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_03230_),
    .X(_00455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20921_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_03230_),
    .X(_00454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20922_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_03230_),
    .X(_00453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20923_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_03228_),
    .X(_00468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20924_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_03228_),
    .X(_00467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20925_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_03228_),
    .X(_00466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20926_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_03228_),
    .X(_00465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20927_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_03228_),
    .X(_00464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20928_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_03228_),
    .X(_00463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20929_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_03228_),
    .X(_00462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20930_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_03228_),
    .X(_00461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20931_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_03252_),
    .X(_00380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20932_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_03252_),
    .X(_00379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20933_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_03252_),
    .X(_00378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20934_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_03252_),
    .X(_00377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20935_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_03252_),
    .X(_00376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20936_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_03252_),
    .X(_00375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20937_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_03252_),
    .X(_00374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20938_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_03252_),
    .X(_00373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20939_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_03253_),
    .X(_00236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20940_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_03253_),
    .X(_00235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20941_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_03253_),
    .X(_00234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20942_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_03253_),
    .X(_00233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20943_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_03253_),
    .X(_00232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20944_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_03253_),
    .X(_00231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20945_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_03253_),
    .X(_00230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20946_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_03253_),
    .X(_00229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20947_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_03251_),
    .X(_00388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20948_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_03251_),
    .X(_00387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20949_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_03251_),
    .X(_00386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20950_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_03251_),
    .X(_00385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20951_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_03251_),
    .X(_00384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20952_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_03251_),
    .X(_00383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20953_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_03251_),
    .X(_00382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20954_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_03251_),
    .X(_00381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20955_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_03250_),
    .X(_00244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20956_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_03250_),
    .X(_00243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20957_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_03250_),
    .X(_00242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20958_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_03250_),
    .X(_00241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20959_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_03250_),
    .X(_00240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20960_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_03250_),
    .X(_00239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20961_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_03250_),
    .X(_00238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20962_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_03250_),
    .X(_00237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20963_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_03249_),
    .X(_00252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20964_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_03249_),
    .X(_00251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20965_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_03249_),
    .X(_00250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20966_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_03249_),
    .X(_00249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20967_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_03249_),
    .X(_00248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20968_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_03249_),
    .X(_00247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20969_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_03249_),
    .X(_00246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20970_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_03249_),
    .X(_00245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20971_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_03247_),
    .X(_00396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20972_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_03247_),
    .X(_00395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20973_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_03247_),
    .X(_00394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20974_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_03247_),
    .X(_00393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20975_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_03247_),
    .X(_00392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20976_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_03247_),
    .X(_00391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20977_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_03247_),
    .X(_00390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20978_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_03247_),
    .X(_00389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20979_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_03248_),
    .X(_00260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20980_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_03248_),
    .X(_00259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20981_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_03248_),
    .X(_00258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20982_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_03248_),
    .X(_00257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20983_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_03248_),
    .X(_00256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20984_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_03248_),
    .X(_00255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20985_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_03248_),
    .X(_00254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20986_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_03248_),
    .X(_00253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20987_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_03244_),
    .X(_00276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20988_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_03244_),
    .X(_00275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20989_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_03244_),
    .X(_00274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20990_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_03244_),
    .X(_00273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20991_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_03244_),
    .X(_00272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20992_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_03244_),
    .X(_00271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20993_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_03244_),
    .X(_00270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20994_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_03244_),
    .X(_00269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20995_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_03211_),
    .X(_00652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20996_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_03211_),
    .X(_00651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20997_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_03211_),
    .X(_00650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20998_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_03211_),
    .X(_00649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _20999_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_03211_),
    .X(_00648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21000_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_03211_),
    .X(_00647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21001_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_03211_),
    .X(_00646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21002_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_03211_),
    .X(_00645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21003_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_03210_),
    .X(_00644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21004_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_03210_),
    .X(_00643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21005_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_03210_),
    .X(_00642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21006_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_03210_),
    .X(_00641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21007_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_03210_),
    .X(_00640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21008_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_03210_),
    .X(_00639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21009_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_03210_),
    .X(_00638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21010_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_03210_),
    .X(_00637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21011_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_03209_),
    .X(_00636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21012_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_03209_),
    .X(_00635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21013_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_03209_),
    .X(_00634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21014_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_03209_),
    .X(_00633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21015_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_03209_),
    .X(_00632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21016_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_03209_),
    .X(_00631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21017_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_03209_),
    .X(_00630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21018_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_03209_),
    .X(_00629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21019_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_03208_),
    .X(_00628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21020_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_03208_),
    .X(_00627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21021_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_03208_),
    .X(_00626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21022_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_03208_),
    .X(_00625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21023_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_03208_),
    .X(_00624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21024_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_03208_),
    .X(_00623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21025_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_03208_),
    .X(_00622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21026_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_03208_),
    .X(_00621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21027_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_03206_),
    .X(_00612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21028_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_03206_),
    .X(_00611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21029_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_03206_),
    .X(_00610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21030_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_03206_),
    .X(_00609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21031_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_03206_),
    .X(_00608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21032_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_03206_),
    .X(_00607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21033_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_03206_),
    .X(_00606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21034_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_03206_),
    .X(_00605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21035_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_03205_),
    .X(_00604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21036_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_03205_),
    .X(_00603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21037_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_03205_),
    .X(_00602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21038_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_03205_),
    .X(_00601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21039_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_03205_),
    .X(_00600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21040_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_03205_),
    .X(_00599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21041_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_03205_),
    .X(_00598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21042_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_03205_),
    .X(_00597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21043_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_03204_),
    .X(_00596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21044_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_03204_),
    .X(_00595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21045_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_03204_),
    .X(_00594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21046_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_03204_),
    .X(_00593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21047_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_03204_),
    .X(_00592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21048_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_03204_),
    .X(_00591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21049_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_03204_),
    .X(_00590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21050_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_03204_),
    .X(_00589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21051_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_03203_),
    .X(_00588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21052_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_03203_),
    .X(_00587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21053_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_03203_),
    .X(_00586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21054_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_03203_),
    .X(_00585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21055_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_03203_),
    .X(_00584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21056_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_03203_),
    .X(_00583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21057_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_03203_),
    .X(_00582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21058_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_03203_),
    .X(_00581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21059_ (.A0(_01982_),
    .A1(io_out[12]),
    .S(_02858_),
    .X(_00012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21060_ (.A0(\design_top.IDATA[18] ),
    .A1(\design_top.core0.S1PTR[3] ),
    .S(\design_top.HLT ),
    .X(_00003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21061_ (.A0(\design_top.IDATA[21] ),
    .A1(\design_top.core0.S2PTR[1] ),
    .S(\design_top.HLT ),
    .X(_00005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21062_ (.A0(_01981_),
    .A1(\design_top.IOMUX[3][31] ),
    .S(_03197_),
    .X(_00037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21063_ (.A0(_01980_),
    .A1(\design_top.IOMUX[3][30] ),
    .S(_03197_),
    .X(_00036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21064_ (.A0(_01979_),
    .A1(\design_top.IOMUX[3][29] ),
    .S(_03197_),
    .X(_00034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21065_ (.A0(_01978_),
    .A1(\design_top.IOMUX[3][28] ),
    .S(_03197_),
    .X(_00033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21066_ (.A0(_01977_),
    .A1(\design_top.IOMUX[3][27] ),
    .S(_03197_),
    .X(_00032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21067_ (.A0(_01976_),
    .A1(\design_top.IOMUX[3][26] ),
    .S(_03197_),
    .X(_00031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21068_ (.A0(_01975_),
    .A1(\design_top.IOMUX[3][25] ),
    .S(_03197_),
    .X(_00030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21069_ (.A0(_01974_),
    .A1(\design_top.IOMUX[3][24] ),
    .S(_03197_),
    .X(_00029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21070_ (.A0(_01973_),
    .A1(\design_top.IOMUX[3][23] ),
    .S(_03197_),
    .X(_00028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21071_ (.A0(_01972_),
    .A1(\design_top.IOMUX[3][22] ),
    .S(_03197_),
    .X(_00027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21072_ (.A0(_01971_),
    .A1(\design_top.IOMUX[3][21] ),
    .S(_03197_),
    .X(_00026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21073_ (.A0(_01970_),
    .A1(\design_top.IOMUX[3][20] ),
    .S(_03197_),
    .X(_00025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21074_ (.A0(_01969_),
    .A1(\design_top.IOMUX[3][19] ),
    .S(_03197_),
    .X(_00023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21075_ (.A0(_01968_),
    .A1(\design_top.IOMUX[3][18] ),
    .S(_03197_),
    .X(_00022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21076_ (.A0(_01967_),
    .A1(\design_top.IOMUX[3][17] ),
    .S(_03197_),
    .X(_00021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21077_ (.A0(_01966_),
    .A1(\design_top.IOMUX[3][16] ),
    .S(_03197_),
    .X(_00020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21078_ (.A0(_01965_),
    .A1(\design_top.IOMUX[3][15] ),
    .S(_03197_),
    .X(_00019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21079_ (.A0(_01964_),
    .A1(\design_top.IOMUX[3][14] ),
    .S(_03197_),
    .X(_00018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21080_ (.A0(_01963_),
    .A1(\design_top.IOMUX[3][13] ),
    .S(_03197_),
    .X(_00017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21081_ (.A0(_01962_),
    .A1(\design_top.IOMUX[3][12] ),
    .S(_03197_),
    .X(_00016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21082_ (.A0(_01961_),
    .A1(\design_top.IOMUX[3][11] ),
    .S(_03197_),
    .X(_00015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21083_ (.A0(_01960_),
    .A1(\design_top.IOMUX[3][10] ),
    .S(_03197_),
    .X(_00014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21084_ (.A0(_01959_),
    .A1(\design_top.IOMUX[3][9] ),
    .S(_03197_),
    .X(_00044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21085_ (.A0(_01958_),
    .A1(\design_top.IOMUX[3][8] ),
    .S(_03197_),
    .X(_00043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21086_ (.A0(_01957_),
    .A1(\design_top.IOMUX[3][7] ),
    .S(_03197_),
    .X(_00042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21087_ (.A0(_01956_),
    .A1(\design_top.IOMUX[3][6] ),
    .S(_03197_),
    .X(_00041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21088_ (.A0(_01955_),
    .A1(\design_top.IOMUX[3][5] ),
    .S(_03197_),
    .X(_00040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21089_ (.A0(_01954_),
    .A1(\design_top.IOMUX[3][4] ),
    .S(_03197_),
    .X(_00039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21090_ (.A0(_01953_),
    .A1(\design_top.IOMUX[3][3] ),
    .S(_03197_),
    .X(_00038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21091_ (.A0(_01952_),
    .A1(\design_top.IOMUX[3][2] ),
    .S(_03197_),
    .X(_00035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21092_ (.A0(_01951_),
    .A1(\design_top.IOMUX[3][1] ),
    .S(_03197_),
    .X(_00024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21093_ (.A0(_01950_),
    .A1(\design_top.IOMUX[3][0] ),
    .S(_03197_),
    .X(_00013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21094_ (.A0(\design_top.IDATA[17] ),
    .A1(\design_top.core0.S1PTR[2] ),
    .S(\design_top.HLT ),
    .X(_00002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21095_ (.A0(\design_top.IDATA[20] ),
    .A1(\design_top.core0.S2PTR[0] ),
    .S(\design_top.HLT ),
    .X(_00004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21096_ (.A0(_01943_),
    .A1(\design_top.DADDR[31] ),
    .S(_02869_),
    .X(_01944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21097_ (.A0(_01944_),
    .A1(_01942_),
    .S(_03195_),
    .X(_00101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21098_ (.A0(_01939_),
    .A1(_01940_),
    .S(_02869_),
    .X(_01941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21099_ (.A0(_01941_),
    .A1(_01938_),
    .S(_03195_),
    .X(_00100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21100_ (.A0(_01935_),
    .A1(_01936_),
    .S(_02869_),
    .X(_01937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21101_ (.A0(_01937_),
    .A1(_01934_),
    .S(_03195_),
    .X(_00098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21102_ (.A0(_01931_),
    .A1(_01932_),
    .S(_02869_),
    .X(_01933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21103_ (.A0(_01933_),
    .A1(_01930_),
    .S(_03195_),
    .X(_00097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21104_ (.A0(_01927_),
    .A1(_01928_),
    .S(_02869_),
    .X(_01929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21105_ (.A0(_01929_),
    .A1(_01926_),
    .S(_03195_),
    .X(_00096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21106_ (.A0(_01923_),
    .A1(_01924_),
    .S(_02869_),
    .X(_01925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21107_ (.A0(_01925_),
    .A1(_01922_),
    .S(_03195_),
    .X(_00095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21108_ (.A0(_01919_),
    .A1(_01920_),
    .S(_02869_),
    .X(_01921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21109_ (.A0(_01921_),
    .A1(_01918_),
    .S(_03195_),
    .X(_00094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21110_ (.A0(_01915_),
    .A1(_01916_),
    .S(_02869_),
    .X(_01917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21111_ (.A0(_01917_),
    .A1(_01914_),
    .S(_03195_),
    .X(_00093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21112_ (.A0(_01911_),
    .A1(_01912_),
    .S(_02869_),
    .X(_01913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21113_ (.A0(_01913_),
    .A1(_01910_),
    .S(_03195_),
    .X(_00092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21114_ (.A0(_01907_),
    .A1(_01908_),
    .S(_02869_),
    .X(_01909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21115_ (.A0(_01909_),
    .A1(_01906_),
    .S(_03195_),
    .X(_00091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21116_ (.A0(_01903_),
    .A1(_01904_),
    .S(_02869_),
    .X(_01905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21117_ (.A0(_01905_),
    .A1(_01902_),
    .S(_03195_),
    .X(_00090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21118_ (.A0(_01899_),
    .A1(_01900_),
    .S(_02869_),
    .X(_01901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21119_ (.A0(_01901_),
    .A1(_01898_),
    .S(_03195_),
    .X(_00089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21120_ (.A0(_01895_),
    .A1(_01896_),
    .S(_02869_),
    .X(_01897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21121_ (.A0(_01897_),
    .A1(_01894_),
    .S(_03195_),
    .X(_00088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21122_ (.A0(_01891_),
    .A1(_01892_),
    .S(_02869_),
    .X(_01893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21123_ (.A0(_01893_),
    .A1(_01890_),
    .S(_03195_),
    .X(_00087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21124_ (.A0(_01887_),
    .A1(_01888_),
    .S(_02869_),
    .X(_01889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21125_ (.A0(_01889_),
    .A1(_01886_),
    .S(_03195_),
    .X(_00086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21126_ (.A0(_01883_),
    .A1(_01884_),
    .S(_02869_),
    .X(_01885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21127_ (.A0(_01885_),
    .A1(_01882_),
    .S(_03195_),
    .X(_00085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21128_ (.A0(_01879_),
    .A1(_01880_),
    .S(_02869_),
    .X(_01881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21129_ (.A0(_01881_),
    .A1(_01878_),
    .S(_03195_),
    .X(_00084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21130_ (.A0(_01875_),
    .A1(_01876_),
    .S(_02869_),
    .X(_01877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21131_ (.A0(_01877_),
    .A1(_01874_),
    .S(_03195_),
    .X(_00083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21132_ (.A0(_01871_),
    .A1(_01872_),
    .S(_02869_),
    .X(_01873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21133_ (.A0(_01873_),
    .A1(_01870_),
    .S(_03195_),
    .X(_00082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21134_ (.A0(_01867_),
    .A1(_01868_),
    .S(_02869_),
    .X(_01869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21135_ (.A0(_01869_),
    .A1(_01866_),
    .S(_03195_),
    .X(_00081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21136_ (.A0(_01863_),
    .A1(_01864_),
    .S(_02869_),
    .X(_01865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21137_ (.A0(_01865_),
    .A1(_01862_),
    .S(_03195_),
    .X(_00080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21138_ (.A0(_01859_),
    .A1(_01860_),
    .S(_02869_),
    .X(_01861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21139_ (.A0(_01861_),
    .A1(_01858_),
    .S(_03195_),
    .X(_00079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21140_ (.A0(_01855_),
    .A1(_01856_),
    .S(_02869_),
    .X(_01857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21141_ (.A0(_01857_),
    .A1(_01854_),
    .S(_03195_),
    .X(_00108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21142_ (.A0(_01851_),
    .A1(_01852_),
    .S(_02869_),
    .X(_01853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21143_ (.A0(_01853_),
    .A1(_01850_),
    .S(_03195_),
    .X(_00107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21144_ (.A0(_01848_),
    .A1(_01847_),
    .S(_02869_),
    .X(_01849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21145_ (.A0(_01849_),
    .A1(_01846_),
    .S(_03195_),
    .X(_00106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21146_ (.A0(_01844_),
    .A1(_03216_),
    .S(_02869_),
    .X(_01845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21147_ (.A0(_01845_),
    .A1(_01843_),
    .S(_03195_),
    .X(_00105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21148_ (.A0(_01841_),
    .A1(_03199_),
    .S(_02869_),
    .X(_01842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21149_ (.A0(_01842_),
    .A1(_01840_),
    .S(_03195_),
    .X(_00104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21150_ (.A0(_01838_),
    .A1(_01837_),
    .S(_02869_),
    .X(_01839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21151_ (.A0(_01839_),
    .A1(_01836_),
    .S(_03195_),
    .X(_00103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21152_ (.A0(_01834_),
    .A1(\design_top.DADDR[3] ),
    .S(_02869_),
    .X(_01835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21153_ (.A0(_01835_),
    .A1(_01833_),
    .S(_03195_),
    .X(_00102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21154_ (.A0(_01831_),
    .A1(\design_top.DADDR[2] ),
    .S(_02869_),
    .X(_01832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21155_ (.A0(_01832_),
    .A1(_01830_),
    .S(_03195_),
    .X(_00099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21156_ (.A0(_01473_),
    .A1(_01474_),
    .S(\design_top.core0.XRES ),
    .X(_00045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21157_ (.A0(_00936_),
    .A1(_00935_),
    .S(_02661_),
    .X(_00011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21158_ (.A0(_00933_),
    .A1(_03196_),
    .S(_00934_),
    .X(_00078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21159_ (.A0(\design_top.IDATA[15] ),
    .A1(\design_top.core0.S1PTR[0] ),
    .S(\design_top.HLT ),
    .X(_00000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21160_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_03245_),
    .X(_00268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21161_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_03245_),
    .X(_00267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21162_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_03245_),
    .X(_00266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21163_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_03245_),
    .X(_00265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21164_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_03245_),
    .X(_00264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21165_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_03245_),
    .X(_00263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21166_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_03245_),
    .X(_00262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21167_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_03245_),
    .X(_00261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21168_ (.A0(_00732_),
    .A1(\design_top.IDATA[20] ),
    .S(_00008_),
    .X(_00733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21169_ (.A0(_00733_),
    .A1(\design_top.IDATA[7] ),
    .S(_00009_),
    .X(_00734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21170_ (.A0(_00734_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21171_ (.A0(_00729_),
    .A1(\design_top.IDATA[30] ),
    .S(_00008_),
    .X(_00730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21172_ (.A0(_00730_),
    .A1(\design_top.IDATA[30] ),
    .S(_00009_),
    .X(_00731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21173_ (.A0(_00731_),
    .A1(\design_top.IDATA[30] ),
    .S(_00010_),
    .X(_00048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21174_ (.A0(_00726_),
    .A1(_00693_),
    .S(_00008_),
    .X(_00727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21175_ (.A0(_00727_),
    .A1(_00693_),
    .S(_00009_),
    .X(_00728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21176_ (.A0(_00728_),
    .A1(_00693_),
    .S(_00010_),
    .X(_00077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21177_ (.A0(_00723_),
    .A1(_03968_),
    .S(_00008_),
    .X(_00724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21178_ (.A0(_00724_),
    .A1(_03968_),
    .S(_00009_),
    .X(_00725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21179_ (.A0(_00725_),
    .A1(_03968_),
    .S(_00010_),
    .X(_00076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21180_ (.A0(_00720_),
    .A1(_03964_),
    .S(_00008_),
    .X(_00721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21181_ (.A0(_00721_),
    .A1(_03964_),
    .S(_00009_),
    .X(_00722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21182_ (.A0(_00722_),
    .A1(_03964_),
    .S(_00010_),
    .X(_00075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21183_ (.A0(_00717_),
    .A1(_03960_),
    .S(_00008_),
    .X(_00718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21184_ (.A0(_00718_),
    .A1(_03960_),
    .S(_00009_),
    .X(_00719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21185_ (.A0(_00719_),
    .A1(_03960_),
    .S(_00010_),
    .X(_00074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21186_ (.A0(_00714_),
    .A1(_03956_),
    .S(_00008_),
    .X(_00715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21187_ (.A0(_00715_),
    .A1(_03956_),
    .S(_00009_),
    .X(_00716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21188_ (.A0(_00716_),
    .A1(_03956_),
    .S(_00010_),
    .X(_00073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21189_ (.A0(_00711_),
    .A1(_03952_),
    .S(_00008_),
    .X(_00712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21190_ (.A0(_00712_),
    .A1(_00710_),
    .S(_00009_),
    .X(_00713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21191_ (.A0(_00713_),
    .A1(_00710_),
    .S(_00010_),
    .X(_00072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21192_ (.A0(_00707_),
    .A1(\design_top.IDATA[23] ),
    .S(_00008_),
    .X(_00708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21193_ (.A0(_00708_),
    .A1(\design_top.IDATA[10] ),
    .S(_00009_),
    .X(_00709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21194_ (.A0(_00709_),
    .A1(\design_top.IDATA[10] ),
    .S(_00010_),
    .X(_00071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21195_ (.A0(_00704_),
    .A1(\design_top.IDATA[22] ),
    .S(_00008_),
    .X(_00705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21196_ (.A0(_00705_),
    .A1(\design_top.IDATA[9] ),
    .S(_00009_),
    .X(_00706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21197_ (.A0(_00706_),
    .A1(\design_top.IDATA[9] ),
    .S(_00010_),
    .X(_00069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21198_ (.A0(_00701_),
    .A1(\design_top.IDATA[21] ),
    .S(_00008_),
    .X(_00702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21199_ (.A0(_00702_),
    .A1(\design_top.IDATA[8] ),
    .S(_00009_),
    .X(_00703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21200_ (.A0(_00703_),
    .A1(\design_top.IDATA[8] ),
    .S(_00010_),
    .X(_00058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21201_ (.A0(_00700_),
    .A1(\design_top.IDATA[7] ),
    .S(_00010_),
    .X(_00047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21202_ (.A0(\design_top.IDATA[16] ),
    .A1(\design_top.core0.S1PTR[1] ),
    .S(\design_top.HLT ),
    .X(_00001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21203_ (.A0(\design_top.IDATA[30] ),
    .A1(\design_top.IDATA[31] ),
    .S(_03914_),
    .X(_00697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21204_ (.A0(_00697_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_00698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21205_ (.A0(_00698_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21206_ (.A0(_00699_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21207_ (.A0(_00693_),
    .A1(\design_top.IDATA[31] ),
    .S(_03914_),
    .X(_00694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21208_ (.A0(_00694_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_00695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21209_ (.A0(_00695_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21210_ (.A0(_00696_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21211_ (.A0(_03968_),
    .A1(\design_top.IDATA[31] ),
    .S(_03914_),
    .X(_03969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21212_ (.A0(_03969_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_03970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21213_ (.A0(_03970_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_03971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21214_ (.A0(_03971_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21215_ (.A0(_03964_),
    .A1(\design_top.IDATA[31] ),
    .S(_03914_),
    .X(_03965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21216_ (.A0(_03965_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_03966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21217_ (.A0(_03966_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_03967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21218_ (.A0(_03967_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21219_ (.A0(_03960_),
    .A1(\design_top.IDATA[31] ),
    .S(_03914_),
    .X(_03961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21220_ (.A0(_03961_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_03962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21221_ (.A0(_03962_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_03963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21222_ (.A0(_03963_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21223_ (.A0(_03956_),
    .A1(\design_top.IDATA[31] ),
    .S(_03914_),
    .X(_03957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21224_ (.A0(_03957_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_03958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21225_ (.A0(_03958_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_03959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21226_ (.A0(_03959_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21227_ (.A0(_03952_),
    .A1(\design_top.IDATA[31] ),
    .S(_03914_),
    .X(_03953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21228_ (.A0(_03953_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_03954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21229_ (.A0(_03954_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_03955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21230_ (.A0(_03955_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21231_ (.A0(\design_top.IDATA[23] ),
    .A1(\design_top.IDATA[31] ),
    .S(_03914_),
    .X(_03949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21232_ (.A0(_03949_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_03950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21233_ (.A0(_03950_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_03951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21234_ (.A0(_03951_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21235_ (.A0(\design_top.IDATA[22] ),
    .A1(\design_top.IDATA[31] ),
    .S(_03914_),
    .X(_03946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21236_ (.A0(_03946_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_03947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21237_ (.A0(_03947_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_03948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21238_ (.A0(_03948_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21239_ (.A0(\design_top.IDATA[21] ),
    .A1(\design_top.IDATA[31] ),
    .S(_03914_),
    .X(_03943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21240_ (.A0(_03943_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_03944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21241_ (.A0(_03944_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_03945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21242_ (.A0(_03945_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21243_ (.A0(\design_top.IDATA[20] ),
    .A1(\design_top.IDATA[31] ),
    .S(_03914_),
    .X(_03940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21244_ (.A0(_03940_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_03941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21245_ (.A0(_03941_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_03942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21246_ (.A0(_03942_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21247_ (.A0(_03936_),
    .A1(\design_top.IDATA[31] ),
    .S(_03914_),
    .X(_03937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21248_ (.A0(_03937_),
    .A1(_03936_),
    .S(_00008_),
    .X(_03938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21249_ (.A0(_03938_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_03939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21250_ (.A0(_03939_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21251_ (.A0(\design_top.IDATA[18] ),
    .A1(\design_top.IDATA[31] ),
    .S(_03914_),
    .X(_03933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21252_ (.A0(_03933_),
    .A1(\design_top.IDATA[18] ),
    .S(_00008_),
    .X(_03934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21253_ (.A0(_03934_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_03935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21254_ (.A0(_03935_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21255_ (.A0(\design_top.IDATA[17] ),
    .A1(\design_top.IDATA[31] ),
    .S(_03914_),
    .X(_03930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21256_ (.A0(_03930_),
    .A1(\design_top.IDATA[17] ),
    .S(_00008_),
    .X(_03931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21257_ (.A0(_03931_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_03932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21258_ (.A0(_03932_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21259_ (.A0(\design_top.IDATA[16] ),
    .A1(\design_top.IDATA[31] ),
    .S(_03914_),
    .X(_03927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21260_ (.A0(_03927_),
    .A1(\design_top.IDATA[16] ),
    .S(_00008_),
    .X(_03928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21261_ (.A0(_03928_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_03929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21262_ (.A0(_03929_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21263_ (.A0(\design_top.IDATA[15] ),
    .A1(\design_top.IDATA[31] ),
    .S(_03914_),
    .X(_03924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21264_ (.A0(_03924_),
    .A1(\design_top.IDATA[15] ),
    .S(_00008_),
    .X(_03925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21265_ (.A0(_03925_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_03926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21266_ (.A0(_03926_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21267_ (.A0(\design_top.IDATA[14] ),
    .A1(\design_top.IDATA[31] ),
    .S(_03914_),
    .X(_03921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21268_ (.A0(_03921_),
    .A1(\design_top.IDATA[14] ),
    .S(_00008_),
    .X(_03922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21269_ (.A0(_03922_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_03923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21270_ (.A0(_03923_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21271_ (.A0(\design_top.IDATA[13] ),
    .A1(\design_top.IDATA[31] ),
    .S(_03914_),
    .X(_03918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21272_ (.A0(_03918_),
    .A1(\design_top.IDATA[13] ),
    .S(_00008_),
    .X(_03919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21273_ (.A0(_03919_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_03920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21274_ (.A0(_03920_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21275_ (.A0(\design_top.IDATA[12] ),
    .A1(\design_top.IDATA[31] ),
    .S(_03914_),
    .X(_03915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21276_ (.A0(_03915_),
    .A1(\design_top.IDATA[12] ),
    .S(_00008_),
    .X(_03916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21277_ (.A0(_03916_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_03917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21278_ (.A0(_03917_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21279_ (.A0(\design_top.IDATA[22] ),
    .A1(\design_top.core0.S2PTR[2] ),
    .S(\design_top.HLT ),
    .X(_00006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _21280_ (.A0(\design_top.IDATA[23] ),
    .A1(\design_top.core0.S2PTR[3] ),
    .S(\design_top.HLT ),
    .X(_00007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21281_ (.A0(\design_top.uart0.UART_XFIFO[0] ),
    .A1(\design_top.uart0.UART_XFIFO[1] ),
    .A2(\design_top.uart0.UART_XFIFO[2] ),
    .A3(\design_top.uart0.UART_XFIFO[3] ),
    .S0(\design_top.uart0.UART_XSTATE[0] ),
    .S1(\design_top.uart0.UART_XSTATE[1] ),
    .X(_01946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21282_ (.A0(\design_top.uart0.UART_XFIFO[4] ),
    .A1(\design_top.uart0.UART_XFIFO[5] ),
    .A2(\design_top.uart0.UART_XFIFO[6] ),
    .A3(\design_top.uart0.UART_XFIFO[7] ),
    .S0(\design_top.uart0.UART_XSTATE[0] ),
    .S1(\design_top.uart0.UART_XSTATE[1] ),
    .X(_01947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21283_ (.A0(_01821_),
    .A1(_02887_),
    .A2(_00852_),
    .A3(_01822_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21284_ (.A0(_01817_),
    .A1(_01814_),
    .A2(_01808_),
    .A3(_01809_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21285_ (.A0(_01800_),
    .A1(_02896_),
    .A2(_00852_),
    .A3(_01801_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21286_ (.A0(_01796_),
    .A1(_01793_),
    .A2(_01788_),
    .A3(_01789_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21287_ (.A0(_01780_),
    .A1(_01766_),
    .A2(_00852_),
    .A3(_01781_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21288_ (.A0(_01776_),
    .A1(_01773_),
    .A2(_01767_),
    .A3(_01768_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21289_ (.A0(_01758_),
    .A1(_02913_),
    .A2(_00852_),
    .A3(_01759_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21290_ (.A0(_01754_),
    .A1(_01751_),
    .A2(_01747_),
    .A3(_01748_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21291_ (.A0(_01739_),
    .A1(_01725_),
    .A2(_00852_),
    .A3(_01740_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21292_ (.A0(_01735_),
    .A1(_01732_),
    .A2(_01726_),
    .A3(_01727_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21293_ (.A0(_01717_),
    .A1(_02930_),
    .A2(_00852_),
    .A3(_01718_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21294_ (.A0(_01713_),
    .A1(_01710_),
    .A2(_01705_),
    .A3(_01706_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21295_ (.A0(_01697_),
    .A1(_01683_),
    .A2(_00852_),
    .A3(_01698_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21296_ (.A0(_01693_),
    .A1(_01690_),
    .A2(_01684_),
    .A3(_01685_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21297_ (.A0(_01675_),
    .A1(_02947_),
    .A2(_00852_),
    .A3(_01676_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21298_ (.A0(_01671_),
    .A1(_01668_),
    .A2(_01665_),
    .A3(_01666_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21299_ (.A0(_01657_),
    .A1(_01643_),
    .A2(_00852_),
    .A3(_01658_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21300_ (.A0(_01653_),
    .A1(_01650_),
    .A2(_01644_),
    .A3(_01645_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21301_ (.A0(_01635_),
    .A1(_02964_),
    .A2(_00852_),
    .A3(_01636_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21302_ (.A0(_01631_),
    .A1(_01628_),
    .A2(_01623_),
    .A3(_01624_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21303_ (.A0(_01615_),
    .A1(_01601_),
    .A2(_00852_),
    .A3(_01616_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21304_ (.A0(_01611_),
    .A1(_01608_),
    .A2(_01602_),
    .A3(_01603_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21305_ (.A0(_01593_),
    .A1(_02981_),
    .A2(_00852_),
    .A3(_01594_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21306_ (.A0(_01589_),
    .A1(_01586_),
    .A2(_01582_),
    .A3(_01583_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21307_ (.A0(_01574_),
    .A1(_01559_),
    .A2(_00852_),
    .A3(_01575_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21308_ (.A0(_01570_),
    .A1(_01567_),
    .A2(_01561_),
    .A3(_01562_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21309_ (.A0(_01551_),
    .A1(_02998_),
    .A2(_00852_),
    .A3(_01552_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21310_ (.A0(_01547_),
    .A1(_01544_),
    .A2(_01539_),
    .A3(_01540_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21311_ (.A0(_01531_),
    .A1(_01517_),
    .A2(_00852_),
    .A3(_01532_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21312_ (.A0(_01527_),
    .A1(_01524_),
    .A2(_01518_),
    .A3(_01519_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21313_ (.A0(_01509_),
    .A1(_03015_),
    .A2(_00852_),
    .A3(_01510_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21314_ (.A0(_01504_),
    .A1(_00823_),
    .A2(_01504_),
    .A3(_02684_),
    .S0(_03103_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21315_ (.A0(_01505_),
    .A1(_01503_),
    .A2(_01501_),
    .A3(_01502_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21316_ (.A0(_01492_),
    .A1(_01476_),
    .A2(_00852_),
    .A3(_01494_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21317_ (.A0(_01485_),
    .A1(_01486_),
    .A2(_01485_),
    .A3(_01487_),
    .S0(_03103_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21318_ (.A0(_01488_),
    .A1(_01484_),
    .A2(_01478_),
    .A3(_01479_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21319_ (.A0(_01465_),
    .A1(_03032_),
    .A2(_00852_),
    .A3(_01467_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21320_ (.A0(_01458_),
    .A1(_01459_),
    .A2(_01458_),
    .A3(_01460_),
    .S0(_03103_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21321_ (.A0(_01461_),
    .A1(_01457_),
    .A2(_01452_),
    .A3(_01453_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21322_ (.A0(_01443_),
    .A1(_01428_),
    .A2(_00852_),
    .A3(_01445_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21323_ (.A0(_01436_),
    .A1(_01437_),
    .A2(_01436_),
    .A3(_01438_),
    .S0(_03103_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21324_ (.A0(_01439_),
    .A1(_01435_),
    .A2(_01429_),
    .A3(_01430_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21325_ (.A0(_01419_),
    .A1(_03048_),
    .A2(_00852_),
    .A3(_01421_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21326_ (.A0(_01412_),
    .A1(_01413_),
    .A2(_01412_),
    .A3(_01414_),
    .S0(_03103_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21327_ (.A0(_01415_),
    .A1(_01411_),
    .A2(_01407_),
    .A3(_01408_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21328_ (.A0(_01398_),
    .A1(_01383_),
    .A2(_00852_),
    .A3(_01400_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21329_ (.A0(_01391_),
    .A1(_01392_),
    .A2(_01391_),
    .A3(_01393_),
    .S0(_03103_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21330_ (.A0(_01394_),
    .A1(_01390_),
    .A2(_01384_),
    .A3(_01385_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21331_ (.A0(_01374_),
    .A1(_03064_),
    .A2(_00852_),
    .A3(_01376_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21332_ (.A0(_01367_),
    .A1(_01368_),
    .A2(_01367_),
    .A3(_01369_),
    .S0(_03103_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21333_ (.A0(_01370_),
    .A1(_01366_),
    .A2(_01361_),
    .A3(_01362_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21334_ (.A0(_01352_),
    .A1(_01337_),
    .A2(_00852_),
    .A3(_01354_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21335_ (.A0(_01345_),
    .A1(_01346_),
    .A2(_01345_),
    .A3(_01347_),
    .S0(_03103_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21336_ (.A0(_01348_),
    .A1(_01344_),
    .A2(_01338_),
    .A3(_01339_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21337_ (.A0(_01328_),
    .A1(_03080_),
    .A2(_00851_),
    .A3(_01330_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21338_ (.A0(_01320_),
    .A1(_01322_),
    .A2(_01320_),
    .A3(_01323_),
    .S0(_03103_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21339_ (.A0(_01324_),
    .A1(_01317_),
    .A2(_01314_),
    .A3(_01315_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21340_ (.A0(_01289_),
    .A1(_01268_),
    .A2(_01307_),
    .A3(_01298_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21341_ (.A0(_01279_),
    .A1(_01282_),
    .A2(_01279_),
    .A3(_01284_),
    .S0(_03103_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21342_ (.A0(_01285_),
    .A1(_01276_),
    .A2(_01270_),
    .A3(_01271_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21343_ (.A0(_01243_),
    .A1(_03096_),
    .A2(_01261_),
    .A3(_01252_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21344_ (.A0(_01233_),
    .A1(_01236_),
    .A2(_01233_),
    .A3(_01238_),
    .S0(_03103_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21345_ (.A0(_01239_),
    .A1(_01230_),
    .A2(_01225_),
    .A3(_01226_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21346_ (.A0(_01201_),
    .A1(_01181_),
    .A2(_01218_),
    .A3(_01209_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21347_ (.A0(_01191_),
    .A1(_01194_),
    .A2(_01191_),
    .A3(_01196_),
    .S0(_03103_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21348_ (.A0(_01197_),
    .A1(_01188_),
    .A2(_01182_),
    .A3(_01183_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21349_ (.A0(_01157_),
    .A1(_03113_),
    .A2(_01174_),
    .A3(_01165_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21350_ (.A0(_01144_),
    .A1(_01150_),
    .A2(_01144_),
    .A3(_01152_),
    .S0(_03103_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21351_ (.A0(_01153_),
    .A1(_01137_),
    .A2(_01133_),
    .A3(_01134_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21352_ (.A0(_01108_),
    .A1(_01078_),
    .A2(_01126_),
    .A3(_01117_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21353_ (.A0(_01093_),
    .A1(_01100_),
    .A2(_01093_),
    .A3(_01103_),
    .S0(_03103_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21354_ (.A0(_01104_),
    .A1(_01086_),
    .A2(_01080_),
    .A3(_01081_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21355_ (.A0(_01053_),
    .A1(_00781_),
    .A2(_01071_),
    .A3(_01061_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21356_ (.A0(_01031_),
    .A1(_01045_),
    .A2(_01031_),
    .A3(_01048_),
    .S0(_03103_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21357_ (.A0(_01049_),
    .A1(_01016_),
    .A2(_01011_),
    .A3(_01012_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_01050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21358_ (.A0(_00983_),
    .A1(_00938_),
    .A2(_01003_),
    .A3(_00992_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_01004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21359_ (.A0(_00831_),
    .A1(_02878_),
    .A2(_00852_),
    .A3(_00842_),
    .S0(_11368_),
    .S1(io_out[12]),
    .X(_00853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21360_ (.A0(_00825_),
    .A1(_00819_),
    .A2(_00782_),
    .A3(_00784_),
    .S0(_11369_),
    .S1(_02852_),
    .X(_00826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21361_ (.A0(\design_top.core0.REG2[0][0] ),
    .A1(\design_top.core0.REG2[1][0] ),
    .A2(\design_top.core0.REG2[2][0] ),
    .A3(\design_top.core0.REG2[3][0] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21362_ (.A0(\design_top.core0.REG2[4][0] ),
    .A1(\design_top.core0.REG2[5][0] ),
    .A2(\design_top.core0.REG2[6][0] ),
    .A3(\design_top.core0.REG2[7][0] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21363_ (.A0(\design_top.core0.REG2[8][0] ),
    .A1(\design_top.core0.REG2[9][0] ),
    .A2(\design_top.core0.REG2[10][0] ),
    .A3(\design_top.core0.REG2[11][0] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21364_ (.A0(\design_top.core0.REG2[12][0] ),
    .A1(\design_top.core0.REG2[13][0] ),
    .A2(\design_top.core0.REG2[14][0] ),
    .A3(\design_top.core0.REG2[15][0] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21365_ (.A0(_03130_),
    .A1(_03131_),
    .A2(_03132_),
    .A3(_03133_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_03134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21366_ (.A0(\design_top.core0.REG2[0][1] ),
    .A1(\design_top.core0.REG2[1][1] ),
    .A2(\design_top.core0.REG2[2][1] ),
    .A3(\design_top.core0.REG2[3][1] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21367_ (.A0(\design_top.core0.REG2[4][1] ),
    .A1(\design_top.core0.REG2[5][1] ),
    .A2(\design_top.core0.REG2[6][1] ),
    .A3(\design_top.core0.REG2[7][1] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21368_ (.A0(\design_top.core0.REG2[8][1] ),
    .A1(\design_top.core0.REG2[9][1] ),
    .A2(\design_top.core0.REG2[10][1] ),
    .A3(\design_top.core0.REG2[11][1] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21369_ (.A0(\design_top.core0.REG2[12][1] ),
    .A1(\design_top.core0.REG2[13][1] ),
    .A2(\design_top.core0.REG2[14][1] ),
    .A3(\design_top.core0.REG2[15][1] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21370_ (.A0(_03123_),
    .A1(_03124_),
    .A2(_03125_),
    .A3(_03126_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_03127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21371_ (.A0(\design_top.core0.REG2[0][2] ),
    .A1(\design_top.core0.REG2[1][2] ),
    .A2(\design_top.core0.REG2[2][2] ),
    .A3(\design_top.core0.REG2[3][2] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21372_ (.A0(\design_top.core0.REG2[4][2] ),
    .A1(\design_top.core0.REG2[5][2] ),
    .A2(\design_top.core0.REG2[6][2] ),
    .A3(\design_top.core0.REG2[7][2] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21373_ (.A0(\design_top.core0.REG2[8][2] ),
    .A1(\design_top.core0.REG2[9][2] ),
    .A2(\design_top.core0.REG2[10][2] ),
    .A3(\design_top.core0.REG2[11][2] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21374_ (.A0(\design_top.core0.REG2[12][2] ),
    .A1(\design_top.core0.REG2[13][2] ),
    .A2(\design_top.core0.REG2[14][2] ),
    .A3(\design_top.core0.REG2[15][2] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21375_ (.A0(_03115_),
    .A1(_03116_),
    .A2(_03117_),
    .A3(_03118_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_03119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21376_ (.A0(\design_top.core0.REG2[0][3] ),
    .A1(\design_top.core0.REG2[1][3] ),
    .A2(\design_top.core0.REG2[2][3] ),
    .A3(\design_top.core0.REG2[3][3] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21377_ (.A0(\design_top.core0.REG2[4][3] ),
    .A1(\design_top.core0.REG2[5][3] ),
    .A2(\design_top.core0.REG2[6][3] ),
    .A3(\design_top.core0.REG2[7][3] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21378_ (.A0(\design_top.core0.REG2[8][3] ),
    .A1(\design_top.core0.REG2[9][3] ),
    .A2(\design_top.core0.REG2[10][3] ),
    .A3(\design_top.core0.REG2[11][3] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21379_ (.A0(\design_top.core0.REG2[12][3] ),
    .A1(\design_top.core0.REG2[13][3] ),
    .A2(\design_top.core0.REG2[14][3] ),
    .A3(\design_top.core0.REG2[15][3] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21380_ (.A0(_03106_),
    .A1(_03107_),
    .A2(_03108_),
    .A3(_03109_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_03110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21381_ (.A0(\design_top.core0.REG2[0][4] ),
    .A1(\design_top.core0.REG2[1][4] ),
    .A2(\design_top.core0.REG2[2][4] ),
    .A3(\design_top.core0.REG2[3][4] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21382_ (.A0(\design_top.core0.REG2[4][4] ),
    .A1(\design_top.core0.REG2[5][4] ),
    .A2(\design_top.core0.REG2[6][4] ),
    .A3(\design_top.core0.REG2[7][4] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21383_ (.A0(\design_top.core0.REG2[8][4] ),
    .A1(\design_top.core0.REG2[9][4] ),
    .A2(\design_top.core0.REG2[10][4] ),
    .A3(\design_top.core0.REG2[11][4] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21384_ (.A0(\design_top.core0.REG2[12][4] ),
    .A1(\design_top.core0.REG2[13][4] ),
    .A2(\design_top.core0.REG2[14][4] ),
    .A3(\design_top.core0.REG2[15][4] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21385_ (.A0(_03098_),
    .A1(_03099_),
    .A2(_03100_),
    .A3(_03101_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_03102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21386_ (.A0(\design_top.core0.REG2[0][5] ),
    .A1(\design_top.core0.REG2[1][5] ),
    .A2(\design_top.core0.REG2[2][5] ),
    .A3(\design_top.core0.REG2[3][5] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21387_ (.A0(\design_top.core0.REG2[4][5] ),
    .A1(\design_top.core0.REG2[5][5] ),
    .A2(\design_top.core0.REG2[6][5] ),
    .A3(\design_top.core0.REG2[7][5] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21388_ (.A0(\design_top.core0.REG2[8][5] ),
    .A1(\design_top.core0.REG2[9][5] ),
    .A2(\design_top.core0.REG2[10][5] ),
    .A3(\design_top.core0.REG2[11][5] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21389_ (.A0(\design_top.core0.REG2[12][5] ),
    .A1(\design_top.core0.REG2[13][5] ),
    .A2(\design_top.core0.REG2[14][5] ),
    .A3(\design_top.core0.REG2[15][5] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21390_ (.A0(_03089_),
    .A1(_03090_),
    .A2(_03091_),
    .A3(_03092_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_03093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21391_ (.A0(\design_top.core0.REG2[0][6] ),
    .A1(\design_top.core0.REG2[1][6] ),
    .A2(\design_top.core0.REG2[2][6] ),
    .A3(\design_top.core0.REG2[3][6] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21392_ (.A0(\design_top.core0.REG2[4][6] ),
    .A1(\design_top.core0.REG2[5][6] ),
    .A2(\design_top.core0.REG2[6][6] ),
    .A3(\design_top.core0.REG2[7][6] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21393_ (.A0(\design_top.core0.REG2[8][6] ),
    .A1(\design_top.core0.REG2[9][6] ),
    .A2(\design_top.core0.REG2[10][6] ),
    .A3(\design_top.core0.REG2[11][6] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21394_ (.A0(\design_top.core0.REG2[12][6] ),
    .A1(\design_top.core0.REG2[13][6] ),
    .A2(\design_top.core0.REG2[14][6] ),
    .A3(\design_top.core0.REG2[15][6] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21395_ (.A0(_03082_),
    .A1(_03083_),
    .A2(_03084_),
    .A3(_03085_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_03086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21396_ (.A0(\design_top.core0.REG2[0][7] ),
    .A1(\design_top.core0.REG2[1][7] ),
    .A2(\design_top.core0.REG2[2][7] ),
    .A3(\design_top.core0.REG2[3][7] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21397_ (.A0(\design_top.core0.REG2[4][7] ),
    .A1(\design_top.core0.REG2[5][7] ),
    .A2(\design_top.core0.REG2[6][7] ),
    .A3(\design_top.core0.REG2[7][7] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21398_ (.A0(\design_top.core0.REG2[8][7] ),
    .A1(\design_top.core0.REG2[9][7] ),
    .A2(\design_top.core0.REG2[10][7] ),
    .A3(\design_top.core0.REG2[11][7] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21399_ (.A0(\design_top.core0.REG2[12][7] ),
    .A1(\design_top.core0.REG2[13][7] ),
    .A2(\design_top.core0.REG2[14][7] ),
    .A3(\design_top.core0.REG2[15][7] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21400_ (.A0(_03073_),
    .A1(_03074_),
    .A2(_03075_),
    .A3(_03076_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_03077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21401_ (.A0(\design_top.core0.REG2[0][8] ),
    .A1(\design_top.core0.REG2[1][8] ),
    .A2(\design_top.core0.REG2[2][8] ),
    .A3(\design_top.core0.REG2[3][8] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21402_ (.A0(\design_top.core0.REG2[4][8] ),
    .A1(\design_top.core0.REG2[5][8] ),
    .A2(\design_top.core0.REG2[6][8] ),
    .A3(\design_top.core0.REG2[7][8] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21403_ (.A0(\design_top.core0.REG2[8][8] ),
    .A1(\design_top.core0.REG2[9][8] ),
    .A2(\design_top.core0.REG2[10][8] ),
    .A3(\design_top.core0.REG2[11][8] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21404_ (.A0(\design_top.core0.REG2[12][8] ),
    .A1(\design_top.core0.REG2[13][8] ),
    .A2(\design_top.core0.REG2[14][8] ),
    .A3(\design_top.core0.REG2[15][8] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21405_ (.A0(_03066_),
    .A1(_03067_),
    .A2(_03068_),
    .A3(_03069_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_03070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21406_ (.A0(\design_top.core0.REG2[0][9] ),
    .A1(\design_top.core0.REG2[1][9] ),
    .A2(\design_top.core0.REG2[2][9] ),
    .A3(\design_top.core0.REG2[3][9] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21407_ (.A0(\design_top.core0.REG2[4][9] ),
    .A1(\design_top.core0.REG2[5][9] ),
    .A2(\design_top.core0.REG2[6][9] ),
    .A3(\design_top.core0.REG2[7][9] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21408_ (.A0(\design_top.core0.REG2[8][9] ),
    .A1(\design_top.core0.REG2[9][9] ),
    .A2(\design_top.core0.REG2[10][9] ),
    .A3(\design_top.core0.REG2[11][9] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21409_ (.A0(\design_top.core0.REG2[12][9] ),
    .A1(\design_top.core0.REG2[13][9] ),
    .A2(\design_top.core0.REG2[14][9] ),
    .A3(\design_top.core0.REG2[15][9] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21410_ (.A0(_03057_),
    .A1(_03058_),
    .A2(_03059_),
    .A3(_03060_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_03061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21411_ (.A0(\design_top.core0.REG2[0][10] ),
    .A1(\design_top.core0.REG2[1][10] ),
    .A2(\design_top.core0.REG2[2][10] ),
    .A3(\design_top.core0.REG2[3][10] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21412_ (.A0(\design_top.core0.REG2[4][10] ),
    .A1(\design_top.core0.REG2[5][10] ),
    .A2(\design_top.core0.REG2[6][10] ),
    .A3(\design_top.core0.REG2[7][10] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21413_ (.A0(\design_top.core0.REG2[8][10] ),
    .A1(\design_top.core0.REG2[9][10] ),
    .A2(\design_top.core0.REG2[10][10] ),
    .A3(\design_top.core0.REG2[11][10] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21414_ (.A0(\design_top.core0.REG2[12][10] ),
    .A1(\design_top.core0.REG2[13][10] ),
    .A2(\design_top.core0.REG2[14][10] ),
    .A3(\design_top.core0.REG2[15][10] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21415_ (.A0(_03050_),
    .A1(_03051_),
    .A2(_03052_),
    .A3(_03053_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_03054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21416_ (.A0(\design_top.core0.REG2[0][11] ),
    .A1(\design_top.core0.REG2[1][11] ),
    .A2(\design_top.core0.REG2[2][11] ),
    .A3(\design_top.core0.REG2[3][11] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21417_ (.A0(\design_top.core0.REG2[4][11] ),
    .A1(\design_top.core0.REG2[5][11] ),
    .A2(\design_top.core0.REG2[6][11] ),
    .A3(\design_top.core0.REG2[7][11] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21418_ (.A0(\design_top.core0.REG2[8][11] ),
    .A1(\design_top.core0.REG2[9][11] ),
    .A2(\design_top.core0.REG2[10][11] ),
    .A3(\design_top.core0.REG2[11][11] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21419_ (.A0(\design_top.core0.REG2[12][11] ),
    .A1(\design_top.core0.REG2[13][11] ),
    .A2(\design_top.core0.REG2[14][11] ),
    .A3(\design_top.core0.REG2[15][11] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21420_ (.A0(_03041_),
    .A1(_03042_),
    .A2(_03043_),
    .A3(_03044_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_03045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21421_ (.A0(\design_top.core0.REG2[0][12] ),
    .A1(\design_top.core0.REG2[1][12] ),
    .A2(\design_top.core0.REG2[2][12] ),
    .A3(\design_top.core0.REG2[3][12] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21422_ (.A0(\design_top.core0.REG2[4][12] ),
    .A1(\design_top.core0.REG2[5][12] ),
    .A2(\design_top.core0.REG2[6][12] ),
    .A3(\design_top.core0.REG2[7][12] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21423_ (.A0(\design_top.core0.REG2[8][12] ),
    .A1(\design_top.core0.REG2[9][12] ),
    .A2(\design_top.core0.REG2[10][12] ),
    .A3(\design_top.core0.REG2[11][12] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21424_ (.A0(\design_top.core0.REG2[12][12] ),
    .A1(\design_top.core0.REG2[13][12] ),
    .A2(\design_top.core0.REG2[14][12] ),
    .A3(\design_top.core0.REG2[15][12] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21425_ (.A0(_03034_),
    .A1(_03035_),
    .A2(_03036_),
    .A3(_03037_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_03038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21426_ (.A0(\design_top.core0.REG2[0][13] ),
    .A1(\design_top.core0.REG2[1][13] ),
    .A2(\design_top.core0.REG2[2][13] ),
    .A3(\design_top.core0.REG2[3][13] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21427_ (.A0(\design_top.core0.REG2[4][13] ),
    .A1(\design_top.core0.REG2[5][13] ),
    .A2(\design_top.core0.REG2[6][13] ),
    .A3(\design_top.core0.REG2[7][13] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21428_ (.A0(\design_top.core0.REG2[8][13] ),
    .A1(\design_top.core0.REG2[9][13] ),
    .A2(\design_top.core0.REG2[10][13] ),
    .A3(\design_top.core0.REG2[11][13] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21429_ (.A0(\design_top.core0.REG2[12][13] ),
    .A1(\design_top.core0.REG2[13][13] ),
    .A2(\design_top.core0.REG2[14][13] ),
    .A3(\design_top.core0.REG2[15][13] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21430_ (.A0(_03025_),
    .A1(_03026_),
    .A2(_03027_),
    .A3(_03028_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_03029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21431_ (.A0(\design_top.core0.REG2[0][14] ),
    .A1(\design_top.core0.REG2[1][14] ),
    .A2(\design_top.core0.REG2[2][14] ),
    .A3(\design_top.core0.REG2[3][14] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21432_ (.A0(\design_top.core0.REG2[4][14] ),
    .A1(\design_top.core0.REG2[5][14] ),
    .A2(\design_top.core0.REG2[6][14] ),
    .A3(\design_top.core0.REG2[7][14] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21433_ (.A0(\design_top.core0.REG2[8][14] ),
    .A1(\design_top.core0.REG2[9][14] ),
    .A2(\design_top.core0.REG2[10][14] ),
    .A3(\design_top.core0.REG2[11][14] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21434_ (.A0(\design_top.core0.REG2[12][14] ),
    .A1(\design_top.core0.REG2[13][14] ),
    .A2(\design_top.core0.REG2[14][14] ),
    .A3(\design_top.core0.REG2[15][14] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21435_ (.A0(_03017_),
    .A1(_03018_),
    .A2(_03019_),
    .A3(_03020_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_03021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21436_ (.A0(\design_top.core0.REG2[0][15] ),
    .A1(\design_top.core0.REG2[1][15] ),
    .A2(\design_top.core0.REG2[2][15] ),
    .A3(\design_top.core0.REG2[3][15] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21437_ (.A0(\design_top.core0.REG2[4][15] ),
    .A1(\design_top.core0.REG2[5][15] ),
    .A2(\design_top.core0.REG2[6][15] ),
    .A3(\design_top.core0.REG2[7][15] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21438_ (.A0(\design_top.core0.REG2[8][15] ),
    .A1(\design_top.core0.REG2[9][15] ),
    .A2(\design_top.core0.REG2[10][15] ),
    .A3(\design_top.core0.REG2[11][15] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21439_ (.A0(\design_top.core0.REG2[12][15] ),
    .A1(\design_top.core0.REG2[13][15] ),
    .A2(\design_top.core0.REG2[14][15] ),
    .A3(\design_top.core0.REG2[15][15] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21440_ (.A0(_03008_),
    .A1(_03009_),
    .A2(_03010_),
    .A3(_03011_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_03012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21441_ (.A0(\design_top.core0.REG2[0][16] ),
    .A1(\design_top.core0.REG2[1][16] ),
    .A2(\design_top.core0.REG2[2][16] ),
    .A3(\design_top.core0.REG2[3][16] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21442_ (.A0(\design_top.core0.REG2[4][16] ),
    .A1(\design_top.core0.REG2[5][16] ),
    .A2(\design_top.core0.REG2[6][16] ),
    .A3(\design_top.core0.REG2[7][16] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21443_ (.A0(\design_top.core0.REG2[8][16] ),
    .A1(\design_top.core0.REG2[9][16] ),
    .A2(\design_top.core0.REG2[10][16] ),
    .A3(\design_top.core0.REG2[11][16] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21444_ (.A0(\design_top.core0.REG2[12][16] ),
    .A1(\design_top.core0.REG2[13][16] ),
    .A2(\design_top.core0.REG2[14][16] ),
    .A3(\design_top.core0.REG2[15][16] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_03003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21445_ (.A0(_03000_),
    .A1(_03001_),
    .A2(_03002_),
    .A3(_03003_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_03004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21446_ (.A0(\design_top.core0.REG2[0][17] ),
    .A1(\design_top.core0.REG2[1][17] ),
    .A2(\design_top.core0.REG2[2][17] ),
    .A3(\design_top.core0.REG2[3][17] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21447_ (.A0(\design_top.core0.REG2[4][17] ),
    .A1(\design_top.core0.REG2[5][17] ),
    .A2(\design_top.core0.REG2[6][17] ),
    .A3(\design_top.core0.REG2[7][17] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21448_ (.A0(\design_top.core0.REG2[8][17] ),
    .A1(\design_top.core0.REG2[9][17] ),
    .A2(\design_top.core0.REG2[10][17] ),
    .A3(\design_top.core0.REG2[11][17] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21449_ (.A0(\design_top.core0.REG2[12][17] ),
    .A1(\design_top.core0.REG2[13][17] ),
    .A2(\design_top.core0.REG2[14][17] ),
    .A3(\design_top.core0.REG2[15][17] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21450_ (.A0(_02991_),
    .A1(_02992_),
    .A2(_02993_),
    .A3(_02994_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_02995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21451_ (.A0(\design_top.core0.REG2[0][18] ),
    .A1(\design_top.core0.REG2[1][18] ),
    .A2(\design_top.core0.REG2[2][18] ),
    .A3(\design_top.core0.REG2[3][18] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21452_ (.A0(\design_top.core0.REG2[4][18] ),
    .A1(\design_top.core0.REG2[5][18] ),
    .A2(\design_top.core0.REG2[6][18] ),
    .A3(\design_top.core0.REG2[7][18] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21453_ (.A0(\design_top.core0.REG2[8][18] ),
    .A1(\design_top.core0.REG2[9][18] ),
    .A2(\design_top.core0.REG2[10][18] ),
    .A3(\design_top.core0.REG2[11][18] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21454_ (.A0(\design_top.core0.REG2[12][18] ),
    .A1(\design_top.core0.REG2[13][18] ),
    .A2(\design_top.core0.REG2[14][18] ),
    .A3(\design_top.core0.REG2[15][18] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21455_ (.A0(_02983_),
    .A1(_02984_),
    .A2(_02985_),
    .A3(_02986_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_02987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21456_ (.A0(\design_top.core0.REG2[0][19] ),
    .A1(\design_top.core0.REG2[1][19] ),
    .A2(\design_top.core0.REG2[2][19] ),
    .A3(\design_top.core0.REG2[3][19] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21457_ (.A0(\design_top.core0.REG2[4][19] ),
    .A1(\design_top.core0.REG2[5][19] ),
    .A2(\design_top.core0.REG2[6][19] ),
    .A3(\design_top.core0.REG2[7][19] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21458_ (.A0(\design_top.core0.REG2[8][19] ),
    .A1(\design_top.core0.REG2[9][19] ),
    .A2(\design_top.core0.REG2[10][19] ),
    .A3(\design_top.core0.REG2[11][19] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21459_ (.A0(\design_top.core0.REG2[12][19] ),
    .A1(\design_top.core0.REG2[13][19] ),
    .A2(\design_top.core0.REG2[14][19] ),
    .A3(\design_top.core0.REG2[15][19] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21460_ (.A0(_02974_),
    .A1(_02975_),
    .A2(_02976_),
    .A3(_02977_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_02978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21461_ (.A0(\design_top.core0.REG2[0][20] ),
    .A1(\design_top.core0.REG2[1][20] ),
    .A2(\design_top.core0.REG2[2][20] ),
    .A3(\design_top.core0.REG2[3][20] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21462_ (.A0(\design_top.core0.REG2[4][20] ),
    .A1(\design_top.core0.REG2[5][20] ),
    .A2(\design_top.core0.REG2[6][20] ),
    .A3(\design_top.core0.REG2[7][20] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21463_ (.A0(\design_top.core0.REG2[8][20] ),
    .A1(\design_top.core0.REG2[9][20] ),
    .A2(\design_top.core0.REG2[10][20] ),
    .A3(\design_top.core0.REG2[11][20] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21464_ (.A0(\design_top.core0.REG2[12][20] ),
    .A1(\design_top.core0.REG2[13][20] ),
    .A2(\design_top.core0.REG2[14][20] ),
    .A3(\design_top.core0.REG2[15][20] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21465_ (.A0(_02966_),
    .A1(_02967_),
    .A2(_02968_),
    .A3(_02969_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_02970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21466_ (.A0(\design_top.core0.REG2[0][21] ),
    .A1(\design_top.core0.REG2[1][21] ),
    .A2(\design_top.core0.REG2[2][21] ),
    .A3(\design_top.core0.REG2[3][21] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21467_ (.A0(\design_top.core0.REG2[4][21] ),
    .A1(\design_top.core0.REG2[5][21] ),
    .A2(\design_top.core0.REG2[6][21] ),
    .A3(\design_top.core0.REG2[7][21] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21468_ (.A0(\design_top.core0.REG2[8][21] ),
    .A1(\design_top.core0.REG2[9][21] ),
    .A2(\design_top.core0.REG2[10][21] ),
    .A3(\design_top.core0.REG2[11][21] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21469_ (.A0(\design_top.core0.REG2[12][21] ),
    .A1(\design_top.core0.REG2[13][21] ),
    .A2(\design_top.core0.REG2[14][21] ),
    .A3(\design_top.core0.REG2[15][21] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21470_ (.A0(_02957_),
    .A1(_02958_),
    .A2(_02959_),
    .A3(_02960_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_02961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21471_ (.A0(\design_top.core0.REG2[0][22] ),
    .A1(\design_top.core0.REG2[1][22] ),
    .A2(\design_top.core0.REG2[2][22] ),
    .A3(\design_top.core0.REG2[3][22] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21472_ (.A0(\design_top.core0.REG2[4][22] ),
    .A1(\design_top.core0.REG2[5][22] ),
    .A2(\design_top.core0.REG2[6][22] ),
    .A3(\design_top.core0.REG2[7][22] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21473_ (.A0(\design_top.core0.REG2[8][22] ),
    .A1(\design_top.core0.REG2[9][22] ),
    .A2(\design_top.core0.REG2[10][22] ),
    .A3(\design_top.core0.REG2[11][22] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21474_ (.A0(\design_top.core0.REG2[12][22] ),
    .A1(\design_top.core0.REG2[13][22] ),
    .A2(\design_top.core0.REG2[14][22] ),
    .A3(\design_top.core0.REG2[15][22] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21475_ (.A0(_02949_),
    .A1(_02950_),
    .A2(_02951_),
    .A3(_02952_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_02953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21476_ (.A0(\design_top.core0.REG2[0][23] ),
    .A1(\design_top.core0.REG2[1][23] ),
    .A2(\design_top.core0.REG2[2][23] ),
    .A3(\design_top.core0.REG2[3][23] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21477_ (.A0(\design_top.core0.REG2[4][23] ),
    .A1(\design_top.core0.REG2[5][23] ),
    .A2(\design_top.core0.REG2[6][23] ),
    .A3(\design_top.core0.REG2[7][23] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21478_ (.A0(\design_top.core0.REG2[8][23] ),
    .A1(\design_top.core0.REG2[9][23] ),
    .A2(\design_top.core0.REG2[10][23] ),
    .A3(\design_top.core0.REG2[11][23] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21479_ (.A0(\design_top.core0.REG2[12][23] ),
    .A1(\design_top.core0.REG2[13][23] ),
    .A2(\design_top.core0.REG2[14][23] ),
    .A3(\design_top.core0.REG2[15][23] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21480_ (.A0(_02940_),
    .A1(_02941_),
    .A2(_02942_),
    .A3(_02943_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_02944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21481_ (.A0(\design_top.core0.REG2[0][24] ),
    .A1(\design_top.core0.REG2[1][24] ),
    .A2(\design_top.core0.REG2[2][24] ),
    .A3(\design_top.core0.REG2[3][24] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21482_ (.A0(\design_top.core0.REG2[4][24] ),
    .A1(\design_top.core0.REG2[5][24] ),
    .A2(\design_top.core0.REG2[6][24] ),
    .A3(\design_top.core0.REG2[7][24] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21483_ (.A0(\design_top.core0.REG2[8][24] ),
    .A1(\design_top.core0.REG2[9][24] ),
    .A2(\design_top.core0.REG2[10][24] ),
    .A3(\design_top.core0.REG2[11][24] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21484_ (.A0(\design_top.core0.REG2[12][24] ),
    .A1(\design_top.core0.REG2[13][24] ),
    .A2(\design_top.core0.REG2[14][24] ),
    .A3(\design_top.core0.REG2[15][24] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21485_ (.A0(_02932_),
    .A1(_02933_),
    .A2(_02934_),
    .A3(_02935_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_02936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21486_ (.A0(\design_top.core0.REG2[0][25] ),
    .A1(\design_top.core0.REG2[1][25] ),
    .A2(\design_top.core0.REG2[2][25] ),
    .A3(\design_top.core0.REG2[3][25] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21487_ (.A0(\design_top.core0.REG2[4][25] ),
    .A1(\design_top.core0.REG2[5][25] ),
    .A2(\design_top.core0.REG2[6][25] ),
    .A3(\design_top.core0.REG2[7][25] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21488_ (.A0(\design_top.core0.REG2[8][25] ),
    .A1(\design_top.core0.REG2[9][25] ),
    .A2(\design_top.core0.REG2[10][25] ),
    .A3(\design_top.core0.REG2[11][25] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21489_ (.A0(\design_top.core0.REG2[12][25] ),
    .A1(\design_top.core0.REG2[13][25] ),
    .A2(\design_top.core0.REG2[14][25] ),
    .A3(\design_top.core0.REG2[15][25] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21490_ (.A0(_02923_),
    .A1(_02924_),
    .A2(_02925_),
    .A3(_02926_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_02927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21491_ (.A0(\design_top.core0.REG2[0][26] ),
    .A1(\design_top.core0.REG2[1][26] ),
    .A2(\design_top.core0.REG2[2][26] ),
    .A3(\design_top.core0.REG2[3][26] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21492_ (.A0(\design_top.core0.REG2[4][26] ),
    .A1(\design_top.core0.REG2[5][26] ),
    .A2(\design_top.core0.REG2[6][26] ),
    .A3(\design_top.core0.REG2[7][26] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21493_ (.A0(\design_top.core0.REG2[8][26] ),
    .A1(\design_top.core0.REG2[9][26] ),
    .A2(\design_top.core0.REG2[10][26] ),
    .A3(\design_top.core0.REG2[11][26] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21494_ (.A0(\design_top.core0.REG2[12][26] ),
    .A1(\design_top.core0.REG2[13][26] ),
    .A2(\design_top.core0.REG2[14][26] ),
    .A3(\design_top.core0.REG2[15][26] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21495_ (.A0(_02915_),
    .A1(_02916_),
    .A2(_02917_),
    .A3(_02918_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_02919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21496_ (.A0(\design_top.core0.REG2[0][27] ),
    .A1(\design_top.core0.REG2[1][27] ),
    .A2(\design_top.core0.REG2[2][27] ),
    .A3(\design_top.core0.REG2[3][27] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21497_ (.A0(\design_top.core0.REG2[4][27] ),
    .A1(\design_top.core0.REG2[5][27] ),
    .A2(\design_top.core0.REG2[6][27] ),
    .A3(\design_top.core0.REG2[7][27] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21498_ (.A0(\design_top.core0.REG2[8][27] ),
    .A1(\design_top.core0.REG2[9][27] ),
    .A2(\design_top.core0.REG2[10][27] ),
    .A3(\design_top.core0.REG2[11][27] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21499_ (.A0(\design_top.core0.REG2[12][27] ),
    .A1(\design_top.core0.REG2[13][27] ),
    .A2(\design_top.core0.REG2[14][27] ),
    .A3(\design_top.core0.REG2[15][27] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21500_ (.A0(_02906_),
    .A1(_02907_),
    .A2(_02908_),
    .A3(_02909_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_02910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21501_ (.A0(\design_top.core0.REG2[0][28] ),
    .A1(\design_top.core0.REG2[1][28] ),
    .A2(\design_top.core0.REG2[2][28] ),
    .A3(\design_top.core0.REG2[3][28] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21502_ (.A0(\design_top.core0.REG2[4][28] ),
    .A1(\design_top.core0.REG2[5][28] ),
    .A2(\design_top.core0.REG2[6][28] ),
    .A3(\design_top.core0.REG2[7][28] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21503_ (.A0(\design_top.core0.REG2[8][28] ),
    .A1(\design_top.core0.REG2[9][28] ),
    .A2(\design_top.core0.REG2[10][28] ),
    .A3(\design_top.core0.REG2[11][28] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21504_ (.A0(\design_top.core0.REG2[12][28] ),
    .A1(\design_top.core0.REG2[13][28] ),
    .A2(\design_top.core0.REG2[14][28] ),
    .A3(\design_top.core0.REG2[15][28] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21505_ (.A0(_02898_),
    .A1(_02899_),
    .A2(_02900_),
    .A3(_02901_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_02902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21506_ (.A0(\design_top.core0.REG2[0][29] ),
    .A1(\design_top.core0.REG2[1][29] ),
    .A2(\design_top.core0.REG2[2][29] ),
    .A3(\design_top.core0.REG2[3][29] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21507_ (.A0(\design_top.core0.REG2[4][29] ),
    .A1(\design_top.core0.REG2[5][29] ),
    .A2(\design_top.core0.REG2[6][29] ),
    .A3(\design_top.core0.REG2[7][29] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21508_ (.A0(\design_top.core0.REG2[8][29] ),
    .A1(\design_top.core0.REG2[9][29] ),
    .A2(\design_top.core0.REG2[10][29] ),
    .A3(\design_top.core0.REG2[11][29] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21509_ (.A0(\design_top.core0.REG2[12][29] ),
    .A1(\design_top.core0.REG2[13][29] ),
    .A2(\design_top.core0.REG2[14][29] ),
    .A3(\design_top.core0.REG2[15][29] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21510_ (.A0(_02889_),
    .A1(_02890_),
    .A2(_02891_),
    .A3(_02892_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_02893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21511_ (.A0(\design_top.core0.REG2[0][30] ),
    .A1(\design_top.core0.REG2[1][30] ),
    .A2(\design_top.core0.REG2[2][30] ),
    .A3(\design_top.core0.REG2[3][30] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21512_ (.A0(\design_top.core0.REG2[4][30] ),
    .A1(\design_top.core0.REG2[5][30] ),
    .A2(\design_top.core0.REG2[6][30] ),
    .A3(\design_top.core0.REG2[7][30] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21513_ (.A0(\design_top.core0.REG2[8][30] ),
    .A1(\design_top.core0.REG2[9][30] ),
    .A2(\design_top.core0.REG2[10][30] ),
    .A3(\design_top.core0.REG2[11][30] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21514_ (.A0(\design_top.core0.REG2[12][30] ),
    .A1(\design_top.core0.REG2[13][30] ),
    .A2(\design_top.core0.REG2[14][30] ),
    .A3(\design_top.core0.REG2[15][30] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21515_ (.A0(_02880_),
    .A1(_02881_),
    .A2(_02882_),
    .A3(_02883_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_02884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21516_ (.A0(\design_top.core0.REG2[0][31] ),
    .A1(\design_top.core0.REG2[1][31] ),
    .A2(\design_top.core0.REG2[2][31] ),
    .A3(\design_top.core0.REG2[3][31] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21517_ (.A0(\design_top.core0.REG2[4][31] ),
    .A1(\design_top.core0.REG2[5][31] ),
    .A2(\design_top.core0.REG2[6][31] ),
    .A3(\design_top.core0.REG2[7][31] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21518_ (.A0(\design_top.core0.REG2[8][31] ),
    .A1(\design_top.core0.REG2[9][31] ),
    .A2(\design_top.core0.REG2[10][31] ),
    .A3(\design_top.core0.REG2[11][31] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21519_ (.A0(\design_top.core0.REG2[12][31] ),
    .A1(\design_top.core0.REG2[13][31] ),
    .A2(\design_top.core0.REG2[14][31] ),
    .A3(\design_top.core0.REG2[15][31] ),
    .S0(_00689_),
    .S1(_00690_),
    .X(_02874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21520_ (.A0(_02871_),
    .A1(_02872_),
    .A2(_02873_),
    .A3(_02874_),
    .S0(_00691_),
    .S1(_00692_),
    .X(_02875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21521_ (.A0(\design_top.core0.REG1[0][4] ),
    .A1(\design_top.core0.REG1[1][4] ),
    .A2(\design_top.core0.REG1[2][4] ),
    .A3(\design_top.core0.REG1[3][4] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21522_ (.A0(\design_top.core0.REG1[4][4] ),
    .A1(\design_top.core0.REG1[5][4] ),
    .A2(\design_top.core0.REG1[6][4] ),
    .A3(\design_top.core0.REG1[7][4] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21523_ (.A0(\design_top.core0.REG1[8][4] ),
    .A1(\design_top.core0.REG1[9][4] ),
    .A2(\design_top.core0.REG1[10][4] ),
    .A3(\design_top.core0.REG1[11][4] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21524_ (.A0(\design_top.core0.REG1[12][4] ),
    .A1(\design_top.core0.REG1[13][4] ),
    .A2(\design_top.core0.REG1[14][4] ),
    .A3(\design_top.core0.REG1[15][4] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21525_ (.A0(_02841_),
    .A1(_02842_),
    .A2(_02843_),
    .A3(_02844_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21526_ (.A0(\design_top.core0.REG1[0][5] ),
    .A1(\design_top.core0.REG1[1][5] ),
    .A2(\design_top.core0.REG1[2][5] ),
    .A3(\design_top.core0.REG1[3][5] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21527_ (.A0(\design_top.core0.REG1[4][5] ),
    .A1(\design_top.core0.REG1[5][5] ),
    .A2(\design_top.core0.REG1[6][5] ),
    .A3(\design_top.core0.REG1[7][5] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21528_ (.A0(\design_top.core0.REG1[8][5] ),
    .A1(\design_top.core0.REG1[9][5] ),
    .A2(\design_top.core0.REG1[10][5] ),
    .A3(\design_top.core0.REG1[11][5] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21529_ (.A0(\design_top.core0.REG1[12][5] ),
    .A1(\design_top.core0.REG1[13][5] ),
    .A2(\design_top.core0.REG1[14][5] ),
    .A3(\design_top.core0.REG1[15][5] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21530_ (.A0(_02835_),
    .A1(_02836_),
    .A2(_02837_),
    .A3(_02838_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21531_ (.A0(\design_top.core0.REG1[0][6] ),
    .A1(\design_top.core0.REG1[1][6] ),
    .A2(\design_top.core0.REG1[2][6] ),
    .A3(\design_top.core0.REG1[3][6] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21532_ (.A0(\design_top.core0.REG1[4][6] ),
    .A1(\design_top.core0.REG1[5][6] ),
    .A2(\design_top.core0.REG1[6][6] ),
    .A3(\design_top.core0.REG1[7][6] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21533_ (.A0(\design_top.core0.REG1[8][6] ),
    .A1(\design_top.core0.REG1[9][6] ),
    .A2(\design_top.core0.REG1[10][6] ),
    .A3(\design_top.core0.REG1[11][6] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21534_ (.A0(\design_top.core0.REG1[12][6] ),
    .A1(\design_top.core0.REG1[13][6] ),
    .A2(\design_top.core0.REG1[14][6] ),
    .A3(\design_top.core0.REG1[15][6] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21535_ (.A0(_02829_),
    .A1(_02830_),
    .A2(_02831_),
    .A3(_02832_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21536_ (.A0(\design_top.core0.REG1[0][7] ),
    .A1(\design_top.core0.REG1[1][7] ),
    .A2(\design_top.core0.REG1[2][7] ),
    .A3(\design_top.core0.REG1[3][7] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21537_ (.A0(\design_top.core0.REG1[4][7] ),
    .A1(\design_top.core0.REG1[5][7] ),
    .A2(\design_top.core0.REG1[6][7] ),
    .A3(\design_top.core0.REG1[7][7] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21538_ (.A0(\design_top.core0.REG1[8][7] ),
    .A1(\design_top.core0.REG1[9][7] ),
    .A2(\design_top.core0.REG1[10][7] ),
    .A3(\design_top.core0.REG1[11][7] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21539_ (.A0(\design_top.core0.REG1[12][7] ),
    .A1(\design_top.core0.REG1[13][7] ),
    .A2(\design_top.core0.REG1[14][7] ),
    .A3(\design_top.core0.REG1[15][7] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21540_ (.A0(_02823_),
    .A1(_02824_),
    .A2(_02825_),
    .A3(_02826_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21541_ (.A0(\design_top.core0.REG1[0][8] ),
    .A1(\design_top.core0.REG1[1][8] ),
    .A2(\design_top.core0.REG1[2][8] ),
    .A3(\design_top.core0.REG1[3][8] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21542_ (.A0(\design_top.core0.REG1[4][8] ),
    .A1(\design_top.core0.REG1[5][8] ),
    .A2(\design_top.core0.REG1[6][8] ),
    .A3(\design_top.core0.REG1[7][8] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21543_ (.A0(\design_top.core0.REG1[8][8] ),
    .A1(\design_top.core0.REG1[9][8] ),
    .A2(\design_top.core0.REG1[10][8] ),
    .A3(\design_top.core0.REG1[11][8] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21544_ (.A0(\design_top.core0.REG1[12][8] ),
    .A1(\design_top.core0.REG1[13][8] ),
    .A2(\design_top.core0.REG1[14][8] ),
    .A3(\design_top.core0.REG1[15][8] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21545_ (.A0(_02817_),
    .A1(_02818_),
    .A2(_02819_),
    .A3(_02820_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21546_ (.A0(\design_top.core0.REG1[0][9] ),
    .A1(\design_top.core0.REG1[1][9] ),
    .A2(\design_top.core0.REG1[2][9] ),
    .A3(\design_top.core0.REG1[3][9] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21547_ (.A0(\design_top.core0.REG1[4][9] ),
    .A1(\design_top.core0.REG1[5][9] ),
    .A2(\design_top.core0.REG1[6][9] ),
    .A3(\design_top.core0.REG1[7][9] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21548_ (.A0(\design_top.core0.REG1[8][9] ),
    .A1(\design_top.core0.REG1[9][9] ),
    .A2(\design_top.core0.REG1[10][9] ),
    .A3(\design_top.core0.REG1[11][9] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21549_ (.A0(\design_top.core0.REG1[12][9] ),
    .A1(\design_top.core0.REG1[13][9] ),
    .A2(\design_top.core0.REG1[14][9] ),
    .A3(\design_top.core0.REG1[15][9] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21550_ (.A0(_02811_),
    .A1(_02812_),
    .A2(_02813_),
    .A3(_02814_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21551_ (.A0(\design_top.core0.REG1[0][10] ),
    .A1(\design_top.core0.REG1[1][10] ),
    .A2(\design_top.core0.REG1[2][10] ),
    .A3(\design_top.core0.REG1[3][10] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21552_ (.A0(\design_top.core0.REG1[4][10] ),
    .A1(\design_top.core0.REG1[5][10] ),
    .A2(\design_top.core0.REG1[6][10] ),
    .A3(\design_top.core0.REG1[7][10] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21553_ (.A0(\design_top.core0.REG1[8][10] ),
    .A1(\design_top.core0.REG1[9][10] ),
    .A2(\design_top.core0.REG1[10][10] ),
    .A3(\design_top.core0.REG1[11][10] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21554_ (.A0(\design_top.core0.REG1[12][10] ),
    .A1(\design_top.core0.REG1[13][10] ),
    .A2(\design_top.core0.REG1[14][10] ),
    .A3(\design_top.core0.REG1[15][10] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21555_ (.A0(_02805_),
    .A1(_02806_),
    .A2(_02807_),
    .A3(_02808_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21556_ (.A0(\design_top.core0.REG1[0][11] ),
    .A1(\design_top.core0.REG1[1][11] ),
    .A2(\design_top.core0.REG1[2][11] ),
    .A3(\design_top.core0.REG1[3][11] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21557_ (.A0(\design_top.core0.REG1[4][11] ),
    .A1(\design_top.core0.REG1[5][11] ),
    .A2(\design_top.core0.REG1[6][11] ),
    .A3(\design_top.core0.REG1[7][11] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21558_ (.A0(\design_top.core0.REG1[8][11] ),
    .A1(\design_top.core0.REG1[9][11] ),
    .A2(\design_top.core0.REG1[10][11] ),
    .A3(\design_top.core0.REG1[11][11] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21559_ (.A0(\design_top.core0.REG1[12][11] ),
    .A1(\design_top.core0.REG1[13][11] ),
    .A2(\design_top.core0.REG1[14][11] ),
    .A3(\design_top.core0.REG1[15][11] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21560_ (.A0(_02799_),
    .A1(_02800_),
    .A2(_02801_),
    .A3(_02802_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21561_ (.A0(\design_top.core0.REG1[0][12] ),
    .A1(\design_top.core0.REG1[1][12] ),
    .A2(\design_top.core0.REG1[2][12] ),
    .A3(\design_top.core0.REG1[3][12] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21562_ (.A0(\design_top.core0.REG1[4][12] ),
    .A1(\design_top.core0.REG1[5][12] ),
    .A2(\design_top.core0.REG1[6][12] ),
    .A3(\design_top.core0.REG1[7][12] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21563_ (.A0(\design_top.core0.REG1[8][12] ),
    .A1(\design_top.core0.REG1[9][12] ),
    .A2(\design_top.core0.REG1[10][12] ),
    .A3(\design_top.core0.REG1[11][12] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21564_ (.A0(\design_top.core0.REG1[12][12] ),
    .A1(\design_top.core0.REG1[13][12] ),
    .A2(\design_top.core0.REG1[14][12] ),
    .A3(\design_top.core0.REG1[15][12] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21565_ (.A0(_02793_),
    .A1(_02794_),
    .A2(_02795_),
    .A3(_02796_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21566_ (.A0(\design_top.core0.REG1[0][13] ),
    .A1(\design_top.core0.REG1[1][13] ),
    .A2(\design_top.core0.REG1[2][13] ),
    .A3(\design_top.core0.REG1[3][13] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21567_ (.A0(\design_top.core0.REG1[4][13] ),
    .A1(\design_top.core0.REG1[5][13] ),
    .A2(\design_top.core0.REG1[6][13] ),
    .A3(\design_top.core0.REG1[7][13] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21568_ (.A0(\design_top.core0.REG1[8][13] ),
    .A1(\design_top.core0.REG1[9][13] ),
    .A2(\design_top.core0.REG1[10][13] ),
    .A3(\design_top.core0.REG1[11][13] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21569_ (.A0(\design_top.core0.REG1[12][13] ),
    .A1(\design_top.core0.REG1[13][13] ),
    .A2(\design_top.core0.REG1[14][13] ),
    .A3(\design_top.core0.REG1[15][13] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21570_ (.A0(_02787_),
    .A1(_02788_),
    .A2(_02789_),
    .A3(_02790_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21571_ (.A0(\design_top.core0.REG1[0][14] ),
    .A1(\design_top.core0.REG1[1][14] ),
    .A2(\design_top.core0.REG1[2][14] ),
    .A3(\design_top.core0.REG1[3][14] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21572_ (.A0(\design_top.core0.REG1[4][14] ),
    .A1(\design_top.core0.REG1[5][14] ),
    .A2(\design_top.core0.REG1[6][14] ),
    .A3(\design_top.core0.REG1[7][14] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21573_ (.A0(\design_top.core0.REG1[8][14] ),
    .A1(\design_top.core0.REG1[9][14] ),
    .A2(\design_top.core0.REG1[10][14] ),
    .A3(\design_top.core0.REG1[11][14] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21574_ (.A0(\design_top.core0.REG1[12][14] ),
    .A1(\design_top.core0.REG1[13][14] ),
    .A2(\design_top.core0.REG1[14][14] ),
    .A3(\design_top.core0.REG1[15][14] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21575_ (.A0(_02781_),
    .A1(_02782_),
    .A2(_02783_),
    .A3(_02784_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21576_ (.A0(\design_top.core0.REG1[0][15] ),
    .A1(\design_top.core0.REG1[1][15] ),
    .A2(\design_top.core0.REG1[2][15] ),
    .A3(\design_top.core0.REG1[3][15] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21577_ (.A0(\design_top.core0.REG1[4][15] ),
    .A1(\design_top.core0.REG1[5][15] ),
    .A2(\design_top.core0.REG1[6][15] ),
    .A3(\design_top.core0.REG1[7][15] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21578_ (.A0(\design_top.core0.REG1[8][15] ),
    .A1(\design_top.core0.REG1[9][15] ),
    .A2(\design_top.core0.REG1[10][15] ),
    .A3(\design_top.core0.REG1[11][15] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21579_ (.A0(\design_top.core0.REG1[12][15] ),
    .A1(\design_top.core0.REG1[13][15] ),
    .A2(\design_top.core0.REG1[14][15] ),
    .A3(\design_top.core0.REG1[15][15] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21580_ (.A0(_02775_),
    .A1(_02776_),
    .A2(_02777_),
    .A3(_02778_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21581_ (.A0(\design_top.core0.REG1[0][16] ),
    .A1(\design_top.core0.REG1[1][16] ),
    .A2(\design_top.core0.REG1[2][16] ),
    .A3(\design_top.core0.REG1[3][16] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21582_ (.A0(\design_top.core0.REG1[4][16] ),
    .A1(\design_top.core0.REG1[5][16] ),
    .A2(\design_top.core0.REG1[6][16] ),
    .A3(\design_top.core0.REG1[7][16] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21583_ (.A0(\design_top.core0.REG1[8][16] ),
    .A1(\design_top.core0.REG1[9][16] ),
    .A2(\design_top.core0.REG1[10][16] ),
    .A3(\design_top.core0.REG1[11][16] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21584_ (.A0(\design_top.core0.REG1[12][16] ),
    .A1(\design_top.core0.REG1[13][16] ),
    .A2(\design_top.core0.REG1[14][16] ),
    .A3(\design_top.core0.REG1[15][16] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21585_ (.A0(_02769_),
    .A1(_02770_),
    .A2(_02771_),
    .A3(_02772_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21586_ (.A0(\design_top.core0.REG1[0][17] ),
    .A1(\design_top.core0.REG1[1][17] ),
    .A2(\design_top.core0.REG1[2][17] ),
    .A3(\design_top.core0.REG1[3][17] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21587_ (.A0(\design_top.core0.REG1[4][17] ),
    .A1(\design_top.core0.REG1[5][17] ),
    .A2(\design_top.core0.REG1[6][17] ),
    .A3(\design_top.core0.REG1[7][17] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21588_ (.A0(\design_top.core0.REG1[8][17] ),
    .A1(\design_top.core0.REG1[9][17] ),
    .A2(\design_top.core0.REG1[10][17] ),
    .A3(\design_top.core0.REG1[11][17] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21589_ (.A0(\design_top.core0.REG1[12][17] ),
    .A1(\design_top.core0.REG1[13][17] ),
    .A2(\design_top.core0.REG1[14][17] ),
    .A3(\design_top.core0.REG1[15][17] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21590_ (.A0(_02763_),
    .A1(_02764_),
    .A2(_02765_),
    .A3(_02766_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21591_ (.A0(\design_top.core0.REG1[0][18] ),
    .A1(\design_top.core0.REG1[1][18] ),
    .A2(\design_top.core0.REG1[2][18] ),
    .A3(\design_top.core0.REG1[3][18] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21592_ (.A0(\design_top.core0.REG1[4][18] ),
    .A1(\design_top.core0.REG1[5][18] ),
    .A2(\design_top.core0.REG1[6][18] ),
    .A3(\design_top.core0.REG1[7][18] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21593_ (.A0(\design_top.core0.REG1[8][18] ),
    .A1(\design_top.core0.REG1[9][18] ),
    .A2(\design_top.core0.REG1[10][18] ),
    .A3(\design_top.core0.REG1[11][18] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21594_ (.A0(\design_top.core0.REG1[12][18] ),
    .A1(\design_top.core0.REG1[13][18] ),
    .A2(\design_top.core0.REG1[14][18] ),
    .A3(\design_top.core0.REG1[15][18] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21595_ (.A0(_02757_),
    .A1(_02758_),
    .A2(_02759_),
    .A3(_02760_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21596_ (.A0(\design_top.core0.REG1[0][19] ),
    .A1(\design_top.core0.REG1[1][19] ),
    .A2(\design_top.core0.REG1[2][19] ),
    .A3(\design_top.core0.REG1[3][19] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21597_ (.A0(\design_top.core0.REG1[4][19] ),
    .A1(\design_top.core0.REG1[5][19] ),
    .A2(\design_top.core0.REG1[6][19] ),
    .A3(\design_top.core0.REG1[7][19] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21598_ (.A0(\design_top.core0.REG1[8][19] ),
    .A1(\design_top.core0.REG1[9][19] ),
    .A2(\design_top.core0.REG1[10][19] ),
    .A3(\design_top.core0.REG1[11][19] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21599_ (.A0(\design_top.core0.REG1[12][19] ),
    .A1(\design_top.core0.REG1[13][19] ),
    .A2(\design_top.core0.REG1[14][19] ),
    .A3(\design_top.core0.REG1[15][19] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21600_ (.A0(_02751_),
    .A1(_02752_),
    .A2(_02753_),
    .A3(_02754_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21601_ (.A0(\design_top.core0.REG1[0][20] ),
    .A1(\design_top.core0.REG1[1][20] ),
    .A2(\design_top.core0.REG1[2][20] ),
    .A3(\design_top.core0.REG1[3][20] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21602_ (.A0(\design_top.core0.REG1[4][20] ),
    .A1(\design_top.core0.REG1[5][20] ),
    .A2(\design_top.core0.REG1[6][20] ),
    .A3(\design_top.core0.REG1[7][20] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21603_ (.A0(\design_top.core0.REG1[8][20] ),
    .A1(\design_top.core0.REG1[9][20] ),
    .A2(\design_top.core0.REG1[10][20] ),
    .A3(\design_top.core0.REG1[11][20] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21604_ (.A0(\design_top.core0.REG1[12][20] ),
    .A1(\design_top.core0.REG1[13][20] ),
    .A2(\design_top.core0.REG1[14][20] ),
    .A3(\design_top.core0.REG1[15][20] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21605_ (.A0(_02745_),
    .A1(_02746_),
    .A2(_02747_),
    .A3(_02748_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21606_ (.A0(\design_top.core0.REG1[0][21] ),
    .A1(\design_top.core0.REG1[1][21] ),
    .A2(\design_top.core0.REG1[2][21] ),
    .A3(\design_top.core0.REG1[3][21] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21607_ (.A0(\design_top.core0.REG1[4][21] ),
    .A1(\design_top.core0.REG1[5][21] ),
    .A2(\design_top.core0.REG1[6][21] ),
    .A3(\design_top.core0.REG1[7][21] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21608_ (.A0(\design_top.core0.REG1[8][21] ),
    .A1(\design_top.core0.REG1[9][21] ),
    .A2(\design_top.core0.REG1[10][21] ),
    .A3(\design_top.core0.REG1[11][21] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21609_ (.A0(\design_top.core0.REG1[12][21] ),
    .A1(\design_top.core0.REG1[13][21] ),
    .A2(\design_top.core0.REG1[14][21] ),
    .A3(\design_top.core0.REG1[15][21] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21610_ (.A0(_02739_),
    .A1(_02740_),
    .A2(_02741_),
    .A3(_02742_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21611_ (.A0(\design_top.core0.REG1[0][22] ),
    .A1(\design_top.core0.REG1[1][22] ),
    .A2(\design_top.core0.REG1[2][22] ),
    .A3(\design_top.core0.REG1[3][22] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21612_ (.A0(\design_top.core0.REG1[4][22] ),
    .A1(\design_top.core0.REG1[5][22] ),
    .A2(\design_top.core0.REG1[6][22] ),
    .A3(\design_top.core0.REG1[7][22] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21613_ (.A0(\design_top.core0.REG1[8][22] ),
    .A1(\design_top.core0.REG1[9][22] ),
    .A2(\design_top.core0.REG1[10][22] ),
    .A3(\design_top.core0.REG1[11][22] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21614_ (.A0(\design_top.core0.REG1[12][22] ),
    .A1(\design_top.core0.REG1[13][22] ),
    .A2(\design_top.core0.REG1[14][22] ),
    .A3(\design_top.core0.REG1[15][22] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21615_ (.A0(_02733_),
    .A1(_02734_),
    .A2(_02735_),
    .A3(_02736_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21616_ (.A0(\design_top.core0.REG1[0][23] ),
    .A1(\design_top.core0.REG1[1][23] ),
    .A2(\design_top.core0.REG1[2][23] ),
    .A3(\design_top.core0.REG1[3][23] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21617_ (.A0(\design_top.core0.REG1[4][23] ),
    .A1(\design_top.core0.REG1[5][23] ),
    .A2(\design_top.core0.REG1[6][23] ),
    .A3(\design_top.core0.REG1[7][23] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21618_ (.A0(\design_top.core0.REG1[8][23] ),
    .A1(\design_top.core0.REG1[9][23] ),
    .A2(\design_top.core0.REG1[10][23] ),
    .A3(\design_top.core0.REG1[11][23] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21619_ (.A0(\design_top.core0.REG1[12][23] ),
    .A1(\design_top.core0.REG1[13][23] ),
    .A2(\design_top.core0.REG1[14][23] ),
    .A3(\design_top.core0.REG1[15][23] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21620_ (.A0(_02727_),
    .A1(_02728_),
    .A2(_02729_),
    .A3(_02730_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21621_ (.A0(\design_top.core0.REG1[0][24] ),
    .A1(\design_top.core0.REG1[1][24] ),
    .A2(\design_top.core0.REG1[2][24] ),
    .A3(\design_top.core0.REG1[3][24] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21622_ (.A0(\design_top.core0.REG1[4][24] ),
    .A1(\design_top.core0.REG1[5][24] ),
    .A2(\design_top.core0.REG1[6][24] ),
    .A3(\design_top.core0.REG1[7][24] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21623_ (.A0(\design_top.core0.REG1[8][24] ),
    .A1(\design_top.core0.REG1[9][24] ),
    .A2(\design_top.core0.REG1[10][24] ),
    .A3(\design_top.core0.REG1[11][24] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21624_ (.A0(\design_top.core0.REG1[12][24] ),
    .A1(\design_top.core0.REG1[13][24] ),
    .A2(\design_top.core0.REG1[14][24] ),
    .A3(\design_top.core0.REG1[15][24] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21625_ (.A0(_02721_),
    .A1(_02722_),
    .A2(_02723_),
    .A3(_02724_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21626_ (.A0(\design_top.core0.REG1[0][25] ),
    .A1(\design_top.core0.REG1[1][25] ),
    .A2(\design_top.core0.REG1[2][25] ),
    .A3(\design_top.core0.REG1[3][25] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21627_ (.A0(\design_top.core0.REG1[4][25] ),
    .A1(\design_top.core0.REG1[5][25] ),
    .A2(\design_top.core0.REG1[6][25] ),
    .A3(\design_top.core0.REG1[7][25] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21628_ (.A0(\design_top.core0.REG1[8][25] ),
    .A1(\design_top.core0.REG1[9][25] ),
    .A2(\design_top.core0.REG1[10][25] ),
    .A3(\design_top.core0.REG1[11][25] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21629_ (.A0(\design_top.core0.REG1[12][25] ),
    .A1(\design_top.core0.REG1[13][25] ),
    .A2(\design_top.core0.REG1[14][25] ),
    .A3(\design_top.core0.REG1[15][25] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21630_ (.A0(_02715_),
    .A1(_02716_),
    .A2(_02717_),
    .A3(_02718_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21631_ (.A0(\design_top.core0.REG1[0][26] ),
    .A1(\design_top.core0.REG1[1][26] ),
    .A2(\design_top.core0.REG1[2][26] ),
    .A3(\design_top.core0.REG1[3][26] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21632_ (.A0(\design_top.core0.REG1[4][26] ),
    .A1(\design_top.core0.REG1[5][26] ),
    .A2(\design_top.core0.REG1[6][26] ),
    .A3(\design_top.core0.REG1[7][26] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21633_ (.A0(\design_top.core0.REG1[8][26] ),
    .A1(\design_top.core0.REG1[9][26] ),
    .A2(\design_top.core0.REG1[10][26] ),
    .A3(\design_top.core0.REG1[11][26] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21634_ (.A0(\design_top.core0.REG1[12][26] ),
    .A1(\design_top.core0.REG1[13][26] ),
    .A2(\design_top.core0.REG1[14][26] ),
    .A3(\design_top.core0.REG1[15][26] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21635_ (.A0(_02709_),
    .A1(_02710_),
    .A2(_02711_),
    .A3(_02712_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21636_ (.A0(\design_top.core0.REG1[0][27] ),
    .A1(\design_top.core0.REG1[1][27] ),
    .A2(\design_top.core0.REG1[2][27] ),
    .A3(\design_top.core0.REG1[3][27] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21637_ (.A0(\design_top.core0.REG1[4][27] ),
    .A1(\design_top.core0.REG1[5][27] ),
    .A2(\design_top.core0.REG1[6][27] ),
    .A3(\design_top.core0.REG1[7][27] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21638_ (.A0(\design_top.core0.REG1[8][27] ),
    .A1(\design_top.core0.REG1[9][27] ),
    .A2(\design_top.core0.REG1[10][27] ),
    .A3(\design_top.core0.REG1[11][27] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21639_ (.A0(\design_top.core0.REG1[12][27] ),
    .A1(\design_top.core0.REG1[13][27] ),
    .A2(\design_top.core0.REG1[14][27] ),
    .A3(\design_top.core0.REG1[15][27] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21640_ (.A0(_02703_),
    .A1(_02704_),
    .A2(_02705_),
    .A3(_02706_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21641_ (.A0(\design_top.core0.REG1[0][28] ),
    .A1(\design_top.core0.REG1[1][28] ),
    .A2(\design_top.core0.REG1[2][28] ),
    .A3(\design_top.core0.REG1[3][28] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21642_ (.A0(\design_top.core0.REG1[4][28] ),
    .A1(\design_top.core0.REG1[5][28] ),
    .A2(\design_top.core0.REG1[6][28] ),
    .A3(\design_top.core0.REG1[7][28] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21643_ (.A0(\design_top.core0.REG1[8][28] ),
    .A1(\design_top.core0.REG1[9][28] ),
    .A2(\design_top.core0.REG1[10][28] ),
    .A3(\design_top.core0.REG1[11][28] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21644_ (.A0(\design_top.core0.REG1[12][28] ),
    .A1(\design_top.core0.REG1[13][28] ),
    .A2(\design_top.core0.REG1[14][28] ),
    .A3(\design_top.core0.REG1[15][28] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21645_ (.A0(_02697_),
    .A1(_02698_),
    .A2(_02699_),
    .A3(_02700_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21646_ (.A0(\design_top.core0.REG1[0][29] ),
    .A1(\design_top.core0.REG1[1][29] ),
    .A2(\design_top.core0.REG1[2][29] ),
    .A3(\design_top.core0.REG1[3][29] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21647_ (.A0(\design_top.core0.REG1[4][29] ),
    .A1(\design_top.core0.REG1[5][29] ),
    .A2(\design_top.core0.REG1[6][29] ),
    .A3(\design_top.core0.REG1[7][29] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21648_ (.A0(\design_top.core0.REG1[8][29] ),
    .A1(\design_top.core0.REG1[9][29] ),
    .A2(\design_top.core0.REG1[10][29] ),
    .A3(\design_top.core0.REG1[11][29] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21649_ (.A0(\design_top.core0.REG1[12][29] ),
    .A1(\design_top.core0.REG1[13][29] ),
    .A2(\design_top.core0.REG1[14][29] ),
    .A3(\design_top.core0.REG1[15][29] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21650_ (.A0(_02691_),
    .A1(_02692_),
    .A2(_02693_),
    .A3(_02694_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21651_ (.A0(\design_top.core0.REG1[0][30] ),
    .A1(\design_top.core0.REG1[1][30] ),
    .A2(\design_top.core0.REG1[2][30] ),
    .A3(\design_top.core0.REG1[3][30] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21652_ (.A0(\design_top.core0.REG1[4][30] ),
    .A1(\design_top.core0.REG1[5][30] ),
    .A2(\design_top.core0.REG1[6][30] ),
    .A3(\design_top.core0.REG1[7][30] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21653_ (.A0(\design_top.core0.REG1[8][30] ),
    .A1(\design_top.core0.REG1[9][30] ),
    .A2(\design_top.core0.REG1[10][30] ),
    .A3(\design_top.core0.REG1[11][30] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21654_ (.A0(\design_top.core0.REG1[12][30] ),
    .A1(\design_top.core0.REG1[13][30] ),
    .A2(\design_top.core0.REG1[14][30] ),
    .A3(\design_top.core0.REG1[15][30] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21655_ (.A0(_02685_),
    .A1(_02686_),
    .A2(_02687_),
    .A3(_02688_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21656_ (.A0(_02664_),
    .A1(_02665_),
    .A2(_02666_),
    .A3(_02667_),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21657_ (.A0(_02669_),
    .A1(_02670_),
    .A2(_02671_),
    .A3(_02672_),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21658_ (.A0(_02674_),
    .A1(_02675_),
    .A2(_02676_),
    .A3(_02677_),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21659_ (.A0(_02679_),
    .A1(_02680_),
    .A2(_02681_),
    .A3(_02682_),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21660_ (.A0(_02668_),
    .A1(_02673_),
    .A2(_02678_),
    .A3(_02683_),
    .S0(_00687_),
    .S1(_00688_),
    .X(_02684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21661_ (.A0(\design_top.core0.REG1[8][3] ),
    .A1(\design_top.core0.REG1[9][3] ),
    .A2(\design_top.core0.REG1[10][3] ),
    .A3(\design_top.core0.REG1[11][3] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21662_ (.A0(\design_top.core0.REG1[12][3] ),
    .A1(\design_top.core0.REG1[13][3] ),
    .A2(\design_top.core0.REG1[14][3] ),
    .A3(\design_top.core0.REG1[15][3] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21663_ (.A0(\design_top.core0.REG1[0][3] ),
    .A1(\design_top.core0.REG1[1][3] ),
    .A2(\design_top.core0.REG1[2][3] ),
    .A3(\design_top.core0.REG1[3][3] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21664_ (.A0(\design_top.core0.REG1[4][3] ),
    .A1(\design_top.core0.REG1[5][3] ),
    .A2(\design_top.core0.REG1[6][3] ),
    .A3(\design_top.core0.REG1[7][3] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21665_ (.A0(\design_top.core0.REG1[8][0] ),
    .A1(\design_top.core0.REG1[9][0] ),
    .A2(\design_top.core0.REG1[10][0] ),
    .A3(\design_top.core0.REG1[11][0] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21666_ (.A0(\design_top.core0.REG1[12][0] ),
    .A1(\design_top.core0.REG1[13][0] ),
    .A2(\design_top.core0.REG1[14][0] ),
    .A3(\design_top.core0.REG1[15][0] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21667_ (.A0(\design_top.core0.REG1[0][0] ),
    .A1(\design_top.core0.REG1[1][0] ),
    .A2(\design_top.core0.REG1[2][0] ),
    .A3(\design_top.core0.REG1[3][0] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21668_ (.A0(\design_top.core0.REG1[4][0] ),
    .A1(\design_top.core0.REG1[5][0] ),
    .A2(\design_top.core0.REG1[6][0] ),
    .A3(\design_top.core0.REG1[7][0] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21669_ (.A0(\design_top.core0.REG1[8][1] ),
    .A1(\design_top.core0.REG1[9][1] ),
    .A2(\design_top.core0.REG1[10][1] ),
    .A3(\design_top.core0.REG1[11][1] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21670_ (.A0(\design_top.core0.REG1[12][1] ),
    .A1(\design_top.core0.REG1[13][1] ),
    .A2(\design_top.core0.REG1[14][1] ),
    .A3(\design_top.core0.REG1[15][1] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21671_ (.A0(\design_top.core0.REG1[0][1] ),
    .A1(\design_top.core0.REG1[1][1] ),
    .A2(\design_top.core0.REG1[2][1] ),
    .A3(\design_top.core0.REG1[3][1] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21672_ (.A0(\design_top.core0.REG1[4][1] ),
    .A1(\design_top.core0.REG1[5][1] ),
    .A2(\design_top.core0.REG1[6][1] ),
    .A3(\design_top.core0.REG1[7][1] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21673_ (.A0(\design_top.core0.REG1[8][2] ),
    .A1(\design_top.core0.REG1[9][2] ),
    .A2(\design_top.core0.REG1[10][2] ),
    .A3(\design_top.core0.REG1[11][2] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21674_ (.A0(\design_top.core0.REG1[12][2] ),
    .A1(\design_top.core0.REG1[13][2] ),
    .A2(\design_top.core0.REG1[14][2] ),
    .A3(\design_top.core0.REG1[15][2] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21675_ (.A0(\design_top.core0.REG1[0][2] ),
    .A1(\design_top.core0.REG1[1][2] ),
    .A2(\design_top.core0.REG1[2][2] ),
    .A3(\design_top.core0.REG1[3][2] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21676_ (.A0(\design_top.core0.REG1[4][2] ),
    .A1(\design_top.core0.REG1[5][2] ),
    .A2(\design_top.core0.REG1[6][2] ),
    .A3(\design_top.core0.REG1[7][2] ),
    .S0(_00685_),
    .S1(_00686_),
    .X(_02629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21677_ (.A0(\design_top.MEM[63][31] ),
    .A1(\design_top.MEM[62][31] ),
    .A2(\design_top.MEM[61][31] ),
    .A3(\design_top.MEM[60][31] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21678_ (.A0(\design_top.MEM[59][31] ),
    .A1(\design_top.MEM[58][31] ),
    .A2(\design_top.MEM[57][31] ),
    .A3(\design_top.MEM[56][31] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21679_ (.A0(\design_top.MEM[55][31] ),
    .A1(\design_top.MEM[54][31] ),
    .A2(\design_top.MEM[53][31] ),
    .A3(\design_top.MEM[52][31] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21680_ (.A0(\design_top.MEM[51][31] ),
    .A1(\design_top.MEM[50][31] ),
    .A2(\design_top.MEM[49][31] ),
    .A3(\design_top.MEM[48][31] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21681_ (.A0(_02621_),
    .A1(_02620_),
    .A2(_02619_),
    .A3(_02618_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21682_ (.A0(\design_top.MEM[47][31] ),
    .A1(\design_top.MEM[46][31] ),
    .A2(\design_top.MEM[45][31] ),
    .A3(\design_top.MEM[44][31] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21683_ (.A0(\design_top.MEM[43][31] ),
    .A1(\design_top.MEM[42][31] ),
    .A2(\design_top.MEM[41][31] ),
    .A3(\design_top.MEM[40][31] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21684_ (.A0(\design_top.MEM[39][31] ),
    .A1(\design_top.MEM[38][31] ),
    .A2(\design_top.MEM[37][31] ),
    .A3(\design_top.MEM[36][31] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21685_ (.A0(\design_top.MEM[35][31] ),
    .A1(\design_top.MEM[34][31] ),
    .A2(\design_top.MEM[33][31] ),
    .A3(\design_top.MEM[32][31] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21686_ (.A0(_02616_),
    .A1(_02615_),
    .A2(_02614_),
    .A3(_02613_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21687_ (.A0(\design_top.MEM[31][31] ),
    .A1(\design_top.MEM[30][31] ),
    .A2(\design_top.MEM[29][31] ),
    .A3(\design_top.MEM[28][31] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21688_ (.A0(\design_top.MEM[27][31] ),
    .A1(\design_top.MEM[26][31] ),
    .A2(\design_top.MEM[25][31] ),
    .A3(\design_top.MEM[24][31] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21689_ (.A0(\design_top.MEM[23][31] ),
    .A1(\design_top.MEM[22][31] ),
    .A2(\design_top.MEM[21][31] ),
    .A3(\design_top.MEM[20][31] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21690_ (.A0(\design_top.MEM[19][31] ),
    .A1(\design_top.MEM[18][31] ),
    .A2(\design_top.MEM[17][31] ),
    .A3(\design_top.MEM[16][31] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21691_ (.A0(_02611_),
    .A1(_02610_),
    .A2(_02609_),
    .A3(_02608_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21692_ (.A0(\design_top.MEM[15][31] ),
    .A1(\design_top.MEM[14][31] ),
    .A2(\design_top.MEM[13][31] ),
    .A3(\design_top.MEM[12][31] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21693_ (.A0(\design_top.MEM[11][31] ),
    .A1(\design_top.MEM[10][31] ),
    .A2(\design_top.MEM[9][31] ),
    .A3(\design_top.MEM[8][31] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21694_ (.A0(\design_top.MEM[7][31] ),
    .A1(\design_top.MEM[6][31] ),
    .A2(\design_top.MEM[5][31] ),
    .A3(\design_top.MEM[4][31] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21695_ (.A0(\design_top.MEM[3][31] ),
    .A1(\design_top.MEM[2][31] ),
    .A2(\design_top.MEM[1][31] ),
    .A3(\design_top.MEM[0][31] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21696_ (.A0(_02606_),
    .A1(_02605_),
    .A2(_02604_),
    .A3(_02603_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21697_ (.A0(_02622_),
    .A1(_02617_),
    .A2(_02612_),
    .A3(_02607_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21698_ (.A0(\design_top.MEM[63][30] ),
    .A1(\design_top.MEM[62][30] ),
    .A2(\design_top.MEM[61][30] ),
    .A3(\design_top.MEM[60][30] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21699_ (.A0(\design_top.MEM[59][30] ),
    .A1(\design_top.MEM[58][30] ),
    .A2(\design_top.MEM[57][30] ),
    .A3(\design_top.MEM[56][30] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21700_ (.A0(\design_top.MEM[55][30] ),
    .A1(\design_top.MEM[54][30] ),
    .A2(\design_top.MEM[53][30] ),
    .A3(\design_top.MEM[52][30] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21701_ (.A0(\design_top.MEM[51][30] ),
    .A1(\design_top.MEM[50][30] ),
    .A2(\design_top.MEM[49][30] ),
    .A3(\design_top.MEM[48][30] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21702_ (.A0(_02601_),
    .A1(_02600_),
    .A2(_02599_),
    .A3(_02598_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21703_ (.A0(\design_top.MEM[47][30] ),
    .A1(\design_top.MEM[46][30] ),
    .A2(\design_top.MEM[45][30] ),
    .A3(\design_top.MEM[44][30] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21704_ (.A0(\design_top.MEM[43][30] ),
    .A1(\design_top.MEM[42][30] ),
    .A2(\design_top.MEM[41][30] ),
    .A3(\design_top.MEM[40][30] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21705_ (.A0(\design_top.MEM[39][30] ),
    .A1(\design_top.MEM[38][30] ),
    .A2(\design_top.MEM[37][30] ),
    .A3(\design_top.MEM[36][30] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21706_ (.A0(\design_top.MEM[35][30] ),
    .A1(\design_top.MEM[34][30] ),
    .A2(\design_top.MEM[33][30] ),
    .A3(\design_top.MEM[32][30] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21707_ (.A0(_02596_),
    .A1(_02595_),
    .A2(_02594_),
    .A3(_02593_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21708_ (.A0(\design_top.MEM[31][30] ),
    .A1(\design_top.MEM[30][30] ),
    .A2(\design_top.MEM[29][30] ),
    .A3(\design_top.MEM[28][30] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21709_ (.A0(\design_top.MEM[27][30] ),
    .A1(\design_top.MEM[26][30] ),
    .A2(\design_top.MEM[25][30] ),
    .A3(\design_top.MEM[24][30] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21710_ (.A0(\design_top.MEM[23][30] ),
    .A1(\design_top.MEM[22][30] ),
    .A2(\design_top.MEM[21][30] ),
    .A3(\design_top.MEM[20][30] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21711_ (.A0(\design_top.MEM[19][30] ),
    .A1(\design_top.MEM[18][30] ),
    .A2(\design_top.MEM[17][30] ),
    .A3(\design_top.MEM[16][30] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21712_ (.A0(_02591_),
    .A1(_02590_),
    .A2(_02589_),
    .A3(_02588_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21713_ (.A0(\design_top.MEM[15][30] ),
    .A1(\design_top.MEM[14][30] ),
    .A2(\design_top.MEM[13][30] ),
    .A3(\design_top.MEM[12][30] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21714_ (.A0(\design_top.MEM[11][30] ),
    .A1(\design_top.MEM[10][30] ),
    .A2(\design_top.MEM[9][30] ),
    .A3(\design_top.MEM[8][30] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21715_ (.A0(\design_top.MEM[7][30] ),
    .A1(\design_top.MEM[6][30] ),
    .A2(\design_top.MEM[5][30] ),
    .A3(\design_top.MEM[4][30] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21716_ (.A0(\design_top.MEM[3][30] ),
    .A1(\design_top.MEM[2][30] ),
    .A2(\design_top.MEM[1][30] ),
    .A3(\design_top.MEM[0][30] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21717_ (.A0(_02586_),
    .A1(_02585_),
    .A2(_02584_),
    .A3(_02583_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21718_ (.A0(_02602_),
    .A1(_02597_),
    .A2(_02592_),
    .A3(_02587_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21719_ (.A0(\design_top.MEM[63][29] ),
    .A1(\design_top.MEM[62][29] ),
    .A2(\design_top.MEM[61][29] ),
    .A3(\design_top.MEM[60][29] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21720_ (.A0(\design_top.MEM[59][29] ),
    .A1(\design_top.MEM[58][29] ),
    .A2(\design_top.MEM[57][29] ),
    .A3(\design_top.MEM[56][29] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21721_ (.A0(\design_top.MEM[55][29] ),
    .A1(\design_top.MEM[54][29] ),
    .A2(\design_top.MEM[53][29] ),
    .A3(\design_top.MEM[52][29] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21722_ (.A0(\design_top.MEM[51][29] ),
    .A1(\design_top.MEM[50][29] ),
    .A2(\design_top.MEM[49][29] ),
    .A3(\design_top.MEM[48][29] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21723_ (.A0(_02581_),
    .A1(_02580_),
    .A2(_02579_),
    .A3(_02578_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21724_ (.A0(\design_top.MEM[47][29] ),
    .A1(\design_top.MEM[46][29] ),
    .A2(\design_top.MEM[45][29] ),
    .A3(\design_top.MEM[44][29] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21725_ (.A0(\design_top.MEM[43][29] ),
    .A1(\design_top.MEM[42][29] ),
    .A2(\design_top.MEM[41][29] ),
    .A3(\design_top.MEM[40][29] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21726_ (.A0(\design_top.MEM[39][29] ),
    .A1(\design_top.MEM[38][29] ),
    .A2(\design_top.MEM[37][29] ),
    .A3(\design_top.MEM[36][29] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21727_ (.A0(\design_top.MEM[35][29] ),
    .A1(\design_top.MEM[34][29] ),
    .A2(\design_top.MEM[33][29] ),
    .A3(\design_top.MEM[32][29] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21728_ (.A0(_02576_),
    .A1(_02575_),
    .A2(_02574_),
    .A3(_02573_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21729_ (.A0(\design_top.MEM[31][29] ),
    .A1(\design_top.MEM[30][29] ),
    .A2(\design_top.MEM[29][29] ),
    .A3(\design_top.MEM[28][29] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21730_ (.A0(\design_top.MEM[27][29] ),
    .A1(\design_top.MEM[26][29] ),
    .A2(\design_top.MEM[25][29] ),
    .A3(\design_top.MEM[24][29] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21731_ (.A0(\design_top.MEM[23][29] ),
    .A1(\design_top.MEM[22][29] ),
    .A2(\design_top.MEM[21][29] ),
    .A3(\design_top.MEM[20][29] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21732_ (.A0(\design_top.MEM[19][29] ),
    .A1(\design_top.MEM[18][29] ),
    .A2(\design_top.MEM[17][29] ),
    .A3(\design_top.MEM[16][29] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21733_ (.A0(_02571_),
    .A1(_02570_),
    .A2(_02569_),
    .A3(_02568_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21734_ (.A0(\design_top.MEM[15][29] ),
    .A1(\design_top.MEM[14][29] ),
    .A2(\design_top.MEM[13][29] ),
    .A3(\design_top.MEM[12][29] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21735_ (.A0(\design_top.MEM[11][29] ),
    .A1(\design_top.MEM[10][29] ),
    .A2(\design_top.MEM[9][29] ),
    .A3(\design_top.MEM[8][29] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21736_ (.A0(\design_top.MEM[7][29] ),
    .A1(\design_top.MEM[6][29] ),
    .A2(\design_top.MEM[5][29] ),
    .A3(\design_top.MEM[4][29] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21737_ (.A0(\design_top.MEM[3][29] ),
    .A1(\design_top.MEM[2][29] ),
    .A2(\design_top.MEM[1][29] ),
    .A3(\design_top.MEM[0][29] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21738_ (.A0(_02566_),
    .A1(_02565_),
    .A2(_02564_),
    .A3(_02563_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21739_ (.A0(_02582_),
    .A1(_02577_),
    .A2(_02572_),
    .A3(_02567_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21740_ (.A0(\design_top.MEM[63][28] ),
    .A1(\design_top.MEM[62][28] ),
    .A2(\design_top.MEM[61][28] ),
    .A3(\design_top.MEM[60][28] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21741_ (.A0(\design_top.MEM[59][28] ),
    .A1(\design_top.MEM[58][28] ),
    .A2(\design_top.MEM[57][28] ),
    .A3(\design_top.MEM[56][28] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21742_ (.A0(\design_top.MEM[55][28] ),
    .A1(\design_top.MEM[54][28] ),
    .A2(\design_top.MEM[53][28] ),
    .A3(\design_top.MEM[52][28] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21743_ (.A0(\design_top.MEM[51][28] ),
    .A1(\design_top.MEM[50][28] ),
    .A2(\design_top.MEM[49][28] ),
    .A3(\design_top.MEM[48][28] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21744_ (.A0(_02561_),
    .A1(_02560_),
    .A2(_02559_),
    .A3(_02558_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21745_ (.A0(\design_top.MEM[47][28] ),
    .A1(\design_top.MEM[46][28] ),
    .A2(\design_top.MEM[45][28] ),
    .A3(\design_top.MEM[44][28] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21746_ (.A0(\design_top.MEM[43][28] ),
    .A1(\design_top.MEM[42][28] ),
    .A2(\design_top.MEM[41][28] ),
    .A3(\design_top.MEM[40][28] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21747_ (.A0(\design_top.MEM[39][28] ),
    .A1(\design_top.MEM[38][28] ),
    .A2(\design_top.MEM[37][28] ),
    .A3(\design_top.MEM[36][28] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21748_ (.A0(\design_top.MEM[35][28] ),
    .A1(\design_top.MEM[34][28] ),
    .A2(\design_top.MEM[33][28] ),
    .A3(\design_top.MEM[32][28] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21749_ (.A0(_02556_),
    .A1(_02555_),
    .A2(_02554_),
    .A3(_02553_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21750_ (.A0(\design_top.MEM[31][28] ),
    .A1(\design_top.MEM[30][28] ),
    .A2(\design_top.MEM[29][28] ),
    .A3(\design_top.MEM[28][28] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21751_ (.A0(\design_top.MEM[27][28] ),
    .A1(\design_top.MEM[26][28] ),
    .A2(\design_top.MEM[25][28] ),
    .A3(\design_top.MEM[24][28] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21752_ (.A0(\design_top.MEM[23][28] ),
    .A1(\design_top.MEM[22][28] ),
    .A2(\design_top.MEM[21][28] ),
    .A3(\design_top.MEM[20][28] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21753_ (.A0(\design_top.MEM[19][28] ),
    .A1(\design_top.MEM[18][28] ),
    .A2(\design_top.MEM[17][28] ),
    .A3(\design_top.MEM[16][28] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21754_ (.A0(_02551_),
    .A1(_02550_),
    .A2(_02549_),
    .A3(_02548_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21755_ (.A0(\design_top.MEM[15][28] ),
    .A1(\design_top.MEM[14][28] ),
    .A2(\design_top.MEM[13][28] ),
    .A3(\design_top.MEM[12][28] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21756_ (.A0(\design_top.MEM[11][28] ),
    .A1(\design_top.MEM[10][28] ),
    .A2(\design_top.MEM[9][28] ),
    .A3(\design_top.MEM[8][28] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21757_ (.A0(\design_top.MEM[7][28] ),
    .A1(\design_top.MEM[6][28] ),
    .A2(\design_top.MEM[5][28] ),
    .A3(\design_top.MEM[4][28] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21758_ (.A0(\design_top.MEM[3][28] ),
    .A1(\design_top.MEM[2][28] ),
    .A2(\design_top.MEM[1][28] ),
    .A3(\design_top.MEM[0][28] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21759_ (.A0(_02546_),
    .A1(_02545_),
    .A2(_02544_),
    .A3(_02543_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21760_ (.A0(_02562_),
    .A1(_02557_),
    .A2(_02552_),
    .A3(_02547_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21761_ (.A0(\design_top.MEM[63][27] ),
    .A1(\design_top.MEM[62][27] ),
    .A2(\design_top.MEM[61][27] ),
    .A3(\design_top.MEM[60][27] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21762_ (.A0(\design_top.MEM[59][27] ),
    .A1(\design_top.MEM[58][27] ),
    .A2(\design_top.MEM[57][27] ),
    .A3(\design_top.MEM[56][27] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21763_ (.A0(\design_top.MEM[55][27] ),
    .A1(\design_top.MEM[54][27] ),
    .A2(\design_top.MEM[53][27] ),
    .A3(\design_top.MEM[52][27] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21764_ (.A0(\design_top.MEM[51][27] ),
    .A1(\design_top.MEM[50][27] ),
    .A2(\design_top.MEM[49][27] ),
    .A3(\design_top.MEM[48][27] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21765_ (.A0(_02541_),
    .A1(_02540_),
    .A2(_02539_),
    .A3(_02538_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21766_ (.A0(\design_top.MEM[47][27] ),
    .A1(\design_top.MEM[46][27] ),
    .A2(\design_top.MEM[45][27] ),
    .A3(\design_top.MEM[44][27] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21767_ (.A0(\design_top.MEM[43][27] ),
    .A1(\design_top.MEM[42][27] ),
    .A2(\design_top.MEM[41][27] ),
    .A3(\design_top.MEM[40][27] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21768_ (.A0(\design_top.MEM[39][27] ),
    .A1(\design_top.MEM[38][27] ),
    .A2(\design_top.MEM[37][27] ),
    .A3(\design_top.MEM[36][27] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21769_ (.A0(\design_top.MEM[35][27] ),
    .A1(\design_top.MEM[34][27] ),
    .A2(\design_top.MEM[33][27] ),
    .A3(\design_top.MEM[32][27] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21770_ (.A0(_02536_),
    .A1(_02535_),
    .A2(_02534_),
    .A3(_02533_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21771_ (.A0(\design_top.MEM[31][27] ),
    .A1(\design_top.MEM[30][27] ),
    .A2(\design_top.MEM[29][27] ),
    .A3(\design_top.MEM[28][27] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21772_ (.A0(\design_top.MEM[27][27] ),
    .A1(\design_top.MEM[26][27] ),
    .A2(\design_top.MEM[25][27] ),
    .A3(\design_top.MEM[24][27] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21773_ (.A0(\design_top.MEM[23][27] ),
    .A1(\design_top.MEM[22][27] ),
    .A2(\design_top.MEM[21][27] ),
    .A3(\design_top.MEM[20][27] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21774_ (.A0(\design_top.MEM[19][27] ),
    .A1(\design_top.MEM[18][27] ),
    .A2(\design_top.MEM[17][27] ),
    .A3(\design_top.MEM[16][27] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21775_ (.A0(_02531_),
    .A1(_02530_),
    .A2(_02529_),
    .A3(_02528_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21776_ (.A0(\design_top.MEM[15][27] ),
    .A1(\design_top.MEM[14][27] ),
    .A2(\design_top.MEM[13][27] ),
    .A3(\design_top.MEM[12][27] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21777_ (.A0(\design_top.MEM[11][27] ),
    .A1(\design_top.MEM[10][27] ),
    .A2(\design_top.MEM[9][27] ),
    .A3(\design_top.MEM[8][27] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21778_ (.A0(\design_top.MEM[7][27] ),
    .A1(\design_top.MEM[6][27] ),
    .A2(\design_top.MEM[5][27] ),
    .A3(\design_top.MEM[4][27] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21779_ (.A0(\design_top.MEM[3][27] ),
    .A1(\design_top.MEM[2][27] ),
    .A2(\design_top.MEM[1][27] ),
    .A3(\design_top.MEM[0][27] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21780_ (.A0(_02526_),
    .A1(_02525_),
    .A2(_02524_),
    .A3(_02523_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21781_ (.A0(_02542_),
    .A1(_02537_),
    .A2(_02532_),
    .A3(_02527_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21782_ (.A0(\design_top.MEM[63][26] ),
    .A1(\design_top.MEM[62][26] ),
    .A2(\design_top.MEM[61][26] ),
    .A3(\design_top.MEM[60][26] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21783_ (.A0(\design_top.MEM[59][26] ),
    .A1(\design_top.MEM[58][26] ),
    .A2(\design_top.MEM[57][26] ),
    .A3(\design_top.MEM[56][26] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21784_ (.A0(\design_top.MEM[55][26] ),
    .A1(\design_top.MEM[54][26] ),
    .A2(\design_top.MEM[53][26] ),
    .A3(\design_top.MEM[52][26] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21785_ (.A0(\design_top.MEM[51][26] ),
    .A1(\design_top.MEM[50][26] ),
    .A2(\design_top.MEM[49][26] ),
    .A3(\design_top.MEM[48][26] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21786_ (.A0(_02521_),
    .A1(_02520_),
    .A2(_02519_),
    .A3(_02518_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21787_ (.A0(\design_top.MEM[47][26] ),
    .A1(\design_top.MEM[46][26] ),
    .A2(\design_top.MEM[45][26] ),
    .A3(\design_top.MEM[44][26] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21788_ (.A0(\design_top.MEM[43][26] ),
    .A1(\design_top.MEM[42][26] ),
    .A2(\design_top.MEM[41][26] ),
    .A3(\design_top.MEM[40][26] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21789_ (.A0(\design_top.MEM[39][26] ),
    .A1(\design_top.MEM[38][26] ),
    .A2(\design_top.MEM[37][26] ),
    .A3(\design_top.MEM[36][26] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21790_ (.A0(\design_top.MEM[35][26] ),
    .A1(\design_top.MEM[34][26] ),
    .A2(\design_top.MEM[33][26] ),
    .A3(\design_top.MEM[32][26] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21791_ (.A0(_02516_),
    .A1(_02515_),
    .A2(_02514_),
    .A3(_02513_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21792_ (.A0(\design_top.MEM[31][26] ),
    .A1(\design_top.MEM[30][26] ),
    .A2(\design_top.MEM[29][26] ),
    .A3(\design_top.MEM[28][26] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21793_ (.A0(\design_top.MEM[27][26] ),
    .A1(\design_top.MEM[26][26] ),
    .A2(\design_top.MEM[25][26] ),
    .A3(\design_top.MEM[24][26] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21794_ (.A0(\design_top.MEM[23][26] ),
    .A1(\design_top.MEM[22][26] ),
    .A2(\design_top.MEM[21][26] ),
    .A3(\design_top.MEM[20][26] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21795_ (.A0(\design_top.MEM[19][26] ),
    .A1(\design_top.MEM[18][26] ),
    .A2(\design_top.MEM[17][26] ),
    .A3(\design_top.MEM[16][26] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21796_ (.A0(_02511_),
    .A1(_02510_),
    .A2(_02509_),
    .A3(_02508_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21797_ (.A0(\design_top.MEM[15][26] ),
    .A1(\design_top.MEM[14][26] ),
    .A2(\design_top.MEM[13][26] ),
    .A3(\design_top.MEM[12][26] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21798_ (.A0(\design_top.MEM[11][26] ),
    .A1(\design_top.MEM[10][26] ),
    .A2(\design_top.MEM[9][26] ),
    .A3(\design_top.MEM[8][26] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21799_ (.A0(\design_top.MEM[7][26] ),
    .A1(\design_top.MEM[6][26] ),
    .A2(\design_top.MEM[5][26] ),
    .A3(\design_top.MEM[4][26] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21800_ (.A0(\design_top.MEM[3][26] ),
    .A1(\design_top.MEM[2][26] ),
    .A2(\design_top.MEM[1][26] ),
    .A3(\design_top.MEM[0][26] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21801_ (.A0(_02506_),
    .A1(_02505_),
    .A2(_02504_),
    .A3(_02503_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21802_ (.A0(_02522_),
    .A1(_02517_),
    .A2(_02512_),
    .A3(_02507_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21803_ (.A0(\design_top.MEM[63][25] ),
    .A1(\design_top.MEM[62][25] ),
    .A2(\design_top.MEM[61][25] ),
    .A3(\design_top.MEM[60][25] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21804_ (.A0(\design_top.MEM[59][25] ),
    .A1(\design_top.MEM[58][25] ),
    .A2(\design_top.MEM[57][25] ),
    .A3(\design_top.MEM[56][25] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21805_ (.A0(\design_top.MEM[55][25] ),
    .A1(\design_top.MEM[54][25] ),
    .A2(\design_top.MEM[53][25] ),
    .A3(\design_top.MEM[52][25] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21806_ (.A0(\design_top.MEM[51][25] ),
    .A1(\design_top.MEM[50][25] ),
    .A2(\design_top.MEM[49][25] ),
    .A3(\design_top.MEM[48][25] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21807_ (.A0(_02501_),
    .A1(_02500_),
    .A2(_02499_),
    .A3(_02498_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21808_ (.A0(\design_top.MEM[47][25] ),
    .A1(\design_top.MEM[46][25] ),
    .A2(\design_top.MEM[45][25] ),
    .A3(\design_top.MEM[44][25] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21809_ (.A0(\design_top.MEM[43][25] ),
    .A1(\design_top.MEM[42][25] ),
    .A2(\design_top.MEM[41][25] ),
    .A3(\design_top.MEM[40][25] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21810_ (.A0(\design_top.MEM[39][25] ),
    .A1(\design_top.MEM[38][25] ),
    .A2(\design_top.MEM[37][25] ),
    .A3(\design_top.MEM[36][25] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21811_ (.A0(\design_top.MEM[35][25] ),
    .A1(\design_top.MEM[34][25] ),
    .A2(\design_top.MEM[33][25] ),
    .A3(\design_top.MEM[32][25] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21812_ (.A0(_02496_),
    .A1(_02495_),
    .A2(_02494_),
    .A3(_02493_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21813_ (.A0(\design_top.MEM[31][25] ),
    .A1(\design_top.MEM[30][25] ),
    .A2(\design_top.MEM[29][25] ),
    .A3(\design_top.MEM[28][25] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21814_ (.A0(\design_top.MEM[27][25] ),
    .A1(\design_top.MEM[26][25] ),
    .A2(\design_top.MEM[25][25] ),
    .A3(\design_top.MEM[24][25] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21815_ (.A0(\design_top.MEM[23][25] ),
    .A1(\design_top.MEM[22][25] ),
    .A2(\design_top.MEM[21][25] ),
    .A3(\design_top.MEM[20][25] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21816_ (.A0(\design_top.MEM[19][25] ),
    .A1(\design_top.MEM[18][25] ),
    .A2(\design_top.MEM[17][25] ),
    .A3(\design_top.MEM[16][25] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21817_ (.A0(_02491_),
    .A1(_02490_),
    .A2(_02489_),
    .A3(_02488_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21818_ (.A0(\design_top.MEM[15][25] ),
    .A1(\design_top.MEM[14][25] ),
    .A2(\design_top.MEM[13][25] ),
    .A3(\design_top.MEM[12][25] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21819_ (.A0(\design_top.MEM[11][25] ),
    .A1(\design_top.MEM[10][25] ),
    .A2(\design_top.MEM[9][25] ),
    .A3(\design_top.MEM[8][25] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21820_ (.A0(\design_top.MEM[7][25] ),
    .A1(\design_top.MEM[6][25] ),
    .A2(\design_top.MEM[5][25] ),
    .A3(\design_top.MEM[4][25] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21821_ (.A0(\design_top.MEM[3][25] ),
    .A1(\design_top.MEM[2][25] ),
    .A2(\design_top.MEM[1][25] ),
    .A3(\design_top.MEM[0][25] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21822_ (.A0(_02486_),
    .A1(_02485_),
    .A2(_02484_),
    .A3(_02483_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21823_ (.A0(_02502_),
    .A1(_02497_),
    .A2(_02492_),
    .A3(_02487_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21824_ (.A0(\design_top.MEM[63][24] ),
    .A1(\design_top.MEM[62][24] ),
    .A2(\design_top.MEM[61][24] ),
    .A3(\design_top.MEM[60][24] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21825_ (.A0(\design_top.MEM[59][24] ),
    .A1(\design_top.MEM[58][24] ),
    .A2(\design_top.MEM[57][24] ),
    .A3(\design_top.MEM[56][24] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21826_ (.A0(\design_top.MEM[55][24] ),
    .A1(\design_top.MEM[54][24] ),
    .A2(\design_top.MEM[53][24] ),
    .A3(\design_top.MEM[52][24] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21827_ (.A0(\design_top.MEM[51][24] ),
    .A1(\design_top.MEM[50][24] ),
    .A2(\design_top.MEM[49][24] ),
    .A3(\design_top.MEM[48][24] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21828_ (.A0(_02481_),
    .A1(_02480_),
    .A2(_02479_),
    .A3(_02478_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21829_ (.A0(\design_top.MEM[47][24] ),
    .A1(\design_top.MEM[46][24] ),
    .A2(\design_top.MEM[45][24] ),
    .A3(\design_top.MEM[44][24] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21830_ (.A0(\design_top.MEM[43][24] ),
    .A1(\design_top.MEM[42][24] ),
    .A2(\design_top.MEM[41][24] ),
    .A3(\design_top.MEM[40][24] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21831_ (.A0(\design_top.MEM[39][24] ),
    .A1(\design_top.MEM[38][24] ),
    .A2(\design_top.MEM[37][24] ),
    .A3(\design_top.MEM[36][24] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21832_ (.A0(\design_top.MEM[35][24] ),
    .A1(\design_top.MEM[34][24] ),
    .A2(\design_top.MEM[33][24] ),
    .A3(\design_top.MEM[32][24] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21833_ (.A0(_02476_),
    .A1(_02475_),
    .A2(_02474_),
    .A3(_02473_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21834_ (.A0(\design_top.MEM[31][24] ),
    .A1(\design_top.MEM[30][24] ),
    .A2(\design_top.MEM[29][24] ),
    .A3(\design_top.MEM[28][24] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21835_ (.A0(\design_top.MEM[27][24] ),
    .A1(\design_top.MEM[26][24] ),
    .A2(\design_top.MEM[25][24] ),
    .A3(\design_top.MEM[24][24] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21836_ (.A0(\design_top.MEM[23][24] ),
    .A1(\design_top.MEM[22][24] ),
    .A2(\design_top.MEM[21][24] ),
    .A3(\design_top.MEM[20][24] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21837_ (.A0(\design_top.MEM[19][24] ),
    .A1(\design_top.MEM[18][24] ),
    .A2(\design_top.MEM[17][24] ),
    .A3(\design_top.MEM[16][24] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21838_ (.A0(_02471_),
    .A1(_02470_),
    .A2(_02469_),
    .A3(_02468_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21839_ (.A0(\design_top.MEM[15][24] ),
    .A1(\design_top.MEM[14][24] ),
    .A2(\design_top.MEM[13][24] ),
    .A3(\design_top.MEM[12][24] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21840_ (.A0(\design_top.MEM[11][24] ),
    .A1(\design_top.MEM[10][24] ),
    .A2(\design_top.MEM[9][24] ),
    .A3(\design_top.MEM[8][24] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21841_ (.A0(\design_top.MEM[7][24] ),
    .A1(\design_top.MEM[6][24] ),
    .A2(\design_top.MEM[5][24] ),
    .A3(\design_top.MEM[4][24] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21842_ (.A0(\design_top.MEM[3][24] ),
    .A1(\design_top.MEM[2][24] ),
    .A2(\design_top.MEM[1][24] ),
    .A3(\design_top.MEM[0][24] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21843_ (.A0(_02466_),
    .A1(_02465_),
    .A2(_02464_),
    .A3(_02463_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21844_ (.A0(_02482_),
    .A1(_02477_),
    .A2(_02472_),
    .A3(_02467_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21845_ (.A0(\design_top.MEM[63][23] ),
    .A1(\design_top.MEM[62][23] ),
    .A2(\design_top.MEM[61][23] ),
    .A3(\design_top.MEM[60][23] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21846_ (.A0(\design_top.MEM[59][23] ),
    .A1(\design_top.MEM[58][23] ),
    .A2(\design_top.MEM[57][23] ),
    .A3(\design_top.MEM[56][23] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21847_ (.A0(\design_top.MEM[55][23] ),
    .A1(\design_top.MEM[54][23] ),
    .A2(\design_top.MEM[53][23] ),
    .A3(\design_top.MEM[52][23] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21848_ (.A0(\design_top.MEM[51][23] ),
    .A1(\design_top.MEM[50][23] ),
    .A2(\design_top.MEM[49][23] ),
    .A3(\design_top.MEM[48][23] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21849_ (.A0(_02461_),
    .A1(_02460_),
    .A2(_02459_),
    .A3(_02458_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21850_ (.A0(\design_top.MEM[47][23] ),
    .A1(\design_top.MEM[46][23] ),
    .A2(\design_top.MEM[45][23] ),
    .A3(\design_top.MEM[44][23] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21851_ (.A0(\design_top.MEM[43][23] ),
    .A1(\design_top.MEM[42][23] ),
    .A2(\design_top.MEM[41][23] ),
    .A3(\design_top.MEM[40][23] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21852_ (.A0(\design_top.MEM[39][23] ),
    .A1(\design_top.MEM[38][23] ),
    .A2(\design_top.MEM[37][23] ),
    .A3(\design_top.MEM[36][23] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21853_ (.A0(\design_top.MEM[35][23] ),
    .A1(\design_top.MEM[34][23] ),
    .A2(\design_top.MEM[33][23] ),
    .A3(\design_top.MEM[32][23] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21854_ (.A0(_02456_),
    .A1(_02455_),
    .A2(_02454_),
    .A3(_02453_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21855_ (.A0(\design_top.MEM[31][23] ),
    .A1(\design_top.MEM[30][23] ),
    .A2(\design_top.MEM[29][23] ),
    .A3(\design_top.MEM[28][23] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21856_ (.A0(\design_top.MEM[27][23] ),
    .A1(\design_top.MEM[26][23] ),
    .A2(\design_top.MEM[25][23] ),
    .A3(\design_top.MEM[24][23] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21857_ (.A0(\design_top.MEM[23][23] ),
    .A1(\design_top.MEM[22][23] ),
    .A2(\design_top.MEM[21][23] ),
    .A3(\design_top.MEM[20][23] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21858_ (.A0(\design_top.MEM[19][23] ),
    .A1(\design_top.MEM[18][23] ),
    .A2(\design_top.MEM[17][23] ),
    .A3(\design_top.MEM[16][23] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21859_ (.A0(_02451_),
    .A1(_02450_),
    .A2(_02449_),
    .A3(_02448_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21860_ (.A0(\design_top.MEM[15][23] ),
    .A1(\design_top.MEM[14][23] ),
    .A2(\design_top.MEM[13][23] ),
    .A3(\design_top.MEM[12][23] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21861_ (.A0(\design_top.MEM[11][23] ),
    .A1(\design_top.MEM[10][23] ),
    .A2(\design_top.MEM[9][23] ),
    .A3(\design_top.MEM[8][23] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21862_ (.A0(\design_top.MEM[7][23] ),
    .A1(\design_top.MEM[6][23] ),
    .A2(\design_top.MEM[5][23] ),
    .A3(\design_top.MEM[4][23] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21863_ (.A0(\design_top.MEM[3][23] ),
    .A1(\design_top.MEM[2][23] ),
    .A2(\design_top.MEM[1][23] ),
    .A3(\design_top.MEM[0][23] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21864_ (.A0(_02446_),
    .A1(_02445_),
    .A2(_02444_),
    .A3(_02443_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21865_ (.A0(_02462_),
    .A1(_02457_),
    .A2(_02452_),
    .A3(_02447_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21866_ (.A0(\design_top.MEM[63][22] ),
    .A1(\design_top.MEM[62][22] ),
    .A2(\design_top.MEM[61][22] ),
    .A3(\design_top.MEM[60][22] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21867_ (.A0(\design_top.MEM[59][22] ),
    .A1(\design_top.MEM[58][22] ),
    .A2(\design_top.MEM[57][22] ),
    .A3(\design_top.MEM[56][22] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21868_ (.A0(\design_top.MEM[55][22] ),
    .A1(\design_top.MEM[54][22] ),
    .A2(\design_top.MEM[53][22] ),
    .A3(\design_top.MEM[52][22] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21869_ (.A0(\design_top.MEM[51][22] ),
    .A1(\design_top.MEM[50][22] ),
    .A2(\design_top.MEM[49][22] ),
    .A3(\design_top.MEM[48][22] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21870_ (.A0(_02441_),
    .A1(_02440_),
    .A2(_02439_),
    .A3(_02438_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21871_ (.A0(\design_top.MEM[47][22] ),
    .A1(\design_top.MEM[46][22] ),
    .A2(\design_top.MEM[45][22] ),
    .A3(\design_top.MEM[44][22] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21872_ (.A0(\design_top.MEM[43][22] ),
    .A1(\design_top.MEM[42][22] ),
    .A2(\design_top.MEM[41][22] ),
    .A3(\design_top.MEM[40][22] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21873_ (.A0(\design_top.MEM[39][22] ),
    .A1(\design_top.MEM[38][22] ),
    .A2(\design_top.MEM[37][22] ),
    .A3(\design_top.MEM[36][22] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21874_ (.A0(\design_top.MEM[35][22] ),
    .A1(\design_top.MEM[34][22] ),
    .A2(\design_top.MEM[33][22] ),
    .A3(\design_top.MEM[32][22] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21875_ (.A0(_02436_),
    .A1(_02435_),
    .A2(_02434_),
    .A3(_02433_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21876_ (.A0(\design_top.MEM[31][22] ),
    .A1(\design_top.MEM[30][22] ),
    .A2(\design_top.MEM[29][22] ),
    .A3(\design_top.MEM[28][22] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21877_ (.A0(\design_top.MEM[27][22] ),
    .A1(\design_top.MEM[26][22] ),
    .A2(\design_top.MEM[25][22] ),
    .A3(\design_top.MEM[24][22] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21878_ (.A0(\design_top.MEM[23][22] ),
    .A1(\design_top.MEM[22][22] ),
    .A2(\design_top.MEM[21][22] ),
    .A3(\design_top.MEM[20][22] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21879_ (.A0(\design_top.MEM[19][22] ),
    .A1(\design_top.MEM[18][22] ),
    .A2(\design_top.MEM[17][22] ),
    .A3(\design_top.MEM[16][22] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21880_ (.A0(_02431_),
    .A1(_02430_),
    .A2(_02429_),
    .A3(_02428_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21881_ (.A0(\design_top.MEM[15][22] ),
    .A1(\design_top.MEM[14][22] ),
    .A2(\design_top.MEM[13][22] ),
    .A3(\design_top.MEM[12][22] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21882_ (.A0(\design_top.MEM[11][22] ),
    .A1(\design_top.MEM[10][22] ),
    .A2(\design_top.MEM[9][22] ),
    .A3(\design_top.MEM[8][22] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21883_ (.A0(\design_top.MEM[7][22] ),
    .A1(\design_top.MEM[6][22] ),
    .A2(\design_top.MEM[5][22] ),
    .A3(\design_top.MEM[4][22] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21884_ (.A0(\design_top.MEM[3][22] ),
    .A1(\design_top.MEM[2][22] ),
    .A2(\design_top.MEM[1][22] ),
    .A3(\design_top.MEM[0][22] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21885_ (.A0(_02426_),
    .A1(_02425_),
    .A2(_02424_),
    .A3(_02423_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21886_ (.A0(_02442_),
    .A1(_02437_),
    .A2(_02432_),
    .A3(_02427_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21887_ (.A0(\design_top.MEM[63][21] ),
    .A1(\design_top.MEM[62][21] ),
    .A2(\design_top.MEM[61][21] ),
    .A3(\design_top.MEM[60][21] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21888_ (.A0(\design_top.MEM[59][21] ),
    .A1(\design_top.MEM[58][21] ),
    .A2(\design_top.MEM[57][21] ),
    .A3(\design_top.MEM[56][21] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21889_ (.A0(\design_top.MEM[55][21] ),
    .A1(\design_top.MEM[54][21] ),
    .A2(\design_top.MEM[53][21] ),
    .A3(\design_top.MEM[52][21] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21890_ (.A0(\design_top.MEM[51][21] ),
    .A1(\design_top.MEM[50][21] ),
    .A2(\design_top.MEM[49][21] ),
    .A3(\design_top.MEM[48][21] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21891_ (.A0(_02421_),
    .A1(_02420_),
    .A2(_02419_),
    .A3(_02418_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21892_ (.A0(\design_top.MEM[47][21] ),
    .A1(\design_top.MEM[46][21] ),
    .A2(\design_top.MEM[45][21] ),
    .A3(\design_top.MEM[44][21] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21893_ (.A0(\design_top.MEM[43][21] ),
    .A1(\design_top.MEM[42][21] ),
    .A2(\design_top.MEM[41][21] ),
    .A3(\design_top.MEM[40][21] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21894_ (.A0(\design_top.MEM[39][21] ),
    .A1(\design_top.MEM[38][21] ),
    .A2(\design_top.MEM[37][21] ),
    .A3(\design_top.MEM[36][21] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21895_ (.A0(\design_top.MEM[35][21] ),
    .A1(\design_top.MEM[34][21] ),
    .A2(\design_top.MEM[33][21] ),
    .A3(\design_top.MEM[32][21] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21896_ (.A0(_02416_),
    .A1(_02415_),
    .A2(_02414_),
    .A3(_02413_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21897_ (.A0(\design_top.MEM[31][21] ),
    .A1(\design_top.MEM[30][21] ),
    .A2(\design_top.MEM[29][21] ),
    .A3(\design_top.MEM[28][21] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21898_ (.A0(\design_top.MEM[27][21] ),
    .A1(\design_top.MEM[26][21] ),
    .A2(\design_top.MEM[25][21] ),
    .A3(\design_top.MEM[24][21] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21899_ (.A0(\design_top.MEM[23][21] ),
    .A1(\design_top.MEM[22][21] ),
    .A2(\design_top.MEM[21][21] ),
    .A3(\design_top.MEM[20][21] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21900_ (.A0(\design_top.MEM[19][21] ),
    .A1(\design_top.MEM[18][21] ),
    .A2(\design_top.MEM[17][21] ),
    .A3(\design_top.MEM[16][21] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21901_ (.A0(_02411_),
    .A1(_02410_),
    .A2(_02409_),
    .A3(_02408_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21902_ (.A0(\design_top.MEM[15][21] ),
    .A1(\design_top.MEM[14][21] ),
    .A2(\design_top.MEM[13][21] ),
    .A3(\design_top.MEM[12][21] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21903_ (.A0(\design_top.MEM[11][21] ),
    .A1(\design_top.MEM[10][21] ),
    .A2(\design_top.MEM[9][21] ),
    .A3(\design_top.MEM[8][21] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21904_ (.A0(\design_top.MEM[7][21] ),
    .A1(\design_top.MEM[6][21] ),
    .A2(\design_top.MEM[5][21] ),
    .A3(\design_top.MEM[4][21] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21905_ (.A0(\design_top.MEM[3][21] ),
    .A1(\design_top.MEM[2][21] ),
    .A2(\design_top.MEM[1][21] ),
    .A3(\design_top.MEM[0][21] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21906_ (.A0(_02406_),
    .A1(_02405_),
    .A2(_02404_),
    .A3(_02403_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21907_ (.A0(_02422_),
    .A1(_02417_),
    .A2(_02412_),
    .A3(_02407_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21908_ (.A0(\design_top.MEM[63][20] ),
    .A1(\design_top.MEM[62][20] ),
    .A2(\design_top.MEM[61][20] ),
    .A3(\design_top.MEM[60][20] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21909_ (.A0(\design_top.MEM[59][20] ),
    .A1(\design_top.MEM[58][20] ),
    .A2(\design_top.MEM[57][20] ),
    .A3(\design_top.MEM[56][20] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21910_ (.A0(\design_top.MEM[55][20] ),
    .A1(\design_top.MEM[54][20] ),
    .A2(\design_top.MEM[53][20] ),
    .A3(\design_top.MEM[52][20] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21911_ (.A0(\design_top.MEM[51][20] ),
    .A1(\design_top.MEM[50][20] ),
    .A2(\design_top.MEM[49][20] ),
    .A3(\design_top.MEM[48][20] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21912_ (.A0(_02401_),
    .A1(_02400_),
    .A2(_02399_),
    .A3(_02398_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21913_ (.A0(\design_top.MEM[47][20] ),
    .A1(\design_top.MEM[46][20] ),
    .A2(\design_top.MEM[45][20] ),
    .A3(\design_top.MEM[44][20] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21914_ (.A0(\design_top.MEM[43][20] ),
    .A1(\design_top.MEM[42][20] ),
    .A2(\design_top.MEM[41][20] ),
    .A3(\design_top.MEM[40][20] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21915_ (.A0(\design_top.MEM[39][20] ),
    .A1(\design_top.MEM[38][20] ),
    .A2(\design_top.MEM[37][20] ),
    .A3(\design_top.MEM[36][20] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21916_ (.A0(\design_top.MEM[35][20] ),
    .A1(\design_top.MEM[34][20] ),
    .A2(\design_top.MEM[33][20] ),
    .A3(\design_top.MEM[32][20] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21917_ (.A0(_02396_),
    .A1(_02395_),
    .A2(_02394_),
    .A3(_02393_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21918_ (.A0(\design_top.MEM[31][20] ),
    .A1(\design_top.MEM[30][20] ),
    .A2(\design_top.MEM[29][20] ),
    .A3(\design_top.MEM[28][20] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21919_ (.A0(\design_top.MEM[27][20] ),
    .A1(\design_top.MEM[26][20] ),
    .A2(\design_top.MEM[25][20] ),
    .A3(\design_top.MEM[24][20] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21920_ (.A0(\design_top.MEM[23][20] ),
    .A1(\design_top.MEM[22][20] ),
    .A2(\design_top.MEM[21][20] ),
    .A3(\design_top.MEM[20][20] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21921_ (.A0(\design_top.MEM[19][20] ),
    .A1(\design_top.MEM[18][20] ),
    .A2(\design_top.MEM[17][20] ),
    .A3(\design_top.MEM[16][20] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21922_ (.A0(_02391_),
    .A1(_02390_),
    .A2(_02389_),
    .A3(_02388_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21923_ (.A0(\design_top.MEM[15][20] ),
    .A1(\design_top.MEM[14][20] ),
    .A2(\design_top.MEM[13][20] ),
    .A3(\design_top.MEM[12][20] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21924_ (.A0(\design_top.MEM[11][20] ),
    .A1(\design_top.MEM[10][20] ),
    .A2(\design_top.MEM[9][20] ),
    .A3(\design_top.MEM[8][20] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21925_ (.A0(\design_top.MEM[7][20] ),
    .A1(\design_top.MEM[6][20] ),
    .A2(\design_top.MEM[5][20] ),
    .A3(\design_top.MEM[4][20] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21926_ (.A0(\design_top.MEM[3][20] ),
    .A1(\design_top.MEM[2][20] ),
    .A2(\design_top.MEM[1][20] ),
    .A3(\design_top.MEM[0][20] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21927_ (.A0(_02386_),
    .A1(_02385_),
    .A2(_02384_),
    .A3(_02383_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21928_ (.A0(_02402_),
    .A1(_02397_),
    .A2(_02392_),
    .A3(_02387_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21929_ (.A0(\design_top.MEM[63][19] ),
    .A1(\design_top.MEM[62][19] ),
    .A2(\design_top.MEM[61][19] ),
    .A3(\design_top.MEM[60][19] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21930_ (.A0(\design_top.MEM[59][19] ),
    .A1(\design_top.MEM[58][19] ),
    .A2(\design_top.MEM[57][19] ),
    .A3(\design_top.MEM[56][19] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21931_ (.A0(\design_top.MEM[55][19] ),
    .A1(\design_top.MEM[54][19] ),
    .A2(\design_top.MEM[53][19] ),
    .A3(\design_top.MEM[52][19] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21932_ (.A0(\design_top.MEM[51][19] ),
    .A1(\design_top.MEM[50][19] ),
    .A2(\design_top.MEM[49][19] ),
    .A3(\design_top.MEM[48][19] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21933_ (.A0(_02381_),
    .A1(_02380_),
    .A2(_02379_),
    .A3(_02378_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21934_ (.A0(\design_top.MEM[47][19] ),
    .A1(\design_top.MEM[46][19] ),
    .A2(\design_top.MEM[45][19] ),
    .A3(\design_top.MEM[44][19] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21935_ (.A0(\design_top.MEM[43][19] ),
    .A1(\design_top.MEM[42][19] ),
    .A2(\design_top.MEM[41][19] ),
    .A3(\design_top.MEM[40][19] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21936_ (.A0(\design_top.MEM[39][19] ),
    .A1(\design_top.MEM[38][19] ),
    .A2(\design_top.MEM[37][19] ),
    .A3(\design_top.MEM[36][19] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21937_ (.A0(\design_top.MEM[35][19] ),
    .A1(\design_top.MEM[34][19] ),
    .A2(\design_top.MEM[33][19] ),
    .A3(\design_top.MEM[32][19] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21938_ (.A0(_02376_),
    .A1(_02375_),
    .A2(_02374_),
    .A3(_02373_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21939_ (.A0(\design_top.MEM[31][19] ),
    .A1(\design_top.MEM[30][19] ),
    .A2(\design_top.MEM[29][19] ),
    .A3(\design_top.MEM[28][19] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21940_ (.A0(\design_top.MEM[27][19] ),
    .A1(\design_top.MEM[26][19] ),
    .A2(\design_top.MEM[25][19] ),
    .A3(\design_top.MEM[24][19] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21941_ (.A0(\design_top.MEM[23][19] ),
    .A1(\design_top.MEM[22][19] ),
    .A2(\design_top.MEM[21][19] ),
    .A3(\design_top.MEM[20][19] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21942_ (.A0(\design_top.MEM[19][19] ),
    .A1(\design_top.MEM[18][19] ),
    .A2(\design_top.MEM[17][19] ),
    .A3(\design_top.MEM[16][19] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21943_ (.A0(_02371_),
    .A1(_02370_),
    .A2(_02369_),
    .A3(_02368_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21944_ (.A0(\design_top.MEM[15][19] ),
    .A1(\design_top.MEM[14][19] ),
    .A2(\design_top.MEM[13][19] ),
    .A3(\design_top.MEM[12][19] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21945_ (.A0(\design_top.MEM[11][19] ),
    .A1(\design_top.MEM[10][19] ),
    .A2(\design_top.MEM[9][19] ),
    .A3(\design_top.MEM[8][19] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21946_ (.A0(\design_top.MEM[7][19] ),
    .A1(\design_top.MEM[6][19] ),
    .A2(\design_top.MEM[5][19] ),
    .A3(\design_top.MEM[4][19] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21947_ (.A0(\design_top.MEM[3][19] ),
    .A1(\design_top.MEM[2][19] ),
    .A2(\design_top.MEM[1][19] ),
    .A3(\design_top.MEM[0][19] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21948_ (.A0(_02366_),
    .A1(_02365_),
    .A2(_02364_),
    .A3(_02363_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21949_ (.A0(_02382_),
    .A1(_02377_),
    .A2(_02372_),
    .A3(_02367_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21950_ (.A0(\design_top.MEM[63][18] ),
    .A1(\design_top.MEM[62][18] ),
    .A2(\design_top.MEM[61][18] ),
    .A3(\design_top.MEM[60][18] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21951_ (.A0(\design_top.MEM[59][18] ),
    .A1(\design_top.MEM[58][18] ),
    .A2(\design_top.MEM[57][18] ),
    .A3(\design_top.MEM[56][18] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21952_ (.A0(\design_top.MEM[55][18] ),
    .A1(\design_top.MEM[54][18] ),
    .A2(\design_top.MEM[53][18] ),
    .A3(\design_top.MEM[52][18] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21953_ (.A0(\design_top.MEM[51][18] ),
    .A1(\design_top.MEM[50][18] ),
    .A2(\design_top.MEM[49][18] ),
    .A3(\design_top.MEM[48][18] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21954_ (.A0(_02361_),
    .A1(_02360_),
    .A2(_02359_),
    .A3(_02358_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21955_ (.A0(\design_top.MEM[47][18] ),
    .A1(\design_top.MEM[46][18] ),
    .A2(\design_top.MEM[45][18] ),
    .A3(\design_top.MEM[44][18] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21956_ (.A0(\design_top.MEM[43][18] ),
    .A1(\design_top.MEM[42][18] ),
    .A2(\design_top.MEM[41][18] ),
    .A3(\design_top.MEM[40][18] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21957_ (.A0(\design_top.MEM[39][18] ),
    .A1(\design_top.MEM[38][18] ),
    .A2(\design_top.MEM[37][18] ),
    .A3(\design_top.MEM[36][18] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21958_ (.A0(\design_top.MEM[35][18] ),
    .A1(\design_top.MEM[34][18] ),
    .A2(\design_top.MEM[33][18] ),
    .A3(\design_top.MEM[32][18] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21959_ (.A0(_02356_),
    .A1(_02355_),
    .A2(_02354_),
    .A3(_02353_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21960_ (.A0(\design_top.MEM[31][18] ),
    .A1(\design_top.MEM[30][18] ),
    .A2(\design_top.MEM[29][18] ),
    .A3(\design_top.MEM[28][18] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21961_ (.A0(\design_top.MEM[27][18] ),
    .A1(\design_top.MEM[26][18] ),
    .A2(\design_top.MEM[25][18] ),
    .A3(\design_top.MEM[24][18] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21962_ (.A0(\design_top.MEM[23][18] ),
    .A1(\design_top.MEM[22][18] ),
    .A2(\design_top.MEM[21][18] ),
    .A3(\design_top.MEM[20][18] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21963_ (.A0(\design_top.MEM[19][18] ),
    .A1(\design_top.MEM[18][18] ),
    .A2(\design_top.MEM[17][18] ),
    .A3(\design_top.MEM[16][18] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21964_ (.A0(_02351_),
    .A1(_02350_),
    .A2(_02349_),
    .A3(_02348_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21965_ (.A0(\design_top.MEM[15][18] ),
    .A1(\design_top.MEM[14][18] ),
    .A2(\design_top.MEM[13][18] ),
    .A3(\design_top.MEM[12][18] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21966_ (.A0(\design_top.MEM[11][18] ),
    .A1(\design_top.MEM[10][18] ),
    .A2(\design_top.MEM[9][18] ),
    .A3(\design_top.MEM[8][18] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21967_ (.A0(\design_top.MEM[7][18] ),
    .A1(\design_top.MEM[6][18] ),
    .A2(\design_top.MEM[5][18] ),
    .A3(\design_top.MEM[4][18] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21968_ (.A0(\design_top.MEM[3][18] ),
    .A1(\design_top.MEM[2][18] ),
    .A2(\design_top.MEM[1][18] ),
    .A3(\design_top.MEM[0][18] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21969_ (.A0(_02346_),
    .A1(_02345_),
    .A2(_02344_),
    .A3(_02343_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21970_ (.A0(_02362_),
    .A1(_02357_),
    .A2(_02352_),
    .A3(_02347_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21971_ (.A0(\design_top.MEM[63][17] ),
    .A1(\design_top.MEM[62][17] ),
    .A2(\design_top.MEM[61][17] ),
    .A3(\design_top.MEM[60][17] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21972_ (.A0(\design_top.MEM[59][17] ),
    .A1(\design_top.MEM[58][17] ),
    .A2(\design_top.MEM[57][17] ),
    .A3(\design_top.MEM[56][17] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21973_ (.A0(\design_top.MEM[55][17] ),
    .A1(\design_top.MEM[54][17] ),
    .A2(\design_top.MEM[53][17] ),
    .A3(\design_top.MEM[52][17] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21974_ (.A0(\design_top.MEM[51][17] ),
    .A1(\design_top.MEM[50][17] ),
    .A2(\design_top.MEM[49][17] ),
    .A3(\design_top.MEM[48][17] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21975_ (.A0(_02341_),
    .A1(_02340_),
    .A2(_02339_),
    .A3(_02338_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21976_ (.A0(\design_top.MEM[47][17] ),
    .A1(\design_top.MEM[46][17] ),
    .A2(\design_top.MEM[45][17] ),
    .A3(\design_top.MEM[44][17] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21977_ (.A0(\design_top.MEM[43][17] ),
    .A1(\design_top.MEM[42][17] ),
    .A2(\design_top.MEM[41][17] ),
    .A3(\design_top.MEM[40][17] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21978_ (.A0(\design_top.MEM[39][17] ),
    .A1(\design_top.MEM[38][17] ),
    .A2(\design_top.MEM[37][17] ),
    .A3(\design_top.MEM[36][17] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21979_ (.A0(\design_top.MEM[35][17] ),
    .A1(\design_top.MEM[34][17] ),
    .A2(\design_top.MEM[33][17] ),
    .A3(\design_top.MEM[32][17] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21980_ (.A0(_02336_),
    .A1(_02335_),
    .A2(_02334_),
    .A3(_02333_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21981_ (.A0(\design_top.MEM[31][17] ),
    .A1(\design_top.MEM[30][17] ),
    .A2(\design_top.MEM[29][17] ),
    .A3(\design_top.MEM[28][17] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21982_ (.A0(\design_top.MEM[27][17] ),
    .A1(\design_top.MEM[26][17] ),
    .A2(\design_top.MEM[25][17] ),
    .A3(\design_top.MEM[24][17] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21983_ (.A0(\design_top.MEM[23][17] ),
    .A1(\design_top.MEM[22][17] ),
    .A2(\design_top.MEM[21][17] ),
    .A3(\design_top.MEM[20][17] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21984_ (.A0(\design_top.MEM[19][17] ),
    .A1(\design_top.MEM[18][17] ),
    .A2(\design_top.MEM[17][17] ),
    .A3(\design_top.MEM[16][17] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21985_ (.A0(_02331_),
    .A1(_02330_),
    .A2(_02329_),
    .A3(_02328_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21986_ (.A0(\design_top.MEM[15][17] ),
    .A1(\design_top.MEM[14][17] ),
    .A2(\design_top.MEM[13][17] ),
    .A3(\design_top.MEM[12][17] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21987_ (.A0(\design_top.MEM[11][17] ),
    .A1(\design_top.MEM[10][17] ),
    .A2(\design_top.MEM[9][17] ),
    .A3(\design_top.MEM[8][17] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21988_ (.A0(\design_top.MEM[7][17] ),
    .A1(\design_top.MEM[6][17] ),
    .A2(\design_top.MEM[5][17] ),
    .A3(\design_top.MEM[4][17] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21989_ (.A0(\design_top.MEM[3][17] ),
    .A1(\design_top.MEM[2][17] ),
    .A2(\design_top.MEM[1][17] ),
    .A3(\design_top.MEM[0][17] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21990_ (.A0(_02326_),
    .A1(_02325_),
    .A2(_02324_),
    .A3(_02323_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21991_ (.A0(_02342_),
    .A1(_02337_),
    .A2(_02332_),
    .A3(_02327_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21992_ (.A0(\design_top.MEM[63][16] ),
    .A1(\design_top.MEM[62][16] ),
    .A2(\design_top.MEM[61][16] ),
    .A3(\design_top.MEM[60][16] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21993_ (.A0(\design_top.MEM[59][16] ),
    .A1(\design_top.MEM[58][16] ),
    .A2(\design_top.MEM[57][16] ),
    .A3(\design_top.MEM[56][16] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21994_ (.A0(\design_top.MEM[55][16] ),
    .A1(\design_top.MEM[54][16] ),
    .A2(\design_top.MEM[53][16] ),
    .A3(\design_top.MEM[52][16] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21995_ (.A0(\design_top.MEM[51][16] ),
    .A1(\design_top.MEM[50][16] ),
    .A2(\design_top.MEM[49][16] ),
    .A3(\design_top.MEM[48][16] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21996_ (.A0(_02321_),
    .A1(_02320_),
    .A2(_02319_),
    .A3(_02318_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21997_ (.A0(\design_top.MEM[47][16] ),
    .A1(\design_top.MEM[46][16] ),
    .A2(\design_top.MEM[45][16] ),
    .A3(\design_top.MEM[44][16] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21998_ (.A0(\design_top.MEM[43][16] ),
    .A1(\design_top.MEM[42][16] ),
    .A2(\design_top.MEM[41][16] ),
    .A3(\design_top.MEM[40][16] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _21999_ (.A0(\design_top.MEM[39][16] ),
    .A1(\design_top.MEM[38][16] ),
    .A2(\design_top.MEM[37][16] ),
    .A3(\design_top.MEM[36][16] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22000_ (.A0(\design_top.MEM[35][16] ),
    .A1(\design_top.MEM[34][16] ),
    .A2(\design_top.MEM[33][16] ),
    .A3(\design_top.MEM[32][16] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22001_ (.A0(_02316_),
    .A1(_02315_),
    .A2(_02314_),
    .A3(_02313_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22002_ (.A0(\design_top.MEM[31][16] ),
    .A1(\design_top.MEM[30][16] ),
    .A2(\design_top.MEM[29][16] ),
    .A3(\design_top.MEM[28][16] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22003_ (.A0(\design_top.MEM[27][16] ),
    .A1(\design_top.MEM[26][16] ),
    .A2(\design_top.MEM[25][16] ),
    .A3(\design_top.MEM[24][16] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22004_ (.A0(\design_top.MEM[23][16] ),
    .A1(\design_top.MEM[22][16] ),
    .A2(\design_top.MEM[21][16] ),
    .A3(\design_top.MEM[20][16] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22005_ (.A0(\design_top.MEM[19][16] ),
    .A1(\design_top.MEM[18][16] ),
    .A2(\design_top.MEM[17][16] ),
    .A3(\design_top.MEM[16][16] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22006_ (.A0(_02311_),
    .A1(_02310_),
    .A2(_02309_),
    .A3(_02308_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22007_ (.A0(\design_top.MEM[15][16] ),
    .A1(\design_top.MEM[14][16] ),
    .A2(\design_top.MEM[13][16] ),
    .A3(\design_top.MEM[12][16] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22008_ (.A0(\design_top.MEM[11][16] ),
    .A1(\design_top.MEM[10][16] ),
    .A2(\design_top.MEM[9][16] ),
    .A3(\design_top.MEM[8][16] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22009_ (.A0(\design_top.MEM[7][16] ),
    .A1(\design_top.MEM[6][16] ),
    .A2(\design_top.MEM[5][16] ),
    .A3(\design_top.MEM[4][16] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22010_ (.A0(\design_top.MEM[3][16] ),
    .A1(\design_top.MEM[2][16] ),
    .A2(\design_top.MEM[1][16] ),
    .A3(\design_top.MEM[0][16] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22011_ (.A0(_02306_),
    .A1(_02305_),
    .A2(_02304_),
    .A3(_02303_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22012_ (.A0(_02322_),
    .A1(_02317_),
    .A2(_02312_),
    .A3(_02307_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22013_ (.A0(\design_top.MEM[63][15] ),
    .A1(\design_top.MEM[62][15] ),
    .A2(\design_top.MEM[61][15] ),
    .A3(\design_top.MEM[60][15] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22014_ (.A0(\design_top.MEM[59][15] ),
    .A1(\design_top.MEM[58][15] ),
    .A2(\design_top.MEM[57][15] ),
    .A3(\design_top.MEM[56][15] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22015_ (.A0(\design_top.MEM[55][15] ),
    .A1(\design_top.MEM[54][15] ),
    .A2(\design_top.MEM[53][15] ),
    .A3(\design_top.MEM[52][15] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22016_ (.A0(\design_top.MEM[51][15] ),
    .A1(\design_top.MEM[50][15] ),
    .A2(\design_top.MEM[49][15] ),
    .A3(\design_top.MEM[48][15] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22017_ (.A0(_02301_),
    .A1(_02300_),
    .A2(_02299_),
    .A3(_02298_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22018_ (.A0(\design_top.MEM[47][15] ),
    .A1(\design_top.MEM[46][15] ),
    .A2(\design_top.MEM[45][15] ),
    .A3(\design_top.MEM[44][15] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22019_ (.A0(\design_top.MEM[43][15] ),
    .A1(\design_top.MEM[42][15] ),
    .A2(\design_top.MEM[41][15] ),
    .A3(\design_top.MEM[40][15] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22020_ (.A0(\design_top.MEM[39][15] ),
    .A1(\design_top.MEM[38][15] ),
    .A2(\design_top.MEM[37][15] ),
    .A3(\design_top.MEM[36][15] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22021_ (.A0(\design_top.MEM[35][15] ),
    .A1(\design_top.MEM[34][15] ),
    .A2(\design_top.MEM[33][15] ),
    .A3(\design_top.MEM[32][15] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22022_ (.A0(_02296_),
    .A1(_02295_),
    .A2(_02294_),
    .A3(_02293_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22023_ (.A0(\design_top.MEM[31][15] ),
    .A1(\design_top.MEM[30][15] ),
    .A2(\design_top.MEM[29][15] ),
    .A3(\design_top.MEM[28][15] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22024_ (.A0(\design_top.MEM[27][15] ),
    .A1(\design_top.MEM[26][15] ),
    .A2(\design_top.MEM[25][15] ),
    .A3(\design_top.MEM[24][15] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22025_ (.A0(\design_top.MEM[23][15] ),
    .A1(\design_top.MEM[22][15] ),
    .A2(\design_top.MEM[21][15] ),
    .A3(\design_top.MEM[20][15] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22026_ (.A0(\design_top.MEM[19][15] ),
    .A1(\design_top.MEM[18][15] ),
    .A2(\design_top.MEM[17][15] ),
    .A3(\design_top.MEM[16][15] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22027_ (.A0(_02291_),
    .A1(_02290_),
    .A2(_02289_),
    .A3(_02288_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22028_ (.A0(\design_top.MEM[15][15] ),
    .A1(\design_top.MEM[14][15] ),
    .A2(\design_top.MEM[13][15] ),
    .A3(\design_top.MEM[12][15] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22029_ (.A0(\design_top.MEM[11][15] ),
    .A1(\design_top.MEM[10][15] ),
    .A2(\design_top.MEM[9][15] ),
    .A3(\design_top.MEM[8][15] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22030_ (.A0(\design_top.MEM[7][15] ),
    .A1(\design_top.MEM[6][15] ),
    .A2(\design_top.MEM[5][15] ),
    .A3(\design_top.MEM[4][15] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22031_ (.A0(\design_top.MEM[3][15] ),
    .A1(\design_top.MEM[2][15] ),
    .A2(\design_top.MEM[1][15] ),
    .A3(\design_top.MEM[0][15] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22032_ (.A0(_02286_),
    .A1(_02285_),
    .A2(_02284_),
    .A3(_02283_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22033_ (.A0(_02302_),
    .A1(_02297_),
    .A2(_02292_),
    .A3(_02287_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22034_ (.A0(\design_top.MEM[63][14] ),
    .A1(\design_top.MEM[62][14] ),
    .A2(\design_top.MEM[61][14] ),
    .A3(\design_top.MEM[60][14] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22035_ (.A0(\design_top.MEM[59][14] ),
    .A1(\design_top.MEM[58][14] ),
    .A2(\design_top.MEM[57][14] ),
    .A3(\design_top.MEM[56][14] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22036_ (.A0(\design_top.MEM[55][14] ),
    .A1(\design_top.MEM[54][14] ),
    .A2(\design_top.MEM[53][14] ),
    .A3(\design_top.MEM[52][14] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22037_ (.A0(\design_top.MEM[51][14] ),
    .A1(\design_top.MEM[50][14] ),
    .A2(\design_top.MEM[49][14] ),
    .A3(\design_top.MEM[48][14] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22038_ (.A0(_02281_),
    .A1(_02280_),
    .A2(_02279_),
    .A3(_02278_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22039_ (.A0(\design_top.MEM[47][14] ),
    .A1(\design_top.MEM[46][14] ),
    .A2(\design_top.MEM[45][14] ),
    .A3(\design_top.MEM[44][14] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22040_ (.A0(\design_top.MEM[43][14] ),
    .A1(\design_top.MEM[42][14] ),
    .A2(\design_top.MEM[41][14] ),
    .A3(\design_top.MEM[40][14] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22041_ (.A0(\design_top.MEM[39][14] ),
    .A1(\design_top.MEM[38][14] ),
    .A2(\design_top.MEM[37][14] ),
    .A3(\design_top.MEM[36][14] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22042_ (.A0(\design_top.MEM[35][14] ),
    .A1(\design_top.MEM[34][14] ),
    .A2(\design_top.MEM[33][14] ),
    .A3(\design_top.MEM[32][14] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22043_ (.A0(_02276_),
    .A1(_02275_),
    .A2(_02274_),
    .A3(_02273_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22044_ (.A0(\design_top.MEM[31][14] ),
    .A1(\design_top.MEM[30][14] ),
    .A2(\design_top.MEM[29][14] ),
    .A3(\design_top.MEM[28][14] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22045_ (.A0(\design_top.MEM[27][14] ),
    .A1(\design_top.MEM[26][14] ),
    .A2(\design_top.MEM[25][14] ),
    .A3(\design_top.MEM[24][14] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22046_ (.A0(\design_top.MEM[23][14] ),
    .A1(\design_top.MEM[22][14] ),
    .A2(\design_top.MEM[21][14] ),
    .A3(\design_top.MEM[20][14] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22047_ (.A0(\design_top.MEM[19][14] ),
    .A1(\design_top.MEM[18][14] ),
    .A2(\design_top.MEM[17][14] ),
    .A3(\design_top.MEM[16][14] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22048_ (.A0(_02271_),
    .A1(_02270_),
    .A2(_02269_),
    .A3(_02268_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22049_ (.A0(\design_top.MEM[15][14] ),
    .A1(\design_top.MEM[14][14] ),
    .A2(\design_top.MEM[13][14] ),
    .A3(\design_top.MEM[12][14] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22050_ (.A0(\design_top.MEM[11][14] ),
    .A1(\design_top.MEM[10][14] ),
    .A2(\design_top.MEM[9][14] ),
    .A3(\design_top.MEM[8][14] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22051_ (.A0(\design_top.MEM[7][14] ),
    .A1(\design_top.MEM[6][14] ),
    .A2(\design_top.MEM[5][14] ),
    .A3(\design_top.MEM[4][14] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22052_ (.A0(\design_top.MEM[3][14] ),
    .A1(\design_top.MEM[2][14] ),
    .A2(\design_top.MEM[1][14] ),
    .A3(\design_top.MEM[0][14] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22053_ (.A0(_02266_),
    .A1(_02265_),
    .A2(_02264_),
    .A3(_02263_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22054_ (.A0(_02282_),
    .A1(_02277_),
    .A2(_02272_),
    .A3(_02267_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22055_ (.A0(\design_top.MEM[63][13] ),
    .A1(\design_top.MEM[62][13] ),
    .A2(\design_top.MEM[61][13] ),
    .A3(\design_top.MEM[60][13] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22056_ (.A0(\design_top.MEM[59][13] ),
    .A1(\design_top.MEM[58][13] ),
    .A2(\design_top.MEM[57][13] ),
    .A3(\design_top.MEM[56][13] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22057_ (.A0(\design_top.MEM[55][13] ),
    .A1(\design_top.MEM[54][13] ),
    .A2(\design_top.MEM[53][13] ),
    .A3(\design_top.MEM[52][13] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22058_ (.A0(\design_top.MEM[51][13] ),
    .A1(\design_top.MEM[50][13] ),
    .A2(\design_top.MEM[49][13] ),
    .A3(\design_top.MEM[48][13] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22059_ (.A0(_02261_),
    .A1(_02260_),
    .A2(_02259_),
    .A3(_02258_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22060_ (.A0(\design_top.MEM[47][13] ),
    .A1(\design_top.MEM[46][13] ),
    .A2(\design_top.MEM[45][13] ),
    .A3(\design_top.MEM[44][13] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22061_ (.A0(\design_top.MEM[43][13] ),
    .A1(\design_top.MEM[42][13] ),
    .A2(\design_top.MEM[41][13] ),
    .A3(\design_top.MEM[40][13] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22062_ (.A0(\design_top.MEM[39][13] ),
    .A1(\design_top.MEM[38][13] ),
    .A2(\design_top.MEM[37][13] ),
    .A3(\design_top.MEM[36][13] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22063_ (.A0(\design_top.MEM[35][13] ),
    .A1(\design_top.MEM[34][13] ),
    .A2(\design_top.MEM[33][13] ),
    .A3(\design_top.MEM[32][13] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22064_ (.A0(_02256_),
    .A1(_02255_),
    .A2(_02254_),
    .A3(_02253_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22065_ (.A0(\design_top.MEM[31][13] ),
    .A1(\design_top.MEM[30][13] ),
    .A2(\design_top.MEM[29][13] ),
    .A3(\design_top.MEM[28][13] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22066_ (.A0(\design_top.MEM[27][13] ),
    .A1(\design_top.MEM[26][13] ),
    .A2(\design_top.MEM[25][13] ),
    .A3(\design_top.MEM[24][13] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22067_ (.A0(\design_top.MEM[23][13] ),
    .A1(\design_top.MEM[22][13] ),
    .A2(\design_top.MEM[21][13] ),
    .A3(\design_top.MEM[20][13] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22068_ (.A0(\design_top.MEM[19][13] ),
    .A1(\design_top.MEM[18][13] ),
    .A2(\design_top.MEM[17][13] ),
    .A3(\design_top.MEM[16][13] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22069_ (.A0(_02251_),
    .A1(_02250_),
    .A2(_02249_),
    .A3(_02248_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22070_ (.A0(\design_top.MEM[15][13] ),
    .A1(\design_top.MEM[14][13] ),
    .A2(\design_top.MEM[13][13] ),
    .A3(\design_top.MEM[12][13] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22071_ (.A0(\design_top.MEM[11][13] ),
    .A1(\design_top.MEM[10][13] ),
    .A2(\design_top.MEM[9][13] ),
    .A3(\design_top.MEM[8][13] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22072_ (.A0(\design_top.MEM[7][13] ),
    .A1(\design_top.MEM[6][13] ),
    .A2(\design_top.MEM[5][13] ),
    .A3(\design_top.MEM[4][13] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22073_ (.A0(\design_top.MEM[3][13] ),
    .A1(\design_top.MEM[2][13] ),
    .A2(\design_top.MEM[1][13] ),
    .A3(\design_top.MEM[0][13] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22074_ (.A0(_02246_),
    .A1(_02245_),
    .A2(_02244_),
    .A3(_02243_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22075_ (.A0(_02262_),
    .A1(_02257_),
    .A2(_02252_),
    .A3(_02247_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22076_ (.A0(\design_top.MEM[63][12] ),
    .A1(\design_top.MEM[62][12] ),
    .A2(\design_top.MEM[61][12] ),
    .A3(\design_top.MEM[60][12] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22077_ (.A0(\design_top.MEM[59][12] ),
    .A1(\design_top.MEM[58][12] ),
    .A2(\design_top.MEM[57][12] ),
    .A3(\design_top.MEM[56][12] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22078_ (.A0(\design_top.MEM[55][12] ),
    .A1(\design_top.MEM[54][12] ),
    .A2(\design_top.MEM[53][12] ),
    .A3(\design_top.MEM[52][12] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22079_ (.A0(\design_top.MEM[51][12] ),
    .A1(\design_top.MEM[50][12] ),
    .A2(\design_top.MEM[49][12] ),
    .A3(\design_top.MEM[48][12] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22080_ (.A0(_02241_),
    .A1(_02240_),
    .A2(_02239_),
    .A3(_02238_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22081_ (.A0(\design_top.MEM[47][12] ),
    .A1(\design_top.MEM[46][12] ),
    .A2(\design_top.MEM[45][12] ),
    .A3(\design_top.MEM[44][12] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22082_ (.A0(\design_top.MEM[43][12] ),
    .A1(\design_top.MEM[42][12] ),
    .A2(\design_top.MEM[41][12] ),
    .A3(\design_top.MEM[40][12] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22083_ (.A0(\design_top.MEM[39][12] ),
    .A1(\design_top.MEM[38][12] ),
    .A2(\design_top.MEM[37][12] ),
    .A3(\design_top.MEM[36][12] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22084_ (.A0(\design_top.MEM[35][12] ),
    .A1(\design_top.MEM[34][12] ),
    .A2(\design_top.MEM[33][12] ),
    .A3(\design_top.MEM[32][12] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22085_ (.A0(_02236_),
    .A1(_02235_),
    .A2(_02234_),
    .A3(_02233_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22086_ (.A0(\design_top.MEM[31][12] ),
    .A1(\design_top.MEM[30][12] ),
    .A2(\design_top.MEM[29][12] ),
    .A3(\design_top.MEM[28][12] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22087_ (.A0(\design_top.MEM[27][12] ),
    .A1(\design_top.MEM[26][12] ),
    .A2(\design_top.MEM[25][12] ),
    .A3(\design_top.MEM[24][12] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22088_ (.A0(\design_top.MEM[23][12] ),
    .A1(\design_top.MEM[22][12] ),
    .A2(\design_top.MEM[21][12] ),
    .A3(\design_top.MEM[20][12] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22089_ (.A0(\design_top.MEM[19][12] ),
    .A1(\design_top.MEM[18][12] ),
    .A2(\design_top.MEM[17][12] ),
    .A3(\design_top.MEM[16][12] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22090_ (.A0(_02231_),
    .A1(_02230_),
    .A2(_02229_),
    .A3(_02228_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22091_ (.A0(\design_top.MEM[15][12] ),
    .A1(\design_top.MEM[14][12] ),
    .A2(\design_top.MEM[13][12] ),
    .A3(\design_top.MEM[12][12] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22092_ (.A0(\design_top.MEM[11][12] ),
    .A1(\design_top.MEM[10][12] ),
    .A2(\design_top.MEM[9][12] ),
    .A3(\design_top.MEM[8][12] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22093_ (.A0(\design_top.MEM[7][12] ),
    .A1(\design_top.MEM[6][12] ),
    .A2(\design_top.MEM[5][12] ),
    .A3(\design_top.MEM[4][12] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22094_ (.A0(\design_top.MEM[3][12] ),
    .A1(\design_top.MEM[2][12] ),
    .A2(\design_top.MEM[1][12] ),
    .A3(\design_top.MEM[0][12] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22095_ (.A0(_02226_),
    .A1(_02225_),
    .A2(_02224_),
    .A3(_02223_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22096_ (.A0(_02242_),
    .A1(_02237_),
    .A2(_02232_),
    .A3(_02227_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22097_ (.A0(\design_top.MEM[63][11] ),
    .A1(\design_top.MEM[62][11] ),
    .A2(\design_top.MEM[61][11] ),
    .A3(\design_top.MEM[60][11] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22098_ (.A0(\design_top.MEM[59][11] ),
    .A1(\design_top.MEM[58][11] ),
    .A2(\design_top.MEM[57][11] ),
    .A3(\design_top.MEM[56][11] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22099_ (.A0(\design_top.MEM[55][11] ),
    .A1(\design_top.MEM[54][11] ),
    .A2(\design_top.MEM[53][11] ),
    .A3(\design_top.MEM[52][11] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22100_ (.A0(\design_top.MEM[51][11] ),
    .A1(\design_top.MEM[50][11] ),
    .A2(\design_top.MEM[49][11] ),
    .A3(\design_top.MEM[48][11] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22101_ (.A0(_02221_),
    .A1(_02220_),
    .A2(_02219_),
    .A3(_02218_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22102_ (.A0(\design_top.MEM[47][11] ),
    .A1(\design_top.MEM[46][11] ),
    .A2(\design_top.MEM[45][11] ),
    .A3(\design_top.MEM[44][11] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22103_ (.A0(\design_top.MEM[43][11] ),
    .A1(\design_top.MEM[42][11] ),
    .A2(\design_top.MEM[41][11] ),
    .A3(\design_top.MEM[40][11] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22104_ (.A0(\design_top.MEM[39][11] ),
    .A1(\design_top.MEM[38][11] ),
    .A2(\design_top.MEM[37][11] ),
    .A3(\design_top.MEM[36][11] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22105_ (.A0(\design_top.MEM[35][11] ),
    .A1(\design_top.MEM[34][11] ),
    .A2(\design_top.MEM[33][11] ),
    .A3(\design_top.MEM[32][11] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22106_ (.A0(_02216_),
    .A1(_02215_),
    .A2(_02214_),
    .A3(_02213_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22107_ (.A0(\design_top.MEM[31][11] ),
    .A1(\design_top.MEM[30][11] ),
    .A2(\design_top.MEM[29][11] ),
    .A3(\design_top.MEM[28][11] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22108_ (.A0(\design_top.MEM[27][11] ),
    .A1(\design_top.MEM[26][11] ),
    .A2(\design_top.MEM[25][11] ),
    .A3(\design_top.MEM[24][11] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22109_ (.A0(\design_top.MEM[23][11] ),
    .A1(\design_top.MEM[22][11] ),
    .A2(\design_top.MEM[21][11] ),
    .A3(\design_top.MEM[20][11] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22110_ (.A0(\design_top.MEM[19][11] ),
    .A1(\design_top.MEM[18][11] ),
    .A2(\design_top.MEM[17][11] ),
    .A3(\design_top.MEM[16][11] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22111_ (.A0(_02211_),
    .A1(_02210_),
    .A2(_02209_),
    .A3(_02208_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22112_ (.A0(\design_top.MEM[15][11] ),
    .A1(\design_top.MEM[14][11] ),
    .A2(\design_top.MEM[13][11] ),
    .A3(\design_top.MEM[12][11] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22113_ (.A0(\design_top.MEM[11][11] ),
    .A1(\design_top.MEM[10][11] ),
    .A2(\design_top.MEM[9][11] ),
    .A3(\design_top.MEM[8][11] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22114_ (.A0(\design_top.MEM[7][11] ),
    .A1(\design_top.MEM[6][11] ),
    .A2(\design_top.MEM[5][11] ),
    .A3(\design_top.MEM[4][11] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22115_ (.A0(\design_top.MEM[3][11] ),
    .A1(\design_top.MEM[2][11] ),
    .A2(\design_top.MEM[1][11] ),
    .A3(\design_top.MEM[0][11] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22116_ (.A0(_02206_),
    .A1(_02205_),
    .A2(_02204_),
    .A3(_02203_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22117_ (.A0(_02222_),
    .A1(_02217_),
    .A2(_02212_),
    .A3(_02207_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22118_ (.A0(\design_top.MEM[63][10] ),
    .A1(\design_top.MEM[62][10] ),
    .A2(\design_top.MEM[61][10] ),
    .A3(\design_top.MEM[60][10] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22119_ (.A0(\design_top.MEM[59][10] ),
    .A1(\design_top.MEM[58][10] ),
    .A2(\design_top.MEM[57][10] ),
    .A3(\design_top.MEM[56][10] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22120_ (.A0(\design_top.MEM[55][10] ),
    .A1(\design_top.MEM[54][10] ),
    .A2(\design_top.MEM[53][10] ),
    .A3(\design_top.MEM[52][10] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22121_ (.A0(\design_top.MEM[51][10] ),
    .A1(\design_top.MEM[50][10] ),
    .A2(\design_top.MEM[49][10] ),
    .A3(\design_top.MEM[48][10] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22122_ (.A0(_02201_),
    .A1(_02200_),
    .A2(_02199_),
    .A3(_02198_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22123_ (.A0(\design_top.MEM[47][10] ),
    .A1(\design_top.MEM[46][10] ),
    .A2(\design_top.MEM[45][10] ),
    .A3(\design_top.MEM[44][10] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22124_ (.A0(\design_top.MEM[43][10] ),
    .A1(\design_top.MEM[42][10] ),
    .A2(\design_top.MEM[41][10] ),
    .A3(\design_top.MEM[40][10] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22125_ (.A0(\design_top.MEM[39][10] ),
    .A1(\design_top.MEM[38][10] ),
    .A2(\design_top.MEM[37][10] ),
    .A3(\design_top.MEM[36][10] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22126_ (.A0(\design_top.MEM[35][10] ),
    .A1(\design_top.MEM[34][10] ),
    .A2(\design_top.MEM[33][10] ),
    .A3(\design_top.MEM[32][10] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22127_ (.A0(_02196_),
    .A1(_02195_),
    .A2(_02194_),
    .A3(_02193_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22128_ (.A0(\design_top.MEM[31][10] ),
    .A1(\design_top.MEM[30][10] ),
    .A2(\design_top.MEM[29][10] ),
    .A3(\design_top.MEM[28][10] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22129_ (.A0(\design_top.MEM[27][10] ),
    .A1(\design_top.MEM[26][10] ),
    .A2(\design_top.MEM[25][10] ),
    .A3(\design_top.MEM[24][10] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22130_ (.A0(\design_top.MEM[23][10] ),
    .A1(\design_top.MEM[22][10] ),
    .A2(\design_top.MEM[21][10] ),
    .A3(\design_top.MEM[20][10] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22131_ (.A0(\design_top.MEM[19][10] ),
    .A1(\design_top.MEM[18][10] ),
    .A2(\design_top.MEM[17][10] ),
    .A3(\design_top.MEM[16][10] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22132_ (.A0(_02191_),
    .A1(_02190_),
    .A2(_02189_),
    .A3(_02188_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22133_ (.A0(\design_top.MEM[15][10] ),
    .A1(\design_top.MEM[14][10] ),
    .A2(\design_top.MEM[13][10] ),
    .A3(\design_top.MEM[12][10] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22134_ (.A0(\design_top.MEM[11][10] ),
    .A1(\design_top.MEM[10][10] ),
    .A2(\design_top.MEM[9][10] ),
    .A3(\design_top.MEM[8][10] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22135_ (.A0(\design_top.MEM[7][10] ),
    .A1(\design_top.MEM[6][10] ),
    .A2(\design_top.MEM[5][10] ),
    .A3(\design_top.MEM[4][10] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22136_ (.A0(\design_top.MEM[3][10] ),
    .A1(\design_top.MEM[2][10] ),
    .A2(\design_top.MEM[1][10] ),
    .A3(\design_top.MEM[0][10] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22137_ (.A0(_02186_),
    .A1(_02185_),
    .A2(_02184_),
    .A3(_02183_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22138_ (.A0(_02202_),
    .A1(_02197_),
    .A2(_02192_),
    .A3(_02187_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22139_ (.A0(\design_top.MEM[63][9] ),
    .A1(\design_top.MEM[62][9] ),
    .A2(\design_top.MEM[61][9] ),
    .A3(\design_top.MEM[60][9] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22140_ (.A0(\design_top.MEM[59][9] ),
    .A1(\design_top.MEM[58][9] ),
    .A2(\design_top.MEM[57][9] ),
    .A3(\design_top.MEM[56][9] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22141_ (.A0(\design_top.MEM[55][9] ),
    .A1(\design_top.MEM[54][9] ),
    .A2(\design_top.MEM[53][9] ),
    .A3(\design_top.MEM[52][9] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22142_ (.A0(\design_top.MEM[51][9] ),
    .A1(\design_top.MEM[50][9] ),
    .A2(\design_top.MEM[49][9] ),
    .A3(\design_top.MEM[48][9] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22143_ (.A0(_02181_),
    .A1(_02180_),
    .A2(_02179_),
    .A3(_02178_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22144_ (.A0(\design_top.MEM[47][9] ),
    .A1(\design_top.MEM[46][9] ),
    .A2(\design_top.MEM[45][9] ),
    .A3(\design_top.MEM[44][9] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22145_ (.A0(\design_top.MEM[43][9] ),
    .A1(\design_top.MEM[42][9] ),
    .A2(\design_top.MEM[41][9] ),
    .A3(\design_top.MEM[40][9] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22146_ (.A0(\design_top.MEM[39][9] ),
    .A1(\design_top.MEM[38][9] ),
    .A2(\design_top.MEM[37][9] ),
    .A3(\design_top.MEM[36][9] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22147_ (.A0(\design_top.MEM[35][9] ),
    .A1(\design_top.MEM[34][9] ),
    .A2(\design_top.MEM[33][9] ),
    .A3(\design_top.MEM[32][9] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22148_ (.A0(_02176_),
    .A1(_02175_),
    .A2(_02174_),
    .A3(_02173_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22149_ (.A0(\design_top.MEM[31][9] ),
    .A1(\design_top.MEM[30][9] ),
    .A2(\design_top.MEM[29][9] ),
    .A3(\design_top.MEM[28][9] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22150_ (.A0(\design_top.MEM[27][9] ),
    .A1(\design_top.MEM[26][9] ),
    .A2(\design_top.MEM[25][9] ),
    .A3(\design_top.MEM[24][9] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22151_ (.A0(\design_top.MEM[23][9] ),
    .A1(\design_top.MEM[22][9] ),
    .A2(\design_top.MEM[21][9] ),
    .A3(\design_top.MEM[20][9] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22152_ (.A0(\design_top.MEM[19][9] ),
    .A1(\design_top.MEM[18][9] ),
    .A2(\design_top.MEM[17][9] ),
    .A3(\design_top.MEM[16][9] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22153_ (.A0(_02171_),
    .A1(_02170_),
    .A2(_02169_),
    .A3(_02168_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22154_ (.A0(\design_top.MEM[15][9] ),
    .A1(\design_top.MEM[14][9] ),
    .A2(\design_top.MEM[13][9] ),
    .A3(\design_top.MEM[12][9] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22155_ (.A0(\design_top.MEM[11][9] ),
    .A1(\design_top.MEM[10][9] ),
    .A2(\design_top.MEM[9][9] ),
    .A3(\design_top.MEM[8][9] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22156_ (.A0(\design_top.MEM[7][9] ),
    .A1(\design_top.MEM[6][9] ),
    .A2(\design_top.MEM[5][9] ),
    .A3(\design_top.MEM[4][9] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22157_ (.A0(\design_top.MEM[3][9] ),
    .A1(\design_top.MEM[2][9] ),
    .A2(\design_top.MEM[1][9] ),
    .A3(\design_top.MEM[0][9] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22158_ (.A0(_02166_),
    .A1(_02165_),
    .A2(_02164_),
    .A3(_02163_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22159_ (.A0(_02182_),
    .A1(_02177_),
    .A2(_02172_),
    .A3(_02167_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22160_ (.A0(\design_top.MEM[63][8] ),
    .A1(\design_top.MEM[62][8] ),
    .A2(\design_top.MEM[61][8] ),
    .A3(\design_top.MEM[60][8] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22161_ (.A0(\design_top.MEM[59][8] ),
    .A1(\design_top.MEM[58][8] ),
    .A2(\design_top.MEM[57][8] ),
    .A3(\design_top.MEM[56][8] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22162_ (.A0(\design_top.MEM[55][8] ),
    .A1(\design_top.MEM[54][8] ),
    .A2(\design_top.MEM[53][8] ),
    .A3(\design_top.MEM[52][8] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22163_ (.A0(\design_top.MEM[51][8] ),
    .A1(\design_top.MEM[50][8] ),
    .A2(\design_top.MEM[49][8] ),
    .A3(\design_top.MEM[48][8] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22164_ (.A0(_02161_),
    .A1(_02160_),
    .A2(_02159_),
    .A3(_02158_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22165_ (.A0(\design_top.MEM[47][8] ),
    .A1(\design_top.MEM[46][8] ),
    .A2(\design_top.MEM[45][8] ),
    .A3(\design_top.MEM[44][8] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22166_ (.A0(\design_top.MEM[43][8] ),
    .A1(\design_top.MEM[42][8] ),
    .A2(\design_top.MEM[41][8] ),
    .A3(\design_top.MEM[40][8] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22167_ (.A0(\design_top.MEM[39][8] ),
    .A1(\design_top.MEM[38][8] ),
    .A2(\design_top.MEM[37][8] ),
    .A3(\design_top.MEM[36][8] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22168_ (.A0(\design_top.MEM[35][8] ),
    .A1(\design_top.MEM[34][8] ),
    .A2(\design_top.MEM[33][8] ),
    .A3(\design_top.MEM[32][8] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22169_ (.A0(_02156_),
    .A1(_02155_),
    .A2(_02154_),
    .A3(_02153_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22170_ (.A0(\design_top.MEM[31][8] ),
    .A1(\design_top.MEM[30][8] ),
    .A2(\design_top.MEM[29][8] ),
    .A3(\design_top.MEM[28][8] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22171_ (.A0(\design_top.MEM[27][8] ),
    .A1(\design_top.MEM[26][8] ),
    .A2(\design_top.MEM[25][8] ),
    .A3(\design_top.MEM[24][8] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22172_ (.A0(\design_top.MEM[23][8] ),
    .A1(\design_top.MEM[22][8] ),
    .A2(\design_top.MEM[21][8] ),
    .A3(\design_top.MEM[20][8] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22173_ (.A0(\design_top.MEM[19][8] ),
    .A1(\design_top.MEM[18][8] ),
    .A2(\design_top.MEM[17][8] ),
    .A3(\design_top.MEM[16][8] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22174_ (.A0(_02151_),
    .A1(_02150_),
    .A2(_02149_),
    .A3(_02148_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22175_ (.A0(\design_top.MEM[15][8] ),
    .A1(\design_top.MEM[14][8] ),
    .A2(\design_top.MEM[13][8] ),
    .A3(\design_top.MEM[12][8] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22176_ (.A0(\design_top.MEM[11][8] ),
    .A1(\design_top.MEM[10][8] ),
    .A2(\design_top.MEM[9][8] ),
    .A3(\design_top.MEM[8][8] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22177_ (.A0(\design_top.MEM[7][8] ),
    .A1(\design_top.MEM[6][8] ),
    .A2(\design_top.MEM[5][8] ),
    .A3(\design_top.MEM[4][8] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22178_ (.A0(\design_top.MEM[3][8] ),
    .A1(\design_top.MEM[2][8] ),
    .A2(\design_top.MEM[1][8] ),
    .A3(\design_top.MEM[0][8] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22179_ (.A0(_02146_),
    .A1(_02145_),
    .A2(_02144_),
    .A3(_02143_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22180_ (.A0(_02162_),
    .A1(_02157_),
    .A2(_02152_),
    .A3(_02147_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22181_ (.A0(\design_top.MEM[63][7] ),
    .A1(\design_top.MEM[62][7] ),
    .A2(\design_top.MEM[61][7] ),
    .A3(\design_top.MEM[60][7] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22182_ (.A0(\design_top.MEM[59][7] ),
    .A1(\design_top.MEM[58][7] ),
    .A2(\design_top.MEM[57][7] ),
    .A3(\design_top.MEM[56][7] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22183_ (.A0(\design_top.MEM[55][7] ),
    .A1(\design_top.MEM[54][7] ),
    .A2(\design_top.MEM[53][7] ),
    .A3(\design_top.MEM[52][7] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22184_ (.A0(\design_top.MEM[51][7] ),
    .A1(\design_top.MEM[50][7] ),
    .A2(\design_top.MEM[49][7] ),
    .A3(\design_top.MEM[48][7] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22185_ (.A0(_02141_),
    .A1(_02140_),
    .A2(_02139_),
    .A3(_02138_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22186_ (.A0(\design_top.MEM[47][7] ),
    .A1(\design_top.MEM[46][7] ),
    .A2(\design_top.MEM[45][7] ),
    .A3(\design_top.MEM[44][7] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22187_ (.A0(\design_top.MEM[43][7] ),
    .A1(\design_top.MEM[42][7] ),
    .A2(\design_top.MEM[41][7] ),
    .A3(\design_top.MEM[40][7] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22188_ (.A0(\design_top.MEM[39][7] ),
    .A1(\design_top.MEM[38][7] ),
    .A2(\design_top.MEM[37][7] ),
    .A3(\design_top.MEM[36][7] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22189_ (.A0(\design_top.MEM[35][7] ),
    .A1(\design_top.MEM[34][7] ),
    .A2(\design_top.MEM[33][7] ),
    .A3(\design_top.MEM[32][7] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22190_ (.A0(_02136_),
    .A1(_02135_),
    .A2(_02134_),
    .A3(_02133_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22191_ (.A0(\design_top.MEM[31][7] ),
    .A1(\design_top.MEM[30][7] ),
    .A2(\design_top.MEM[29][7] ),
    .A3(\design_top.MEM[28][7] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22192_ (.A0(\design_top.MEM[27][7] ),
    .A1(\design_top.MEM[26][7] ),
    .A2(\design_top.MEM[25][7] ),
    .A3(\design_top.MEM[24][7] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22193_ (.A0(\design_top.MEM[23][7] ),
    .A1(\design_top.MEM[22][7] ),
    .A2(\design_top.MEM[21][7] ),
    .A3(\design_top.MEM[20][7] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22194_ (.A0(\design_top.MEM[19][7] ),
    .A1(\design_top.MEM[18][7] ),
    .A2(\design_top.MEM[17][7] ),
    .A3(\design_top.MEM[16][7] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22195_ (.A0(_02131_),
    .A1(_02130_),
    .A2(_02129_),
    .A3(_02128_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22196_ (.A0(\design_top.MEM[15][7] ),
    .A1(\design_top.MEM[14][7] ),
    .A2(\design_top.MEM[13][7] ),
    .A3(\design_top.MEM[12][7] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22197_ (.A0(\design_top.MEM[11][7] ),
    .A1(\design_top.MEM[10][7] ),
    .A2(\design_top.MEM[9][7] ),
    .A3(\design_top.MEM[8][7] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22198_ (.A0(\design_top.MEM[7][7] ),
    .A1(\design_top.MEM[6][7] ),
    .A2(\design_top.MEM[5][7] ),
    .A3(\design_top.MEM[4][7] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22199_ (.A0(\design_top.MEM[3][7] ),
    .A1(\design_top.MEM[2][7] ),
    .A2(\design_top.MEM[1][7] ),
    .A3(\design_top.MEM[0][7] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22200_ (.A0(_02126_),
    .A1(_02125_),
    .A2(_02124_),
    .A3(_02123_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22201_ (.A0(_02142_),
    .A1(_02137_),
    .A2(_02132_),
    .A3(_02127_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22202_ (.A0(\design_top.MEM[63][6] ),
    .A1(\design_top.MEM[62][6] ),
    .A2(\design_top.MEM[61][6] ),
    .A3(\design_top.MEM[60][6] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22203_ (.A0(\design_top.MEM[59][6] ),
    .A1(\design_top.MEM[58][6] ),
    .A2(\design_top.MEM[57][6] ),
    .A3(\design_top.MEM[56][6] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22204_ (.A0(\design_top.MEM[55][6] ),
    .A1(\design_top.MEM[54][6] ),
    .A2(\design_top.MEM[53][6] ),
    .A3(\design_top.MEM[52][6] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22205_ (.A0(\design_top.MEM[51][6] ),
    .A1(\design_top.MEM[50][6] ),
    .A2(\design_top.MEM[49][6] ),
    .A3(\design_top.MEM[48][6] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22206_ (.A0(_02121_),
    .A1(_02120_),
    .A2(_02119_),
    .A3(_02118_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22207_ (.A0(\design_top.MEM[47][6] ),
    .A1(\design_top.MEM[46][6] ),
    .A2(\design_top.MEM[45][6] ),
    .A3(\design_top.MEM[44][6] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22208_ (.A0(\design_top.MEM[43][6] ),
    .A1(\design_top.MEM[42][6] ),
    .A2(\design_top.MEM[41][6] ),
    .A3(\design_top.MEM[40][6] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22209_ (.A0(\design_top.MEM[39][6] ),
    .A1(\design_top.MEM[38][6] ),
    .A2(\design_top.MEM[37][6] ),
    .A3(\design_top.MEM[36][6] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22210_ (.A0(\design_top.MEM[35][6] ),
    .A1(\design_top.MEM[34][6] ),
    .A2(\design_top.MEM[33][6] ),
    .A3(\design_top.MEM[32][6] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22211_ (.A0(_02116_),
    .A1(_02115_),
    .A2(_02114_),
    .A3(_02113_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22212_ (.A0(\design_top.MEM[31][6] ),
    .A1(\design_top.MEM[30][6] ),
    .A2(\design_top.MEM[29][6] ),
    .A3(\design_top.MEM[28][6] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22213_ (.A0(\design_top.MEM[27][6] ),
    .A1(\design_top.MEM[26][6] ),
    .A2(\design_top.MEM[25][6] ),
    .A3(\design_top.MEM[24][6] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22214_ (.A0(\design_top.MEM[23][6] ),
    .A1(\design_top.MEM[22][6] ),
    .A2(\design_top.MEM[21][6] ),
    .A3(\design_top.MEM[20][6] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22215_ (.A0(\design_top.MEM[19][6] ),
    .A1(\design_top.MEM[18][6] ),
    .A2(\design_top.MEM[17][6] ),
    .A3(\design_top.MEM[16][6] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22216_ (.A0(_02111_),
    .A1(_02110_),
    .A2(_02109_),
    .A3(_02108_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22217_ (.A0(\design_top.MEM[15][6] ),
    .A1(\design_top.MEM[14][6] ),
    .A2(\design_top.MEM[13][6] ),
    .A3(\design_top.MEM[12][6] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22218_ (.A0(\design_top.MEM[11][6] ),
    .A1(\design_top.MEM[10][6] ),
    .A2(\design_top.MEM[9][6] ),
    .A3(\design_top.MEM[8][6] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22219_ (.A0(\design_top.MEM[7][6] ),
    .A1(\design_top.MEM[6][6] ),
    .A2(\design_top.MEM[5][6] ),
    .A3(\design_top.MEM[4][6] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22220_ (.A0(\design_top.MEM[3][6] ),
    .A1(\design_top.MEM[2][6] ),
    .A2(\design_top.MEM[1][6] ),
    .A3(\design_top.MEM[0][6] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22221_ (.A0(_02106_),
    .A1(_02105_),
    .A2(_02104_),
    .A3(_02103_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22222_ (.A0(_02122_),
    .A1(_02117_),
    .A2(_02112_),
    .A3(_02107_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22223_ (.A0(\design_top.MEM[63][5] ),
    .A1(\design_top.MEM[62][5] ),
    .A2(\design_top.MEM[61][5] ),
    .A3(\design_top.MEM[60][5] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22224_ (.A0(\design_top.MEM[59][5] ),
    .A1(\design_top.MEM[58][5] ),
    .A2(\design_top.MEM[57][5] ),
    .A3(\design_top.MEM[56][5] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22225_ (.A0(\design_top.MEM[55][5] ),
    .A1(\design_top.MEM[54][5] ),
    .A2(\design_top.MEM[53][5] ),
    .A3(\design_top.MEM[52][5] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22226_ (.A0(\design_top.MEM[51][5] ),
    .A1(\design_top.MEM[50][5] ),
    .A2(\design_top.MEM[49][5] ),
    .A3(\design_top.MEM[48][5] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22227_ (.A0(_02101_),
    .A1(_02100_),
    .A2(_02099_),
    .A3(_02098_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22228_ (.A0(\design_top.MEM[47][5] ),
    .A1(\design_top.MEM[46][5] ),
    .A2(\design_top.MEM[45][5] ),
    .A3(\design_top.MEM[44][5] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22229_ (.A0(\design_top.MEM[43][5] ),
    .A1(\design_top.MEM[42][5] ),
    .A2(\design_top.MEM[41][5] ),
    .A3(\design_top.MEM[40][5] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22230_ (.A0(\design_top.MEM[39][5] ),
    .A1(\design_top.MEM[38][5] ),
    .A2(\design_top.MEM[37][5] ),
    .A3(\design_top.MEM[36][5] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22231_ (.A0(\design_top.MEM[35][5] ),
    .A1(\design_top.MEM[34][5] ),
    .A2(\design_top.MEM[33][5] ),
    .A3(\design_top.MEM[32][5] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22232_ (.A0(_02096_),
    .A1(_02095_),
    .A2(_02094_),
    .A3(_02093_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22233_ (.A0(\design_top.MEM[31][5] ),
    .A1(\design_top.MEM[30][5] ),
    .A2(\design_top.MEM[29][5] ),
    .A3(\design_top.MEM[28][5] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22234_ (.A0(\design_top.MEM[27][5] ),
    .A1(\design_top.MEM[26][5] ),
    .A2(\design_top.MEM[25][5] ),
    .A3(\design_top.MEM[24][5] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22235_ (.A0(\design_top.MEM[23][5] ),
    .A1(\design_top.MEM[22][5] ),
    .A2(\design_top.MEM[21][5] ),
    .A3(\design_top.MEM[20][5] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22236_ (.A0(\design_top.MEM[19][5] ),
    .A1(\design_top.MEM[18][5] ),
    .A2(\design_top.MEM[17][5] ),
    .A3(\design_top.MEM[16][5] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22237_ (.A0(_02091_),
    .A1(_02090_),
    .A2(_02089_),
    .A3(_02088_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22238_ (.A0(\design_top.MEM[15][5] ),
    .A1(\design_top.MEM[14][5] ),
    .A2(\design_top.MEM[13][5] ),
    .A3(\design_top.MEM[12][5] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22239_ (.A0(\design_top.MEM[11][5] ),
    .A1(\design_top.MEM[10][5] ),
    .A2(\design_top.MEM[9][5] ),
    .A3(\design_top.MEM[8][5] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22240_ (.A0(\design_top.MEM[7][5] ),
    .A1(\design_top.MEM[6][5] ),
    .A2(\design_top.MEM[5][5] ),
    .A3(\design_top.MEM[4][5] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22241_ (.A0(\design_top.MEM[3][5] ),
    .A1(\design_top.MEM[2][5] ),
    .A2(\design_top.MEM[1][5] ),
    .A3(\design_top.MEM[0][5] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22242_ (.A0(_02086_),
    .A1(_02085_),
    .A2(_02084_),
    .A3(_02083_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22243_ (.A0(_02102_),
    .A1(_02097_),
    .A2(_02092_),
    .A3(_02087_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22244_ (.A0(\design_top.MEM[63][4] ),
    .A1(\design_top.MEM[62][4] ),
    .A2(\design_top.MEM[61][4] ),
    .A3(\design_top.MEM[60][4] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22245_ (.A0(\design_top.MEM[59][4] ),
    .A1(\design_top.MEM[58][4] ),
    .A2(\design_top.MEM[57][4] ),
    .A3(\design_top.MEM[56][4] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22246_ (.A0(\design_top.MEM[55][4] ),
    .A1(\design_top.MEM[54][4] ),
    .A2(\design_top.MEM[53][4] ),
    .A3(\design_top.MEM[52][4] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22247_ (.A0(\design_top.MEM[51][4] ),
    .A1(\design_top.MEM[50][4] ),
    .A2(\design_top.MEM[49][4] ),
    .A3(\design_top.MEM[48][4] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22248_ (.A0(_02081_),
    .A1(_02080_),
    .A2(_02079_),
    .A3(_02078_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22249_ (.A0(\design_top.MEM[47][4] ),
    .A1(\design_top.MEM[46][4] ),
    .A2(\design_top.MEM[45][4] ),
    .A3(\design_top.MEM[44][4] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22250_ (.A0(\design_top.MEM[43][4] ),
    .A1(\design_top.MEM[42][4] ),
    .A2(\design_top.MEM[41][4] ),
    .A3(\design_top.MEM[40][4] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22251_ (.A0(\design_top.MEM[39][4] ),
    .A1(\design_top.MEM[38][4] ),
    .A2(\design_top.MEM[37][4] ),
    .A3(\design_top.MEM[36][4] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22252_ (.A0(\design_top.MEM[35][4] ),
    .A1(\design_top.MEM[34][4] ),
    .A2(\design_top.MEM[33][4] ),
    .A3(\design_top.MEM[32][4] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22253_ (.A0(_02076_),
    .A1(_02075_),
    .A2(_02074_),
    .A3(_02073_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22254_ (.A0(\design_top.MEM[31][4] ),
    .A1(\design_top.MEM[30][4] ),
    .A2(\design_top.MEM[29][4] ),
    .A3(\design_top.MEM[28][4] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22255_ (.A0(\design_top.MEM[27][4] ),
    .A1(\design_top.MEM[26][4] ),
    .A2(\design_top.MEM[25][4] ),
    .A3(\design_top.MEM[24][4] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22256_ (.A0(\design_top.MEM[23][4] ),
    .A1(\design_top.MEM[22][4] ),
    .A2(\design_top.MEM[21][4] ),
    .A3(\design_top.MEM[20][4] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22257_ (.A0(\design_top.MEM[19][4] ),
    .A1(\design_top.MEM[18][4] ),
    .A2(\design_top.MEM[17][4] ),
    .A3(\design_top.MEM[16][4] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22258_ (.A0(_02071_),
    .A1(_02070_),
    .A2(_02069_),
    .A3(_02068_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22259_ (.A0(\design_top.MEM[15][4] ),
    .A1(\design_top.MEM[14][4] ),
    .A2(\design_top.MEM[13][4] ),
    .A3(\design_top.MEM[12][4] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22260_ (.A0(\design_top.MEM[11][4] ),
    .A1(\design_top.MEM[10][4] ),
    .A2(\design_top.MEM[9][4] ),
    .A3(\design_top.MEM[8][4] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22261_ (.A0(\design_top.MEM[7][4] ),
    .A1(\design_top.MEM[6][4] ),
    .A2(\design_top.MEM[5][4] ),
    .A3(\design_top.MEM[4][4] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22262_ (.A0(\design_top.MEM[3][4] ),
    .A1(\design_top.MEM[2][4] ),
    .A2(\design_top.MEM[1][4] ),
    .A3(\design_top.MEM[0][4] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22263_ (.A0(_02066_),
    .A1(_02065_),
    .A2(_02064_),
    .A3(_02063_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22264_ (.A0(_02082_),
    .A1(_02077_),
    .A2(_02072_),
    .A3(_02067_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22265_ (.A0(\design_top.MEM[63][3] ),
    .A1(\design_top.MEM[62][3] ),
    .A2(\design_top.MEM[61][3] ),
    .A3(\design_top.MEM[60][3] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22266_ (.A0(\design_top.MEM[59][3] ),
    .A1(\design_top.MEM[58][3] ),
    .A2(\design_top.MEM[57][3] ),
    .A3(\design_top.MEM[56][3] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22267_ (.A0(\design_top.MEM[55][3] ),
    .A1(\design_top.MEM[54][3] ),
    .A2(\design_top.MEM[53][3] ),
    .A3(\design_top.MEM[52][3] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22268_ (.A0(\design_top.MEM[51][3] ),
    .A1(\design_top.MEM[50][3] ),
    .A2(\design_top.MEM[49][3] ),
    .A3(\design_top.MEM[48][3] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22269_ (.A0(_02061_),
    .A1(_02060_),
    .A2(_02059_),
    .A3(_02058_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22270_ (.A0(\design_top.MEM[47][3] ),
    .A1(\design_top.MEM[46][3] ),
    .A2(\design_top.MEM[45][3] ),
    .A3(\design_top.MEM[44][3] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22271_ (.A0(\design_top.MEM[43][3] ),
    .A1(\design_top.MEM[42][3] ),
    .A2(\design_top.MEM[41][3] ),
    .A3(\design_top.MEM[40][3] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22272_ (.A0(\design_top.MEM[39][3] ),
    .A1(\design_top.MEM[38][3] ),
    .A2(\design_top.MEM[37][3] ),
    .A3(\design_top.MEM[36][3] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22273_ (.A0(\design_top.MEM[35][3] ),
    .A1(\design_top.MEM[34][3] ),
    .A2(\design_top.MEM[33][3] ),
    .A3(\design_top.MEM[32][3] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22274_ (.A0(_02056_),
    .A1(_02055_),
    .A2(_02054_),
    .A3(_02053_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22275_ (.A0(\design_top.MEM[31][3] ),
    .A1(\design_top.MEM[30][3] ),
    .A2(\design_top.MEM[29][3] ),
    .A3(\design_top.MEM[28][3] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22276_ (.A0(\design_top.MEM[27][3] ),
    .A1(\design_top.MEM[26][3] ),
    .A2(\design_top.MEM[25][3] ),
    .A3(\design_top.MEM[24][3] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22277_ (.A0(\design_top.MEM[23][3] ),
    .A1(\design_top.MEM[22][3] ),
    .A2(\design_top.MEM[21][3] ),
    .A3(\design_top.MEM[20][3] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22278_ (.A0(\design_top.MEM[19][3] ),
    .A1(\design_top.MEM[18][3] ),
    .A2(\design_top.MEM[17][3] ),
    .A3(\design_top.MEM[16][3] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22279_ (.A0(_02051_),
    .A1(_02050_),
    .A2(_02049_),
    .A3(_02048_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22280_ (.A0(\design_top.MEM[15][3] ),
    .A1(\design_top.MEM[14][3] ),
    .A2(\design_top.MEM[13][3] ),
    .A3(\design_top.MEM[12][3] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22281_ (.A0(\design_top.MEM[11][3] ),
    .A1(\design_top.MEM[10][3] ),
    .A2(\design_top.MEM[9][3] ),
    .A3(\design_top.MEM[8][3] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22282_ (.A0(\design_top.MEM[7][3] ),
    .A1(\design_top.MEM[6][3] ),
    .A2(\design_top.MEM[5][3] ),
    .A3(\design_top.MEM[4][3] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22283_ (.A0(\design_top.MEM[3][3] ),
    .A1(\design_top.MEM[2][3] ),
    .A2(\design_top.MEM[1][3] ),
    .A3(\design_top.MEM[0][3] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22284_ (.A0(_02046_),
    .A1(_02045_),
    .A2(_02044_),
    .A3(_02043_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22285_ (.A0(_02062_),
    .A1(_02057_),
    .A2(_02052_),
    .A3(_02047_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22286_ (.A0(\design_top.MEM[63][2] ),
    .A1(\design_top.MEM[62][2] ),
    .A2(\design_top.MEM[61][2] ),
    .A3(\design_top.MEM[60][2] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22287_ (.A0(\design_top.MEM[59][2] ),
    .A1(\design_top.MEM[58][2] ),
    .A2(\design_top.MEM[57][2] ),
    .A3(\design_top.MEM[56][2] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22288_ (.A0(\design_top.MEM[55][2] ),
    .A1(\design_top.MEM[54][2] ),
    .A2(\design_top.MEM[53][2] ),
    .A3(\design_top.MEM[52][2] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22289_ (.A0(\design_top.MEM[51][2] ),
    .A1(\design_top.MEM[50][2] ),
    .A2(\design_top.MEM[49][2] ),
    .A3(\design_top.MEM[48][2] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22290_ (.A0(_02041_),
    .A1(_02040_),
    .A2(_02039_),
    .A3(_02038_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22291_ (.A0(\design_top.MEM[47][2] ),
    .A1(\design_top.MEM[46][2] ),
    .A2(\design_top.MEM[45][2] ),
    .A3(\design_top.MEM[44][2] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22292_ (.A0(\design_top.MEM[43][2] ),
    .A1(\design_top.MEM[42][2] ),
    .A2(\design_top.MEM[41][2] ),
    .A3(\design_top.MEM[40][2] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22293_ (.A0(\design_top.MEM[39][2] ),
    .A1(\design_top.MEM[38][2] ),
    .A2(\design_top.MEM[37][2] ),
    .A3(\design_top.MEM[36][2] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22294_ (.A0(\design_top.MEM[35][2] ),
    .A1(\design_top.MEM[34][2] ),
    .A2(\design_top.MEM[33][2] ),
    .A3(\design_top.MEM[32][2] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22295_ (.A0(_02036_),
    .A1(_02035_),
    .A2(_02034_),
    .A3(_02033_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22296_ (.A0(\design_top.MEM[31][2] ),
    .A1(\design_top.MEM[30][2] ),
    .A2(\design_top.MEM[29][2] ),
    .A3(\design_top.MEM[28][2] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22297_ (.A0(\design_top.MEM[27][2] ),
    .A1(\design_top.MEM[26][2] ),
    .A2(\design_top.MEM[25][2] ),
    .A3(\design_top.MEM[24][2] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22298_ (.A0(\design_top.MEM[23][2] ),
    .A1(\design_top.MEM[22][2] ),
    .A2(\design_top.MEM[21][2] ),
    .A3(\design_top.MEM[20][2] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22299_ (.A0(\design_top.MEM[19][2] ),
    .A1(\design_top.MEM[18][2] ),
    .A2(\design_top.MEM[17][2] ),
    .A3(\design_top.MEM[16][2] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22300_ (.A0(_02031_),
    .A1(_02030_),
    .A2(_02029_),
    .A3(_02028_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22301_ (.A0(\design_top.MEM[15][2] ),
    .A1(\design_top.MEM[14][2] ),
    .A2(\design_top.MEM[13][2] ),
    .A3(\design_top.MEM[12][2] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22302_ (.A0(\design_top.MEM[11][2] ),
    .A1(\design_top.MEM[10][2] ),
    .A2(\design_top.MEM[9][2] ),
    .A3(\design_top.MEM[8][2] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22303_ (.A0(\design_top.MEM[7][2] ),
    .A1(\design_top.MEM[6][2] ),
    .A2(\design_top.MEM[5][2] ),
    .A3(\design_top.MEM[4][2] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22304_ (.A0(\design_top.MEM[3][2] ),
    .A1(\design_top.MEM[2][2] ),
    .A2(\design_top.MEM[1][2] ),
    .A3(\design_top.MEM[0][2] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22305_ (.A0(_02026_),
    .A1(_02025_),
    .A2(_02024_),
    .A3(_02023_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22306_ (.A0(_02042_),
    .A1(_02037_),
    .A2(_02032_),
    .A3(_02027_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22307_ (.A0(\design_top.MEM[63][1] ),
    .A1(\design_top.MEM[62][1] ),
    .A2(\design_top.MEM[61][1] ),
    .A3(\design_top.MEM[60][1] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22308_ (.A0(\design_top.MEM[59][1] ),
    .A1(\design_top.MEM[58][1] ),
    .A2(\design_top.MEM[57][1] ),
    .A3(\design_top.MEM[56][1] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22309_ (.A0(\design_top.MEM[55][1] ),
    .A1(\design_top.MEM[54][1] ),
    .A2(\design_top.MEM[53][1] ),
    .A3(\design_top.MEM[52][1] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22310_ (.A0(\design_top.MEM[51][1] ),
    .A1(\design_top.MEM[50][1] ),
    .A2(\design_top.MEM[49][1] ),
    .A3(\design_top.MEM[48][1] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22311_ (.A0(_02021_),
    .A1(_02020_),
    .A2(_02019_),
    .A3(_02018_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22312_ (.A0(\design_top.MEM[47][1] ),
    .A1(\design_top.MEM[46][1] ),
    .A2(\design_top.MEM[45][1] ),
    .A3(\design_top.MEM[44][1] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22313_ (.A0(\design_top.MEM[43][1] ),
    .A1(\design_top.MEM[42][1] ),
    .A2(\design_top.MEM[41][1] ),
    .A3(\design_top.MEM[40][1] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22314_ (.A0(\design_top.MEM[39][1] ),
    .A1(\design_top.MEM[38][1] ),
    .A2(\design_top.MEM[37][1] ),
    .A3(\design_top.MEM[36][1] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22315_ (.A0(\design_top.MEM[35][1] ),
    .A1(\design_top.MEM[34][1] ),
    .A2(\design_top.MEM[33][1] ),
    .A3(\design_top.MEM[32][1] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22316_ (.A0(_02016_),
    .A1(_02015_),
    .A2(_02014_),
    .A3(_02013_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22317_ (.A0(\design_top.MEM[31][1] ),
    .A1(\design_top.MEM[30][1] ),
    .A2(\design_top.MEM[29][1] ),
    .A3(\design_top.MEM[28][1] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22318_ (.A0(\design_top.MEM[27][1] ),
    .A1(\design_top.MEM[26][1] ),
    .A2(\design_top.MEM[25][1] ),
    .A3(\design_top.MEM[24][1] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22319_ (.A0(\design_top.MEM[23][1] ),
    .A1(\design_top.MEM[22][1] ),
    .A2(\design_top.MEM[21][1] ),
    .A3(\design_top.MEM[20][1] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22320_ (.A0(\design_top.MEM[19][1] ),
    .A1(\design_top.MEM[18][1] ),
    .A2(\design_top.MEM[17][1] ),
    .A3(\design_top.MEM[16][1] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22321_ (.A0(_02011_),
    .A1(_02010_),
    .A2(_02009_),
    .A3(_02008_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22322_ (.A0(\design_top.MEM[15][1] ),
    .A1(\design_top.MEM[14][1] ),
    .A2(\design_top.MEM[13][1] ),
    .A3(\design_top.MEM[12][1] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22323_ (.A0(\design_top.MEM[11][1] ),
    .A1(\design_top.MEM[10][1] ),
    .A2(\design_top.MEM[9][1] ),
    .A3(\design_top.MEM[8][1] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22324_ (.A0(\design_top.MEM[7][1] ),
    .A1(\design_top.MEM[6][1] ),
    .A2(\design_top.MEM[5][1] ),
    .A3(\design_top.MEM[4][1] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22325_ (.A0(\design_top.MEM[3][1] ),
    .A1(\design_top.MEM[2][1] ),
    .A2(\design_top.MEM[1][1] ),
    .A3(\design_top.MEM[0][1] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22326_ (.A0(_02006_),
    .A1(_02005_),
    .A2(_02004_),
    .A3(_02003_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22327_ (.A0(_02022_),
    .A1(_02017_),
    .A2(_02012_),
    .A3(_02007_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22328_ (.A0(\design_top.MEM[63][0] ),
    .A1(\design_top.MEM[62][0] ),
    .A2(\design_top.MEM[61][0] ),
    .A3(\design_top.MEM[60][0] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22329_ (.A0(\design_top.MEM[59][0] ),
    .A1(\design_top.MEM[58][0] ),
    .A2(\design_top.MEM[57][0] ),
    .A3(\design_top.MEM[56][0] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_02000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22330_ (.A0(\design_top.MEM[55][0] ),
    .A1(\design_top.MEM[54][0] ),
    .A2(\design_top.MEM[53][0] ),
    .A3(\design_top.MEM[52][0] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_01999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22331_ (.A0(\design_top.MEM[51][0] ),
    .A1(\design_top.MEM[50][0] ),
    .A2(\design_top.MEM[49][0] ),
    .A3(\design_top.MEM[48][0] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_01998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22332_ (.A0(_02001_),
    .A1(_02000_),
    .A2(_01999_),
    .A3(_01998_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_02002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22333_ (.A0(\design_top.MEM[47][0] ),
    .A1(\design_top.MEM[46][0] ),
    .A2(\design_top.MEM[45][0] ),
    .A3(\design_top.MEM[44][0] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_01996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22334_ (.A0(\design_top.MEM[43][0] ),
    .A1(\design_top.MEM[42][0] ),
    .A2(\design_top.MEM[41][0] ),
    .A3(\design_top.MEM[40][0] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_01995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22335_ (.A0(\design_top.MEM[39][0] ),
    .A1(\design_top.MEM[38][0] ),
    .A2(\design_top.MEM[37][0] ),
    .A3(\design_top.MEM[36][0] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_01994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22336_ (.A0(\design_top.MEM[35][0] ),
    .A1(\design_top.MEM[34][0] ),
    .A2(\design_top.MEM[33][0] ),
    .A3(\design_top.MEM[32][0] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_01993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22337_ (.A0(_01996_),
    .A1(_01995_),
    .A2(_01994_),
    .A3(_01993_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_01997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22338_ (.A0(\design_top.MEM[31][0] ),
    .A1(\design_top.MEM[30][0] ),
    .A2(\design_top.MEM[29][0] ),
    .A3(\design_top.MEM[28][0] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_01991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22339_ (.A0(\design_top.MEM[27][0] ),
    .A1(\design_top.MEM[26][0] ),
    .A2(\design_top.MEM[25][0] ),
    .A3(\design_top.MEM[24][0] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_01990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22340_ (.A0(\design_top.MEM[23][0] ),
    .A1(\design_top.MEM[22][0] ),
    .A2(\design_top.MEM[21][0] ),
    .A3(\design_top.MEM[20][0] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_01989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22341_ (.A0(\design_top.MEM[19][0] ),
    .A1(\design_top.MEM[18][0] ),
    .A2(\design_top.MEM[17][0] ),
    .A3(\design_top.MEM[16][0] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_01988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22342_ (.A0(_01991_),
    .A1(_01990_),
    .A2(_01989_),
    .A3(_01988_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_01992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22343_ (.A0(\design_top.MEM[15][0] ),
    .A1(\design_top.MEM[14][0] ),
    .A2(\design_top.MEM[13][0] ),
    .A3(\design_top.MEM[12][0] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_01986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22344_ (.A0(\design_top.MEM[11][0] ),
    .A1(\design_top.MEM[10][0] ),
    .A2(\design_top.MEM[9][0] ),
    .A3(\design_top.MEM[8][0] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_01985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22345_ (.A0(\design_top.MEM[7][0] ),
    .A1(\design_top.MEM[6][0] ),
    .A2(\design_top.MEM[5][0] ),
    .A3(\design_top.MEM[4][0] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_01984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22346_ (.A0(\design_top.MEM[3][0] ),
    .A1(\design_top.MEM[2][0] ),
    .A2(\design_top.MEM[1][0] ),
    .A3(\design_top.MEM[0][0] ),
    .S0(_02651_),
    .S1(_02660_),
    .X(_01983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22347_ (.A0(_01986_),
    .A1(_01985_),
    .A2(_01984_),
    .A3(_01983_),
    .S0(_02859_),
    .S1(_02860_),
    .X(_01987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22348_ (.A0(_02002_),
    .A1(_01997_),
    .A2(_01992_),
    .A3(_01987_),
    .S0(_02861_),
    .S1(_02862_),
    .X(_00109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22349_ (.A0(\design_top.MEM[0][31] ),
    .A1(\design_top.MEM[1][31] ),
    .A2(\design_top.MEM[2][31] ),
    .A3(\design_top.MEM[3][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22350_ (.A0(\design_top.MEM[4][31] ),
    .A1(\design_top.MEM[5][31] ),
    .A2(\design_top.MEM[6][31] ),
    .A3(\design_top.MEM[7][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22351_ (.A0(\design_top.MEM[8][31] ),
    .A1(\design_top.MEM[9][31] ),
    .A2(\design_top.MEM[10][31] ),
    .A3(\design_top.MEM[11][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22352_ (.A0(\design_top.MEM[12][31] ),
    .A1(\design_top.MEM[13][31] ),
    .A2(\design_top.MEM[14][31] ),
    .A3(\design_top.MEM[15][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22353_ (.A0(_03894_),
    .A1(_03895_),
    .A2(_03896_),
    .A3(_03897_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22354_ (.A0(\design_top.MEM[16][31] ),
    .A1(\design_top.MEM[17][31] ),
    .A2(\design_top.MEM[18][31] ),
    .A3(\design_top.MEM[19][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22355_ (.A0(\design_top.MEM[20][31] ),
    .A1(\design_top.MEM[21][31] ),
    .A2(\design_top.MEM[22][31] ),
    .A3(\design_top.MEM[23][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22356_ (.A0(\design_top.MEM[24][31] ),
    .A1(\design_top.MEM[25][31] ),
    .A2(\design_top.MEM[26][31] ),
    .A3(\design_top.MEM[27][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22357_ (.A0(\design_top.MEM[28][31] ),
    .A1(\design_top.MEM[29][31] ),
    .A2(\design_top.MEM[30][31] ),
    .A3(\design_top.MEM[31][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22358_ (.A0(_03899_),
    .A1(_03900_),
    .A2(_03901_),
    .A3(_03902_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22359_ (.A0(\design_top.MEM[32][31] ),
    .A1(\design_top.MEM[33][31] ),
    .A2(\design_top.MEM[34][31] ),
    .A3(\design_top.MEM[35][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22360_ (.A0(\design_top.MEM[36][31] ),
    .A1(\design_top.MEM[37][31] ),
    .A2(\design_top.MEM[38][31] ),
    .A3(\design_top.MEM[39][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22361_ (.A0(\design_top.MEM[40][31] ),
    .A1(\design_top.MEM[41][31] ),
    .A2(\design_top.MEM[42][31] ),
    .A3(\design_top.MEM[43][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22362_ (.A0(\design_top.MEM[44][31] ),
    .A1(\design_top.MEM[45][31] ),
    .A2(\design_top.MEM[46][31] ),
    .A3(\design_top.MEM[47][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22363_ (.A0(_03904_),
    .A1(_03905_),
    .A2(_03906_),
    .A3(_03907_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22364_ (.A0(\design_top.MEM[48][31] ),
    .A1(\design_top.MEM[49][31] ),
    .A2(\design_top.MEM[50][31] ),
    .A3(\design_top.MEM[51][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22365_ (.A0(\design_top.MEM[52][31] ),
    .A1(\design_top.MEM[53][31] ),
    .A2(\design_top.MEM[54][31] ),
    .A3(\design_top.MEM[55][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22366_ (.A0(\design_top.MEM[56][31] ),
    .A1(\design_top.MEM[57][31] ),
    .A2(\design_top.MEM[58][31] ),
    .A3(\design_top.MEM[59][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22367_ (.A0(\design_top.MEM[60][31] ),
    .A1(\design_top.MEM[61][31] ),
    .A2(\design_top.MEM[62][31] ),
    .A3(\design_top.MEM[63][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22368_ (.A0(_03909_),
    .A1(_03910_),
    .A2(_03911_),
    .A3(_03912_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22369_ (.A0(_03898_),
    .A1(_03903_),
    .A2(_03908_),
    .A3(_03913_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22370_ (.A0(\design_top.MEM[0][30] ),
    .A1(\design_top.MEM[1][30] ),
    .A2(\design_top.MEM[2][30] ),
    .A3(\design_top.MEM[3][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22371_ (.A0(\design_top.MEM[4][30] ),
    .A1(\design_top.MEM[5][30] ),
    .A2(\design_top.MEM[6][30] ),
    .A3(\design_top.MEM[7][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22372_ (.A0(\design_top.MEM[8][30] ),
    .A1(\design_top.MEM[9][30] ),
    .A2(\design_top.MEM[10][30] ),
    .A3(\design_top.MEM[11][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22373_ (.A0(\design_top.MEM[12][30] ),
    .A1(\design_top.MEM[13][30] ),
    .A2(\design_top.MEM[14][30] ),
    .A3(\design_top.MEM[15][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22374_ (.A0(_03874_),
    .A1(_03875_),
    .A2(_03876_),
    .A3(_03877_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22375_ (.A0(\design_top.MEM[16][30] ),
    .A1(\design_top.MEM[17][30] ),
    .A2(\design_top.MEM[18][30] ),
    .A3(\design_top.MEM[19][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22376_ (.A0(\design_top.MEM[20][30] ),
    .A1(\design_top.MEM[21][30] ),
    .A2(\design_top.MEM[22][30] ),
    .A3(\design_top.MEM[23][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22377_ (.A0(\design_top.MEM[24][30] ),
    .A1(\design_top.MEM[25][30] ),
    .A2(\design_top.MEM[26][30] ),
    .A3(\design_top.MEM[27][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22378_ (.A0(\design_top.MEM[28][30] ),
    .A1(\design_top.MEM[29][30] ),
    .A2(\design_top.MEM[30][30] ),
    .A3(\design_top.MEM[31][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22379_ (.A0(_03879_),
    .A1(_03880_),
    .A2(_03881_),
    .A3(_03882_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22380_ (.A0(\design_top.MEM[32][30] ),
    .A1(\design_top.MEM[33][30] ),
    .A2(\design_top.MEM[34][30] ),
    .A3(\design_top.MEM[35][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22381_ (.A0(\design_top.MEM[36][30] ),
    .A1(\design_top.MEM[37][30] ),
    .A2(\design_top.MEM[38][30] ),
    .A3(\design_top.MEM[39][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22382_ (.A0(\design_top.MEM[40][30] ),
    .A1(\design_top.MEM[41][30] ),
    .A2(\design_top.MEM[42][30] ),
    .A3(\design_top.MEM[43][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22383_ (.A0(\design_top.MEM[44][30] ),
    .A1(\design_top.MEM[45][30] ),
    .A2(\design_top.MEM[46][30] ),
    .A3(\design_top.MEM[47][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22384_ (.A0(_03884_),
    .A1(_03885_),
    .A2(_03886_),
    .A3(_03887_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22385_ (.A0(\design_top.MEM[48][30] ),
    .A1(\design_top.MEM[49][30] ),
    .A2(\design_top.MEM[50][30] ),
    .A3(\design_top.MEM[51][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22386_ (.A0(\design_top.MEM[52][30] ),
    .A1(\design_top.MEM[53][30] ),
    .A2(\design_top.MEM[54][30] ),
    .A3(\design_top.MEM[55][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22387_ (.A0(\design_top.MEM[56][30] ),
    .A1(\design_top.MEM[57][30] ),
    .A2(\design_top.MEM[58][30] ),
    .A3(\design_top.MEM[59][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22388_ (.A0(\design_top.MEM[60][30] ),
    .A1(\design_top.MEM[61][30] ),
    .A2(\design_top.MEM[62][30] ),
    .A3(\design_top.MEM[63][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22389_ (.A0(_03889_),
    .A1(_03890_),
    .A2(_03891_),
    .A3(_03892_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22390_ (.A0(_03878_),
    .A1(_03883_),
    .A2(_03888_),
    .A3(_03893_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22391_ (.A0(\design_top.MEM[0][29] ),
    .A1(\design_top.MEM[1][29] ),
    .A2(\design_top.MEM[2][29] ),
    .A3(\design_top.MEM[3][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22392_ (.A0(\design_top.MEM[4][29] ),
    .A1(\design_top.MEM[5][29] ),
    .A2(\design_top.MEM[6][29] ),
    .A3(\design_top.MEM[7][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22393_ (.A0(\design_top.MEM[8][29] ),
    .A1(\design_top.MEM[9][29] ),
    .A2(\design_top.MEM[10][29] ),
    .A3(\design_top.MEM[11][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22394_ (.A0(\design_top.MEM[12][29] ),
    .A1(\design_top.MEM[13][29] ),
    .A2(\design_top.MEM[14][29] ),
    .A3(\design_top.MEM[15][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22395_ (.A0(_03854_),
    .A1(_03855_),
    .A2(_03856_),
    .A3(_03857_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22396_ (.A0(\design_top.MEM[16][29] ),
    .A1(\design_top.MEM[17][29] ),
    .A2(\design_top.MEM[18][29] ),
    .A3(\design_top.MEM[19][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22397_ (.A0(\design_top.MEM[20][29] ),
    .A1(\design_top.MEM[21][29] ),
    .A2(\design_top.MEM[22][29] ),
    .A3(\design_top.MEM[23][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22398_ (.A0(\design_top.MEM[24][29] ),
    .A1(\design_top.MEM[25][29] ),
    .A2(\design_top.MEM[26][29] ),
    .A3(\design_top.MEM[27][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22399_ (.A0(\design_top.MEM[28][29] ),
    .A1(\design_top.MEM[29][29] ),
    .A2(\design_top.MEM[30][29] ),
    .A3(\design_top.MEM[31][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22400_ (.A0(_03859_),
    .A1(_03860_),
    .A2(_03861_),
    .A3(_03862_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22401_ (.A0(\design_top.MEM[32][29] ),
    .A1(\design_top.MEM[33][29] ),
    .A2(\design_top.MEM[34][29] ),
    .A3(\design_top.MEM[35][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22402_ (.A0(\design_top.MEM[36][29] ),
    .A1(\design_top.MEM[37][29] ),
    .A2(\design_top.MEM[38][29] ),
    .A3(\design_top.MEM[39][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22403_ (.A0(\design_top.MEM[40][29] ),
    .A1(\design_top.MEM[41][29] ),
    .A2(\design_top.MEM[42][29] ),
    .A3(\design_top.MEM[43][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22404_ (.A0(\design_top.MEM[44][29] ),
    .A1(\design_top.MEM[45][29] ),
    .A2(\design_top.MEM[46][29] ),
    .A3(\design_top.MEM[47][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22405_ (.A0(_03864_),
    .A1(_03865_),
    .A2(_03866_),
    .A3(_03867_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22406_ (.A0(\design_top.MEM[48][29] ),
    .A1(\design_top.MEM[49][29] ),
    .A2(\design_top.MEM[50][29] ),
    .A3(\design_top.MEM[51][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22407_ (.A0(\design_top.MEM[52][29] ),
    .A1(\design_top.MEM[53][29] ),
    .A2(\design_top.MEM[54][29] ),
    .A3(\design_top.MEM[55][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22408_ (.A0(\design_top.MEM[56][29] ),
    .A1(\design_top.MEM[57][29] ),
    .A2(\design_top.MEM[58][29] ),
    .A3(\design_top.MEM[59][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22409_ (.A0(\design_top.MEM[60][29] ),
    .A1(\design_top.MEM[61][29] ),
    .A2(\design_top.MEM[62][29] ),
    .A3(\design_top.MEM[63][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22410_ (.A0(_03869_),
    .A1(_03870_),
    .A2(_03871_),
    .A3(_03872_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22411_ (.A0(_03858_),
    .A1(_03863_),
    .A2(_03868_),
    .A3(_03873_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22412_ (.A0(\design_top.MEM[0][28] ),
    .A1(\design_top.MEM[1][28] ),
    .A2(\design_top.MEM[2][28] ),
    .A3(\design_top.MEM[3][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22413_ (.A0(\design_top.MEM[4][28] ),
    .A1(\design_top.MEM[5][28] ),
    .A2(\design_top.MEM[6][28] ),
    .A3(\design_top.MEM[7][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22414_ (.A0(\design_top.MEM[8][28] ),
    .A1(\design_top.MEM[9][28] ),
    .A2(\design_top.MEM[10][28] ),
    .A3(\design_top.MEM[11][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22415_ (.A0(\design_top.MEM[12][28] ),
    .A1(\design_top.MEM[13][28] ),
    .A2(\design_top.MEM[14][28] ),
    .A3(\design_top.MEM[15][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22416_ (.A0(_03834_),
    .A1(_03835_),
    .A2(_03836_),
    .A3(_03837_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22417_ (.A0(\design_top.MEM[16][28] ),
    .A1(\design_top.MEM[17][28] ),
    .A2(\design_top.MEM[18][28] ),
    .A3(\design_top.MEM[19][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22418_ (.A0(\design_top.MEM[20][28] ),
    .A1(\design_top.MEM[21][28] ),
    .A2(\design_top.MEM[22][28] ),
    .A3(\design_top.MEM[23][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22419_ (.A0(\design_top.MEM[24][28] ),
    .A1(\design_top.MEM[25][28] ),
    .A2(\design_top.MEM[26][28] ),
    .A3(\design_top.MEM[27][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22420_ (.A0(\design_top.MEM[28][28] ),
    .A1(\design_top.MEM[29][28] ),
    .A2(\design_top.MEM[30][28] ),
    .A3(\design_top.MEM[31][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22421_ (.A0(_03839_),
    .A1(_03840_),
    .A2(_03841_),
    .A3(_03842_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22422_ (.A0(\design_top.MEM[32][28] ),
    .A1(\design_top.MEM[33][28] ),
    .A2(\design_top.MEM[34][28] ),
    .A3(\design_top.MEM[35][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22423_ (.A0(\design_top.MEM[36][28] ),
    .A1(\design_top.MEM[37][28] ),
    .A2(\design_top.MEM[38][28] ),
    .A3(\design_top.MEM[39][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22424_ (.A0(\design_top.MEM[40][28] ),
    .A1(\design_top.MEM[41][28] ),
    .A2(\design_top.MEM[42][28] ),
    .A3(\design_top.MEM[43][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22425_ (.A0(\design_top.MEM[44][28] ),
    .A1(\design_top.MEM[45][28] ),
    .A2(\design_top.MEM[46][28] ),
    .A3(\design_top.MEM[47][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22426_ (.A0(_03844_),
    .A1(_03845_),
    .A2(_03846_),
    .A3(_03847_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22427_ (.A0(\design_top.MEM[48][28] ),
    .A1(\design_top.MEM[49][28] ),
    .A2(\design_top.MEM[50][28] ),
    .A3(\design_top.MEM[51][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22428_ (.A0(\design_top.MEM[52][28] ),
    .A1(\design_top.MEM[53][28] ),
    .A2(\design_top.MEM[54][28] ),
    .A3(\design_top.MEM[55][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22429_ (.A0(\design_top.MEM[56][28] ),
    .A1(\design_top.MEM[57][28] ),
    .A2(\design_top.MEM[58][28] ),
    .A3(\design_top.MEM[59][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22430_ (.A0(\design_top.MEM[60][28] ),
    .A1(\design_top.MEM[61][28] ),
    .A2(\design_top.MEM[62][28] ),
    .A3(\design_top.MEM[63][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22431_ (.A0(_03849_),
    .A1(_03850_),
    .A2(_03851_),
    .A3(_03852_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22432_ (.A0(_03838_),
    .A1(_03843_),
    .A2(_03848_),
    .A3(_03853_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22433_ (.A0(\design_top.MEM[0][27] ),
    .A1(\design_top.MEM[1][27] ),
    .A2(\design_top.MEM[2][27] ),
    .A3(\design_top.MEM[3][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22434_ (.A0(\design_top.MEM[4][27] ),
    .A1(\design_top.MEM[5][27] ),
    .A2(\design_top.MEM[6][27] ),
    .A3(\design_top.MEM[7][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22435_ (.A0(\design_top.MEM[8][27] ),
    .A1(\design_top.MEM[9][27] ),
    .A2(\design_top.MEM[10][27] ),
    .A3(\design_top.MEM[11][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22436_ (.A0(\design_top.MEM[12][27] ),
    .A1(\design_top.MEM[13][27] ),
    .A2(\design_top.MEM[14][27] ),
    .A3(\design_top.MEM[15][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22437_ (.A0(_03814_),
    .A1(_03815_),
    .A2(_03816_),
    .A3(_03817_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22438_ (.A0(\design_top.MEM[16][27] ),
    .A1(\design_top.MEM[17][27] ),
    .A2(\design_top.MEM[18][27] ),
    .A3(\design_top.MEM[19][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22439_ (.A0(\design_top.MEM[20][27] ),
    .A1(\design_top.MEM[21][27] ),
    .A2(\design_top.MEM[22][27] ),
    .A3(\design_top.MEM[23][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22440_ (.A0(\design_top.MEM[24][27] ),
    .A1(\design_top.MEM[25][27] ),
    .A2(\design_top.MEM[26][27] ),
    .A3(\design_top.MEM[27][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22441_ (.A0(\design_top.MEM[28][27] ),
    .A1(\design_top.MEM[29][27] ),
    .A2(\design_top.MEM[30][27] ),
    .A3(\design_top.MEM[31][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22442_ (.A0(_03819_),
    .A1(_03820_),
    .A2(_03821_),
    .A3(_03822_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22443_ (.A0(\design_top.MEM[32][27] ),
    .A1(\design_top.MEM[33][27] ),
    .A2(\design_top.MEM[34][27] ),
    .A3(\design_top.MEM[35][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22444_ (.A0(\design_top.MEM[36][27] ),
    .A1(\design_top.MEM[37][27] ),
    .A2(\design_top.MEM[38][27] ),
    .A3(\design_top.MEM[39][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22445_ (.A0(\design_top.MEM[40][27] ),
    .A1(\design_top.MEM[41][27] ),
    .A2(\design_top.MEM[42][27] ),
    .A3(\design_top.MEM[43][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22446_ (.A0(\design_top.MEM[44][27] ),
    .A1(\design_top.MEM[45][27] ),
    .A2(\design_top.MEM[46][27] ),
    .A3(\design_top.MEM[47][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22447_ (.A0(_03824_),
    .A1(_03825_),
    .A2(_03826_),
    .A3(_03827_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22448_ (.A0(\design_top.MEM[48][27] ),
    .A1(\design_top.MEM[49][27] ),
    .A2(\design_top.MEM[50][27] ),
    .A3(\design_top.MEM[51][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22449_ (.A0(\design_top.MEM[52][27] ),
    .A1(\design_top.MEM[53][27] ),
    .A2(\design_top.MEM[54][27] ),
    .A3(\design_top.MEM[55][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22450_ (.A0(\design_top.MEM[56][27] ),
    .A1(\design_top.MEM[57][27] ),
    .A2(\design_top.MEM[58][27] ),
    .A3(\design_top.MEM[59][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22451_ (.A0(\design_top.MEM[60][27] ),
    .A1(\design_top.MEM[61][27] ),
    .A2(\design_top.MEM[62][27] ),
    .A3(\design_top.MEM[63][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22452_ (.A0(_03829_),
    .A1(_03830_),
    .A2(_03831_),
    .A3(_03832_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22453_ (.A0(_03818_),
    .A1(_03823_),
    .A2(_03828_),
    .A3(_03833_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22454_ (.A0(\design_top.MEM[0][26] ),
    .A1(\design_top.MEM[1][26] ),
    .A2(\design_top.MEM[2][26] ),
    .A3(\design_top.MEM[3][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22455_ (.A0(\design_top.MEM[4][26] ),
    .A1(\design_top.MEM[5][26] ),
    .A2(\design_top.MEM[6][26] ),
    .A3(\design_top.MEM[7][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22456_ (.A0(\design_top.MEM[8][26] ),
    .A1(\design_top.MEM[9][26] ),
    .A2(\design_top.MEM[10][26] ),
    .A3(\design_top.MEM[11][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22457_ (.A0(\design_top.MEM[12][26] ),
    .A1(\design_top.MEM[13][26] ),
    .A2(\design_top.MEM[14][26] ),
    .A3(\design_top.MEM[15][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22458_ (.A0(_03794_),
    .A1(_03795_),
    .A2(_03796_),
    .A3(_03797_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22459_ (.A0(\design_top.MEM[16][26] ),
    .A1(\design_top.MEM[17][26] ),
    .A2(\design_top.MEM[18][26] ),
    .A3(\design_top.MEM[19][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22460_ (.A0(\design_top.MEM[20][26] ),
    .A1(\design_top.MEM[21][26] ),
    .A2(\design_top.MEM[22][26] ),
    .A3(\design_top.MEM[23][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22461_ (.A0(\design_top.MEM[24][26] ),
    .A1(\design_top.MEM[25][26] ),
    .A2(\design_top.MEM[26][26] ),
    .A3(\design_top.MEM[27][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22462_ (.A0(\design_top.MEM[28][26] ),
    .A1(\design_top.MEM[29][26] ),
    .A2(\design_top.MEM[30][26] ),
    .A3(\design_top.MEM[31][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22463_ (.A0(_03799_),
    .A1(_03800_),
    .A2(_03801_),
    .A3(_03802_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22464_ (.A0(\design_top.MEM[32][26] ),
    .A1(\design_top.MEM[33][26] ),
    .A2(\design_top.MEM[34][26] ),
    .A3(\design_top.MEM[35][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22465_ (.A0(\design_top.MEM[36][26] ),
    .A1(\design_top.MEM[37][26] ),
    .A2(\design_top.MEM[38][26] ),
    .A3(\design_top.MEM[39][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22466_ (.A0(\design_top.MEM[40][26] ),
    .A1(\design_top.MEM[41][26] ),
    .A2(\design_top.MEM[42][26] ),
    .A3(\design_top.MEM[43][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22467_ (.A0(\design_top.MEM[44][26] ),
    .A1(\design_top.MEM[45][26] ),
    .A2(\design_top.MEM[46][26] ),
    .A3(\design_top.MEM[47][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22468_ (.A0(_03804_),
    .A1(_03805_),
    .A2(_03806_),
    .A3(_03807_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22469_ (.A0(\design_top.MEM[48][26] ),
    .A1(\design_top.MEM[49][26] ),
    .A2(\design_top.MEM[50][26] ),
    .A3(\design_top.MEM[51][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22470_ (.A0(\design_top.MEM[52][26] ),
    .A1(\design_top.MEM[53][26] ),
    .A2(\design_top.MEM[54][26] ),
    .A3(\design_top.MEM[55][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22471_ (.A0(\design_top.MEM[56][26] ),
    .A1(\design_top.MEM[57][26] ),
    .A2(\design_top.MEM[58][26] ),
    .A3(\design_top.MEM[59][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22472_ (.A0(\design_top.MEM[60][26] ),
    .A1(\design_top.MEM[61][26] ),
    .A2(\design_top.MEM[62][26] ),
    .A3(\design_top.MEM[63][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22473_ (.A0(_03809_),
    .A1(_03810_),
    .A2(_03811_),
    .A3(_03812_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22474_ (.A0(_03798_),
    .A1(_03803_),
    .A2(_03808_),
    .A3(_03813_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22475_ (.A0(\design_top.MEM[0][25] ),
    .A1(\design_top.MEM[1][25] ),
    .A2(\design_top.MEM[2][25] ),
    .A3(\design_top.MEM[3][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22476_ (.A0(\design_top.MEM[4][25] ),
    .A1(\design_top.MEM[5][25] ),
    .A2(\design_top.MEM[6][25] ),
    .A3(\design_top.MEM[7][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22477_ (.A0(\design_top.MEM[8][25] ),
    .A1(\design_top.MEM[9][25] ),
    .A2(\design_top.MEM[10][25] ),
    .A3(\design_top.MEM[11][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22478_ (.A0(\design_top.MEM[12][25] ),
    .A1(\design_top.MEM[13][25] ),
    .A2(\design_top.MEM[14][25] ),
    .A3(\design_top.MEM[15][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22479_ (.A0(_03774_),
    .A1(_03775_),
    .A2(_03776_),
    .A3(_03777_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22480_ (.A0(\design_top.MEM[16][25] ),
    .A1(\design_top.MEM[17][25] ),
    .A2(\design_top.MEM[18][25] ),
    .A3(\design_top.MEM[19][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22481_ (.A0(\design_top.MEM[20][25] ),
    .A1(\design_top.MEM[21][25] ),
    .A2(\design_top.MEM[22][25] ),
    .A3(\design_top.MEM[23][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22482_ (.A0(\design_top.MEM[24][25] ),
    .A1(\design_top.MEM[25][25] ),
    .A2(\design_top.MEM[26][25] ),
    .A3(\design_top.MEM[27][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22483_ (.A0(\design_top.MEM[28][25] ),
    .A1(\design_top.MEM[29][25] ),
    .A2(\design_top.MEM[30][25] ),
    .A3(\design_top.MEM[31][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22484_ (.A0(_03779_),
    .A1(_03780_),
    .A2(_03781_),
    .A3(_03782_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22485_ (.A0(\design_top.MEM[32][25] ),
    .A1(\design_top.MEM[33][25] ),
    .A2(\design_top.MEM[34][25] ),
    .A3(\design_top.MEM[35][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22486_ (.A0(\design_top.MEM[36][25] ),
    .A1(\design_top.MEM[37][25] ),
    .A2(\design_top.MEM[38][25] ),
    .A3(\design_top.MEM[39][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22487_ (.A0(\design_top.MEM[40][25] ),
    .A1(\design_top.MEM[41][25] ),
    .A2(\design_top.MEM[42][25] ),
    .A3(\design_top.MEM[43][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22488_ (.A0(\design_top.MEM[44][25] ),
    .A1(\design_top.MEM[45][25] ),
    .A2(\design_top.MEM[46][25] ),
    .A3(\design_top.MEM[47][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22489_ (.A0(_03784_),
    .A1(_03785_),
    .A2(_03786_),
    .A3(_03787_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22490_ (.A0(\design_top.MEM[48][25] ),
    .A1(\design_top.MEM[49][25] ),
    .A2(\design_top.MEM[50][25] ),
    .A3(\design_top.MEM[51][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22491_ (.A0(\design_top.MEM[52][25] ),
    .A1(\design_top.MEM[53][25] ),
    .A2(\design_top.MEM[54][25] ),
    .A3(\design_top.MEM[55][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22492_ (.A0(\design_top.MEM[56][25] ),
    .A1(\design_top.MEM[57][25] ),
    .A2(\design_top.MEM[58][25] ),
    .A3(\design_top.MEM[59][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22493_ (.A0(\design_top.MEM[60][25] ),
    .A1(\design_top.MEM[61][25] ),
    .A2(\design_top.MEM[62][25] ),
    .A3(\design_top.MEM[63][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22494_ (.A0(_03789_),
    .A1(_03790_),
    .A2(_03791_),
    .A3(_03792_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22495_ (.A0(_03778_),
    .A1(_03783_),
    .A2(_03788_),
    .A3(_03793_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22496_ (.A0(\design_top.MEM[0][24] ),
    .A1(\design_top.MEM[1][24] ),
    .A2(\design_top.MEM[2][24] ),
    .A3(\design_top.MEM[3][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22497_ (.A0(\design_top.MEM[4][24] ),
    .A1(\design_top.MEM[5][24] ),
    .A2(\design_top.MEM[6][24] ),
    .A3(\design_top.MEM[7][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22498_ (.A0(\design_top.MEM[8][24] ),
    .A1(\design_top.MEM[9][24] ),
    .A2(\design_top.MEM[10][24] ),
    .A3(\design_top.MEM[11][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22499_ (.A0(\design_top.MEM[12][24] ),
    .A1(\design_top.MEM[13][24] ),
    .A2(\design_top.MEM[14][24] ),
    .A3(\design_top.MEM[15][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22500_ (.A0(_03754_),
    .A1(_03755_),
    .A2(_03756_),
    .A3(_03757_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22501_ (.A0(\design_top.MEM[16][24] ),
    .A1(\design_top.MEM[17][24] ),
    .A2(\design_top.MEM[18][24] ),
    .A3(\design_top.MEM[19][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22502_ (.A0(\design_top.MEM[20][24] ),
    .A1(\design_top.MEM[21][24] ),
    .A2(\design_top.MEM[22][24] ),
    .A3(\design_top.MEM[23][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22503_ (.A0(\design_top.MEM[24][24] ),
    .A1(\design_top.MEM[25][24] ),
    .A2(\design_top.MEM[26][24] ),
    .A3(\design_top.MEM[27][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22504_ (.A0(\design_top.MEM[28][24] ),
    .A1(\design_top.MEM[29][24] ),
    .A2(\design_top.MEM[30][24] ),
    .A3(\design_top.MEM[31][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22505_ (.A0(_03759_),
    .A1(_03760_),
    .A2(_03761_),
    .A3(_03762_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22506_ (.A0(\design_top.MEM[32][24] ),
    .A1(\design_top.MEM[33][24] ),
    .A2(\design_top.MEM[34][24] ),
    .A3(\design_top.MEM[35][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22507_ (.A0(\design_top.MEM[36][24] ),
    .A1(\design_top.MEM[37][24] ),
    .A2(\design_top.MEM[38][24] ),
    .A3(\design_top.MEM[39][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22508_ (.A0(\design_top.MEM[40][24] ),
    .A1(\design_top.MEM[41][24] ),
    .A2(\design_top.MEM[42][24] ),
    .A3(\design_top.MEM[43][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22509_ (.A0(\design_top.MEM[44][24] ),
    .A1(\design_top.MEM[45][24] ),
    .A2(\design_top.MEM[46][24] ),
    .A3(\design_top.MEM[47][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22510_ (.A0(_03764_),
    .A1(_03765_),
    .A2(_03766_),
    .A3(_03767_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22511_ (.A0(\design_top.MEM[48][24] ),
    .A1(\design_top.MEM[49][24] ),
    .A2(\design_top.MEM[50][24] ),
    .A3(\design_top.MEM[51][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22512_ (.A0(\design_top.MEM[52][24] ),
    .A1(\design_top.MEM[53][24] ),
    .A2(\design_top.MEM[54][24] ),
    .A3(\design_top.MEM[55][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22513_ (.A0(\design_top.MEM[56][24] ),
    .A1(\design_top.MEM[57][24] ),
    .A2(\design_top.MEM[58][24] ),
    .A3(\design_top.MEM[59][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22514_ (.A0(\design_top.MEM[60][24] ),
    .A1(\design_top.MEM[61][24] ),
    .A2(\design_top.MEM[62][24] ),
    .A3(\design_top.MEM[63][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22515_ (.A0(_03769_),
    .A1(_03770_),
    .A2(_03771_),
    .A3(_03772_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22516_ (.A0(_03758_),
    .A1(_03763_),
    .A2(_03768_),
    .A3(_03773_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22517_ (.A0(\design_top.MEM[0][23] ),
    .A1(\design_top.MEM[1][23] ),
    .A2(\design_top.MEM[2][23] ),
    .A3(\design_top.MEM[3][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22518_ (.A0(\design_top.MEM[4][23] ),
    .A1(\design_top.MEM[5][23] ),
    .A2(\design_top.MEM[6][23] ),
    .A3(\design_top.MEM[7][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22519_ (.A0(\design_top.MEM[8][23] ),
    .A1(\design_top.MEM[9][23] ),
    .A2(\design_top.MEM[10][23] ),
    .A3(\design_top.MEM[11][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22520_ (.A0(\design_top.MEM[12][23] ),
    .A1(\design_top.MEM[13][23] ),
    .A2(\design_top.MEM[14][23] ),
    .A3(\design_top.MEM[15][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22521_ (.A0(_03734_),
    .A1(_03735_),
    .A2(_03736_),
    .A3(_03737_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22522_ (.A0(\design_top.MEM[16][23] ),
    .A1(\design_top.MEM[17][23] ),
    .A2(\design_top.MEM[18][23] ),
    .A3(\design_top.MEM[19][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22523_ (.A0(\design_top.MEM[20][23] ),
    .A1(\design_top.MEM[21][23] ),
    .A2(\design_top.MEM[22][23] ),
    .A3(\design_top.MEM[23][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22524_ (.A0(\design_top.MEM[24][23] ),
    .A1(\design_top.MEM[25][23] ),
    .A2(\design_top.MEM[26][23] ),
    .A3(\design_top.MEM[27][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22525_ (.A0(\design_top.MEM[28][23] ),
    .A1(\design_top.MEM[29][23] ),
    .A2(\design_top.MEM[30][23] ),
    .A3(\design_top.MEM[31][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22526_ (.A0(_03739_),
    .A1(_03740_),
    .A2(_03741_),
    .A3(_03742_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22527_ (.A0(\design_top.MEM[32][23] ),
    .A1(\design_top.MEM[33][23] ),
    .A2(\design_top.MEM[34][23] ),
    .A3(\design_top.MEM[35][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22528_ (.A0(\design_top.MEM[36][23] ),
    .A1(\design_top.MEM[37][23] ),
    .A2(\design_top.MEM[38][23] ),
    .A3(\design_top.MEM[39][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22529_ (.A0(\design_top.MEM[40][23] ),
    .A1(\design_top.MEM[41][23] ),
    .A2(\design_top.MEM[42][23] ),
    .A3(\design_top.MEM[43][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22530_ (.A0(\design_top.MEM[44][23] ),
    .A1(\design_top.MEM[45][23] ),
    .A2(\design_top.MEM[46][23] ),
    .A3(\design_top.MEM[47][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22531_ (.A0(_03744_),
    .A1(_03745_),
    .A2(_03746_),
    .A3(_03747_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22532_ (.A0(\design_top.MEM[48][23] ),
    .A1(\design_top.MEM[49][23] ),
    .A2(\design_top.MEM[50][23] ),
    .A3(\design_top.MEM[51][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22533_ (.A0(\design_top.MEM[52][23] ),
    .A1(\design_top.MEM[53][23] ),
    .A2(\design_top.MEM[54][23] ),
    .A3(\design_top.MEM[55][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22534_ (.A0(\design_top.MEM[56][23] ),
    .A1(\design_top.MEM[57][23] ),
    .A2(\design_top.MEM[58][23] ),
    .A3(\design_top.MEM[59][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22535_ (.A0(\design_top.MEM[60][23] ),
    .A1(\design_top.MEM[61][23] ),
    .A2(\design_top.MEM[62][23] ),
    .A3(\design_top.MEM[63][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22536_ (.A0(_03749_),
    .A1(_03750_),
    .A2(_03751_),
    .A3(_03752_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22537_ (.A0(_03738_),
    .A1(_03743_),
    .A2(_03748_),
    .A3(_03753_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22538_ (.A0(\design_top.MEM[0][22] ),
    .A1(\design_top.MEM[1][22] ),
    .A2(\design_top.MEM[2][22] ),
    .A3(\design_top.MEM[3][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22539_ (.A0(\design_top.MEM[4][22] ),
    .A1(\design_top.MEM[5][22] ),
    .A2(\design_top.MEM[6][22] ),
    .A3(\design_top.MEM[7][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22540_ (.A0(\design_top.MEM[8][22] ),
    .A1(\design_top.MEM[9][22] ),
    .A2(\design_top.MEM[10][22] ),
    .A3(\design_top.MEM[11][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22541_ (.A0(\design_top.MEM[12][22] ),
    .A1(\design_top.MEM[13][22] ),
    .A2(\design_top.MEM[14][22] ),
    .A3(\design_top.MEM[15][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22542_ (.A0(_03714_),
    .A1(_03715_),
    .A2(_03716_),
    .A3(_03717_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22543_ (.A0(\design_top.MEM[16][22] ),
    .A1(\design_top.MEM[17][22] ),
    .A2(\design_top.MEM[18][22] ),
    .A3(\design_top.MEM[19][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22544_ (.A0(\design_top.MEM[20][22] ),
    .A1(\design_top.MEM[21][22] ),
    .A2(\design_top.MEM[22][22] ),
    .A3(\design_top.MEM[23][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22545_ (.A0(\design_top.MEM[24][22] ),
    .A1(\design_top.MEM[25][22] ),
    .A2(\design_top.MEM[26][22] ),
    .A3(\design_top.MEM[27][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22546_ (.A0(\design_top.MEM[28][22] ),
    .A1(\design_top.MEM[29][22] ),
    .A2(\design_top.MEM[30][22] ),
    .A3(\design_top.MEM[31][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22547_ (.A0(_03719_),
    .A1(_03720_),
    .A2(_03721_),
    .A3(_03722_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22548_ (.A0(\design_top.MEM[32][22] ),
    .A1(\design_top.MEM[33][22] ),
    .A2(\design_top.MEM[34][22] ),
    .A3(\design_top.MEM[35][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22549_ (.A0(\design_top.MEM[36][22] ),
    .A1(\design_top.MEM[37][22] ),
    .A2(\design_top.MEM[38][22] ),
    .A3(\design_top.MEM[39][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22550_ (.A0(\design_top.MEM[40][22] ),
    .A1(\design_top.MEM[41][22] ),
    .A2(\design_top.MEM[42][22] ),
    .A3(\design_top.MEM[43][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22551_ (.A0(\design_top.MEM[44][22] ),
    .A1(\design_top.MEM[45][22] ),
    .A2(\design_top.MEM[46][22] ),
    .A3(\design_top.MEM[47][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22552_ (.A0(_03724_),
    .A1(_03725_),
    .A2(_03726_),
    .A3(_03727_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22553_ (.A0(\design_top.MEM[48][22] ),
    .A1(\design_top.MEM[49][22] ),
    .A2(\design_top.MEM[50][22] ),
    .A3(\design_top.MEM[51][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22554_ (.A0(\design_top.MEM[52][22] ),
    .A1(\design_top.MEM[53][22] ),
    .A2(\design_top.MEM[54][22] ),
    .A3(\design_top.MEM[55][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22555_ (.A0(\design_top.MEM[56][22] ),
    .A1(\design_top.MEM[57][22] ),
    .A2(\design_top.MEM[58][22] ),
    .A3(\design_top.MEM[59][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22556_ (.A0(\design_top.MEM[60][22] ),
    .A1(\design_top.MEM[61][22] ),
    .A2(\design_top.MEM[62][22] ),
    .A3(\design_top.MEM[63][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22557_ (.A0(_03729_),
    .A1(_03730_),
    .A2(_03731_),
    .A3(_03732_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22558_ (.A0(_03718_),
    .A1(_03723_),
    .A2(_03728_),
    .A3(_03733_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22559_ (.A0(\design_top.MEM[0][21] ),
    .A1(\design_top.MEM[1][21] ),
    .A2(\design_top.MEM[2][21] ),
    .A3(\design_top.MEM[3][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22560_ (.A0(\design_top.MEM[4][21] ),
    .A1(\design_top.MEM[5][21] ),
    .A2(\design_top.MEM[6][21] ),
    .A3(\design_top.MEM[7][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22561_ (.A0(\design_top.MEM[8][21] ),
    .A1(\design_top.MEM[9][21] ),
    .A2(\design_top.MEM[10][21] ),
    .A3(\design_top.MEM[11][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22562_ (.A0(\design_top.MEM[12][21] ),
    .A1(\design_top.MEM[13][21] ),
    .A2(\design_top.MEM[14][21] ),
    .A3(\design_top.MEM[15][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22563_ (.A0(_03694_),
    .A1(_03695_),
    .A2(_03696_),
    .A3(_03697_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22564_ (.A0(\design_top.MEM[16][21] ),
    .A1(\design_top.MEM[17][21] ),
    .A2(\design_top.MEM[18][21] ),
    .A3(\design_top.MEM[19][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22565_ (.A0(\design_top.MEM[20][21] ),
    .A1(\design_top.MEM[21][21] ),
    .A2(\design_top.MEM[22][21] ),
    .A3(\design_top.MEM[23][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22566_ (.A0(\design_top.MEM[24][21] ),
    .A1(\design_top.MEM[25][21] ),
    .A2(\design_top.MEM[26][21] ),
    .A3(\design_top.MEM[27][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22567_ (.A0(\design_top.MEM[28][21] ),
    .A1(\design_top.MEM[29][21] ),
    .A2(\design_top.MEM[30][21] ),
    .A3(\design_top.MEM[31][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22568_ (.A0(_03699_),
    .A1(_03700_),
    .A2(_03701_),
    .A3(_03702_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22569_ (.A0(\design_top.MEM[32][21] ),
    .A1(\design_top.MEM[33][21] ),
    .A2(\design_top.MEM[34][21] ),
    .A3(\design_top.MEM[35][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22570_ (.A0(\design_top.MEM[36][21] ),
    .A1(\design_top.MEM[37][21] ),
    .A2(\design_top.MEM[38][21] ),
    .A3(\design_top.MEM[39][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22571_ (.A0(\design_top.MEM[40][21] ),
    .A1(\design_top.MEM[41][21] ),
    .A2(\design_top.MEM[42][21] ),
    .A3(\design_top.MEM[43][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22572_ (.A0(\design_top.MEM[44][21] ),
    .A1(\design_top.MEM[45][21] ),
    .A2(\design_top.MEM[46][21] ),
    .A3(\design_top.MEM[47][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22573_ (.A0(_03704_),
    .A1(_03705_),
    .A2(_03706_),
    .A3(_03707_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22574_ (.A0(\design_top.MEM[48][21] ),
    .A1(\design_top.MEM[49][21] ),
    .A2(\design_top.MEM[50][21] ),
    .A3(\design_top.MEM[51][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22575_ (.A0(\design_top.MEM[52][21] ),
    .A1(\design_top.MEM[53][21] ),
    .A2(\design_top.MEM[54][21] ),
    .A3(\design_top.MEM[55][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22576_ (.A0(\design_top.MEM[56][21] ),
    .A1(\design_top.MEM[57][21] ),
    .A2(\design_top.MEM[58][21] ),
    .A3(\design_top.MEM[59][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22577_ (.A0(\design_top.MEM[60][21] ),
    .A1(\design_top.MEM[61][21] ),
    .A2(\design_top.MEM[62][21] ),
    .A3(\design_top.MEM[63][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22578_ (.A0(_03709_),
    .A1(_03710_),
    .A2(_03711_),
    .A3(_03712_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22579_ (.A0(_03698_),
    .A1(_03703_),
    .A2(_03708_),
    .A3(_03713_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22580_ (.A0(\design_top.MEM[0][20] ),
    .A1(\design_top.MEM[1][20] ),
    .A2(\design_top.MEM[2][20] ),
    .A3(\design_top.MEM[3][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22581_ (.A0(\design_top.MEM[4][20] ),
    .A1(\design_top.MEM[5][20] ),
    .A2(\design_top.MEM[6][20] ),
    .A3(\design_top.MEM[7][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22582_ (.A0(\design_top.MEM[8][20] ),
    .A1(\design_top.MEM[9][20] ),
    .A2(\design_top.MEM[10][20] ),
    .A3(\design_top.MEM[11][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22583_ (.A0(\design_top.MEM[12][20] ),
    .A1(\design_top.MEM[13][20] ),
    .A2(\design_top.MEM[14][20] ),
    .A3(\design_top.MEM[15][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22584_ (.A0(_03674_),
    .A1(_03675_),
    .A2(_03676_),
    .A3(_03677_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22585_ (.A0(\design_top.MEM[16][20] ),
    .A1(\design_top.MEM[17][20] ),
    .A2(\design_top.MEM[18][20] ),
    .A3(\design_top.MEM[19][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22586_ (.A0(\design_top.MEM[20][20] ),
    .A1(\design_top.MEM[21][20] ),
    .A2(\design_top.MEM[22][20] ),
    .A3(\design_top.MEM[23][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22587_ (.A0(\design_top.MEM[24][20] ),
    .A1(\design_top.MEM[25][20] ),
    .A2(\design_top.MEM[26][20] ),
    .A3(\design_top.MEM[27][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22588_ (.A0(\design_top.MEM[28][20] ),
    .A1(\design_top.MEM[29][20] ),
    .A2(\design_top.MEM[30][20] ),
    .A3(\design_top.MEM[31][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22589_ (.A0(_03679_),
    .A1(_03680_),
    .A2(_03681_),
    .A3(_03682_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22590_ (.A0(\design_top.MEM[32][20] ),
    .A1(\design_top.MEM[33][20] ),
    .A2(\design_top.MEM[34][20] ),
    .A3(\design_top.MEM[35][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22591_ (.A0(\design_top.MEM[36][20] ),
    .A1(\design_top.MEM[37][20] ),
    .A2(\design_top.MEM[38][20] ),
    .A3(\design_top.MEM[39][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22592_ (.A0(\design_top.MEM[40][20] ),
    .A1(\design_top.MEM[41][20] ),
    .A2(\design_top.MEM[42][20] ),
    .A3(\design_top.MEM[43][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22593_ (.A0(\design_top.MEM[44][20] ),
    .A1(\design_top.MEM[45][20] ),
    .A2(\design_top.MEM[46][20] ),
    .A3(\design_top.MEM[47][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22594_ (.A0(_03684_),
    .A1(_03685_),
    .A2(_03686_),
    .A3(_03687_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22595_ (.A0(\design_top.MEM[48][20] ),
    .A1(\design_top.MEM[49][20] ),
    .A2(\design_top.MEM[50][20] ),
    .A3(\design_top.MEM[51][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22596_ (.A0(\design_top.MEM[52][20] ),
    .A1(\design_top.MEM[53][20] ),
    .A2(\design_top.MEM[54][20] ),
    .A3(\design_top.MEM[55][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22597_ (.A0(\design_top.MEM[56][20] ),
    .A1(\design_top.MEM[57][20] ),
    .A2(\design_top.MEM[58][20] ),
    .A3(\design_top.MEM[59][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22598_ (.A0(\design_top.MEM[60][20] ),
    .A1(\design_top.MEM[61][20] ),
    .A2(\design_top.MEM[62][20] ),
    .A3(\design_top.MEM[63][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22599_ (.A0(_03689_),
    .A1(_03690_),
    .A2(_03691_),
    .A3(_03692_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22600_ (.A0(_03678_),
    .A1(_03683_),
    .A2(_03688_),
    .A3(_03693_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22601_ (.A0(\design_top.MEM[0][19] ),
    .A1(\design_top.MEM[1][19] ),
    .A2(\design_top.MEM[2][19] ),
    .A3(\design_top.MEM[3][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22602_ (.A0(\design_top.MEM[4][19] ),
    .A1(\design_top.MEM[5][19] ),
    .A2(\design_top.MEM[6][19] ),
    .A3(\design_top.MEM[7][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22603_ (.A0(\design_top.MEM[8][19] ),
    .A1(\design_top.MEM[9][19] ),
    .A2(\design_top.MEM[10][19] ),
    .A3(\design_top.MEM[11][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22604_ (.A0(\design_top.MEM[12][19] ),
    .A1(\design_top.MEM[13][19] ),
    .A2(\design_top.MEM[14][19] ),
    .A3(\design_top.MEM[15][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22605_ (.A0(_03654_),
    .A1(_03655_),
    .A2(_03656_),
    .A3(_03657_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22606_ (.A0(\design_top.MEM[16][19] ),
    .A1(\design_top.MEM[17][19] ),
    .A2(\design_top.MEM[18][19] ),
    .A3(\design_top.MEM[19][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22607_ (.A0(\design_top.MEM[20][19] ),
    .A1(\design_top.MEM[21][19] ),
    .A2(\design_top.MEM[22][19] ),
    .A3(\design_top.MEM[23][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22608_ (.A0(\design_top.MEM[24][19] ),
    .A1(\design_top.MEM[25][19] ),
    .A2(\design_top.MEM[26][19] ),
    .A3(\design_top.MEM[27][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22609_ (.A0(\design_top.MEM[28][19] ),
    .A1(\design_top.MEM[29][19] ),
    .A2(\design_top.MEM[30][19] ),
    .A3(\design_top.MEM[31][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22610_ (.A0(_03659_),
    .A1(_03660_),
    .A2(_03661_),
    .A3(_03662_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22611_ (.A0(\design_top.MEM[32][19] ),
    .A1(\design_top.MEM[33][19] ),
    .A2(\design_top.MEM[34][19] ),
    .A3(\design_top.MEM[35][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22612_ (.A0(\design_top.MEM[36][19] ),
    .A1(\design_top.MEM[37][19] ),
    .A2(\design_top.MEM[38][19] ),
    .A3(\design_top.MEM[39][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22613_ (.A0(\design_top.MEM[40][19] ),
    .A1(\design_top.MEM[41][19] ),
    .A2(\design_top.MEM[42][19] ),
    .A3(\design_top.MEM[43][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22614_ (.A0(\design_top.MEM[44][19] ),
    .A1(\design_top.MEM[45][19] ),
    .A2(\design_top.MEM[46][19] ),
    .A3(\design_top.MEM[47][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22615_ (.A0(_03664_),
    .A1(_03665_),
    .A2(_03666_),
    .A3(_03667_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22616_ (.A0(\design_top.MEM[48][19] ),
    .A1(\design_top.MEM[49][19] ),
    .A2(\design_top.MEM[50][19] ),
    .A3(\design_top.MEM[51][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22617_ (.A0(\design_top.MEM[52][19] ),
    .A1(\design_top.MEM[53][19] ),
    .A2(\design_top.MEM[54][19] ),
    .A3(\design_top.MEM[55][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22618_ (.A0(\design_top.MEM[56][19] ),
    .A1(\design_top.MEM[57][19] ),
    .A2(\design_top.MEM[58][19] ),
    .A3(\design_top.MEM[59][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22619_ (.A0(\design_top.MEM[60][19] ),
    .A1(\design_top.MEM[61][19] ),
    .A2(\design_top.MEM[62][19] ),
    .A3(\design_top.MEM[63][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22620_ (.A0(_03669_),
    .A1(_03670_),
    .A2(_03671_),
    .A3(_03672_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22621_ (.A0(_03658_),
    .A1(_03663_),
    .A2(_03668_),
    .A3(_03673_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22622_ (.A0(\design_top.MEM[0][18] ),
    .A1(\design_top.MEM[1][18] ),
    .A2(\design_top.MEM[2][18] ),
    .A3(\design_top.MEM[3][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22623_ (.A0(\design_top.MEM[4][18] ),
    .A1(\design_top.MEM[5][18] ),
    .A2(\design_top.MEM[6][18] ),
    .A3(\design_top.MEM[7][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22624_ (.A0(\design_top.MEM[8][18] ),
    .A1(\design_top.MEM[9][18] ),
    .A2(\design_top.MEM[10][18] ),
    .A3(\design_top.MEM[11][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22625_ (.A0(\design_top.MEM[12][18] ),
    .A1(\design_top.MEM[13][18] ),
    .A2(\design_top.MEM[14][18] ),
    .A3(\design_top.MEM[15][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22626_ (.A0(_03634_),
    .A1(_03635_),
    .A2(_03636_),
    .A3(_03637_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22627_ (.A0(\design_top.MEM[16][18] ),
    .A1(\design_top.MEM[17][18] ),
    .A2(\design_top.MEM[18][18] ),
    .A3(\design_top.MEM[19][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22628_ (.A0(\design_top.MEM[20][18] ),
    .A1(\design_top.MEM[21][18] ),
    .A2(\design_top.MEM[22][18] ),
    .A3(\design_top.MEM[23][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22629_ (.A0(\design_top.MEM[24][18] ),
    .A1(\design_top.MEM[25][18] ),
    .A2(\design_top.MEM[26][18] ),
    .A3(\design_top.MEM[27][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22630_ (.A0(\design_top.MEM[28][18] ),
    .A1(\design_top.MEM[29][18] ),
    .A2(\design_top.MEM[30][18] ),
    .A3(\design_top.MEM[31][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22631_ (.A0(_03639_),
    .A1(_03640_),
    .A2(_03641_),
    .A3(_03642_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22632_ (.A0(\design_top.MEM[32][18] ),
    .A1(\design_top.MEM[33][18] ),
    .A2(\design_top.MEM[34][18] ),
    .A3(\design_top.MEM[35][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22633_ (.A0(\design_top.MEM[36][18] ),
    .A1(\design_top.MEM[37][18] ),
    .A2(\design_top.MEM[38][18] ),
    .A3(\design_top.MEM[39][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22634_ (.A0(\design_top.MEM[40][18] ),
    .A1(\design_top.MEM[41][18] ),
    .A2(\design_top.MEM[42][18] ),
    .A3(\design_top.MEM[43][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22635_ (.A0(\design_top.MEM[44][18] ),
    .A1(\design_top.MEM[45][18] ),
    .A2(\design_top.MEM[46][18] ),
    .A3(\design_top.MEM[47][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22636_ (.A0(_03644_),
    .A1(_03645_),
    .A2(_03646_),
    .A3(_03647_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22637_ (.A0(\design_top.MEM[48][18] ),
    .A1(\design_top.MEM[49][18] ),
    .A2(\design_top.MEM[50][18] ),
    .A3(\design_top.MEM[51][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22638_ (.A0(\design_top.MEM[52][18] ),
    .A1(\design_top.MEM[53][18] ),
    .A2(\design_top.MEM[54][18] ),
    .A3(\design_top.MEM[55][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22639_ (.A0(\design_top.MEM[56][18] ),
    .A1(\design_top.MEM[57][18] ),
    .A2(\design_top.MEM[58][18] ),
    .A3(\design_top.MEM[59][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22640_ (.A0(\design_top.MEM[60][18] ),
    .A1(\design_top.MEM[61][18] ),
    .A2(\design_top.MEM[62][18] ),
    .A3(\design_top.MEM[63][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22641_ (.A0(_03649_),
    .A1(_03650_),
    .A2(_03651_),
    .A3(_03652_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22642_ (.A0(_03638_),
    .A1(_03643_),
    .A2(_03648_),
    .A3(_03653_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22643_ (.A0(\design_top.MEM[0][17] ),
    .A1(\design_top.MEM[1][17] ),
    .A2(\design_top.MEM[2][17] ),
    .A3(\design_top.MEM[3][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22644_ (.A0(\design_top.MEM[4][17] ),
    .A1(\design_top.MEM[5][17] ),
    .A2(\design_top.MEM[6][17] ),
    .A3(\design_top.MEM[7][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22645_ (.A0(\design_top.MEM[8][17] ),
    .A1(\design_top.MEM[9][17] ),
    .A2(\design_top.MEM[10][17] ),
    .A3(\design_top.MEM[11][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22646_ (.A0(\design_top.MEM[12][17] ),
    .A1(\design_top.MEM[13][17] ),
    .A2(\design_top.MEM[14][17] ),
    .A3(\design_top.MEM[15][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22647_ (.A0(_03614_),
    .A1(_03615_),
    .A2(_03616_),
    .A3(_03617_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22648_ (.A0(\design_top.MEM[16][17] ),
    .A1(\design_top.MEM[17][17] ),
    .A2(\design_top.MEM[18][17] ),
    .A3(\design_top.MEM[19][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22649_ (.A0(\design_top.MEM[20][17] ),
    .A1(\design_top.MEM[21][17] ),
    .A2(\design_top.MEM[22][17] ),
    .A3(\design_top.MEM[23][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22650_ (.A0(\design_top.MEM[24][17] ),
    .A1(\design_top.MEM[25][17] ),
    .A2(\design_top.MEM[26][17] ),
    .A3(\design_top.MEM[27][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22651_ (.A0(\design_top.MEM[28][17] ),
    .A1(\design_top.MEM[29][17] ),
    .A2(\design_top.MEM[30][17] ),
    .A3(\design_top.MEM[31][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22652_ (.A0(_03619_),
    .A1(_03620_),
    .A2(_03621_),
    .A3(_03622_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22653_ (.A0(\design_top.MEM[32][17] ),
    .A1(\design_top.MEM[33][17] ),
    .A2(\design_top.MEM[34][17] ),
    .A3(\design_top.MEM[35][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22654_ (.A0(\design_top.MEM[36][17] ),
    .A1(\design_top.MEM[37][17] ),
    .A2(\design_top.MEM[38][17] ),
    .A3(\design_top.MEM[39][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22655_ (.A0(\design_top.MEM[40][17] ),
    .A1(\design_top.MEM[41][17] ),
    .A2(\design_top.MEM[42][17] ),
    .A3(\design_top.MEM[43][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22656_ (.A0(\design_top.MEM[44][17] ),
    .A1(\design_top.MEM[45][17] ),
    .A2(\design_top.MEM[46][17] ),
    .A3(\design_top.MEM[47][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22657_ (.A0(_03624_),
    .A1(_03625_),
    .A2(_03626_),
    .A3(_03627_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22658_ (.A0(\design_top.MEM[48][17] ),
    .A1(\design_top.MEM[49][17] ),
    .A2(\design_top.MEM[50][17] ),
    .A3(\design_top.MEM[51][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22659_ (.A0(\design_top.MEM[52][17] ),
    .A1(\design_top.MEM[53][17] ),
    .A2(\design_top.MEM[54][17] ),
    .A3(\design_top.MEM[55][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22660_ (.A0(\design_top.MEM[56][17] ),
    .A1(\design_top.MEM[57][17] ),
    .A2(\design_top.MEM[58][17] ),
    .A3(\design_top.MEM[59][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22661_ (.A0(\design_top.MEM[60][17] ),
    .A1(\design_top.MEM[61][17] ),
    .A2(\design_top.MEM[62][17] ),
    .A3(\design_top.MEM[63][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22662_ (.A0(_03629_),
    .A1(_03630_),
    .A2(_03631_),
    .A3(_03632_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22663_ (.A0(_03618_),
    .A1(_03623_),
    .A2(_03628_),
    .A3(_03633_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22664_ (.A0(\design_top.MEM[0][16] ),
    .A1(\design_top.MEM[1][16] ),
    .A2(\design_top.MEM[2][16] ),
    .A3(\design_top.MEM[3][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22665_ (.A0(\design_top.MEM[4][16] ),
    .A1(\design_top.MEM[5][16] ),
    .A2(\design_top.MEM[6][16] ),
    .A3(\design_top.MEM[7][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22666_ (.A0(\design_top.MEM[8][16] ),
    .A1(\design_top.MEM[9][16] ),
    .A2(\design_top.MEM[10][16] ),
    .A3(\design_top.MEM[11][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22667_ (.A0(\design_top.MEM[12][16] ),
    .A1(\design_top.MEM[13][16] ),
    .A2(\design_top.MEM[14][16] ),
    .A3(\design_top.MEM[15][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22668_ (.A0(_03594_),
    .A1(_03595_),
    .A2(_03596_),
    .A3(_03597_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22669_ (.A0(\design_top.MEM[16][16] ),
    .A1(\design_top.MEM[17][16] ),
    .A2(\design_top.MEM[18][16] ),
    .A3(\design_top.MEM[19][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22670_ (.A0(\design_top.MEM[20][16] ),
    .A1(\design_top.MEM[21][16] ),
    .A2(\design_top.MEM[22][16] ),
    .A3(\design_top.MEM[23][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22671_ (.A0(\design_top.MEM[24][16] ),
    .A1(\design_top.MEM[25][16] ),
    .A2(\design_top.MEM[26][16] ),
    .A3(\design_top.MEM[27][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22672_ (.A0(\design_top.MEM[28][16] ),
    .A1(\design_top.MEM[29][16] ),
    .A2(\design_top.MEM[30][16] ),
    .A3(\design_top.MEM[31][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22673_ (.A0(_03599_),
    .A1(_03600_),
    .A2(_03601_),
    .A3(_03602_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22674_ (.A0(\design_top.MEM[32][16] ),
    .A1(\design_top.MEM[33][16] ),
    .A2(\design_top.MEM[34][16] ),
    .A3(\design_top.MEM[35][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22675_ (.A0(\design_top.MEM[36][16] ),
    .A1(\design_top.MEM[37][16] ),
    .A2(\design_top.MEM[38][16] ),
    .A3(\design_top.MEM[39][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22676_ (.A0(\design_top.MEM[40][16] ),
    .A1(\design_top.MEM[41][16] ),
    .A2(\design_top.MEM[42][16] ),
    .A3(\design_top.MEM[43][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22677_ (.A0(\design_top.MEM[44][16] ),
    .A1(\design_top.MEM[45][16] ),
    .A2(\design_top.MEM[46][16] ),
    .A3(\design_top.MEM[47][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22678_ (.A0(_03604_),
    .A1(_03605_),
    .A2(_03606_),
    .A3(_03607_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22679_ (.A0(\design_top.MEM[48][16] ),
    .A1(\design_top.MEM[49][16] ),
    .A2(\design_top.MEM[50][16] ),
    .A3(\design_top.MEM[51][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22680_ (.A0(\design_top.MEM[52][16] ),
    .A1(\design_top.MEM[53][16] ),
    .A2(\design_top.MEM[54][16] ),
    .A3(\design_top.MEM[55][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22681_ (.A0(\design_top.MEM[56][16] ),
    .A1(\design_top.MEM[57][16] ),
    .A2(\design_top.MEM[58][16] ),
    .A3(\design_top.MEM[59][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22682_ (.A0(\design_top.MEM[60][16] ),
    .A1(\design_top.MEM[61][16] ),
    .A2(\design_top.MEM[62][16] ),
    .A3(\design_top.MEM[63][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22683_ (.A0(_03609_),
    .A1(_03610_),
    .A2(_03611_),
    .A3(_03612_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22684_ (.A0(_03598_),
    .A1(_03603_),
    .A2(_03608_),
    .A3(_03613_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22685_ (.A0(\design_top.MEM[0][15] ),
    .A1(\design_top.MEM[1][15] ),
    .A2(\design_top.MEM[2][15] ),
    .A3(\design_top.MEM[3][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22686_ (.A0(\design_top.MEM[4][15] ),
    .A1(\design_top.MEM[5][15] ),
    .A2(\design_top.MEM[6][15] ),
    .A3(\design_top.MEM[7][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22687_ (.A0(\design_top.MEM[8][15] ),
    .A1(\design_top.MEM[9][15] ),
    .A2(\design_top.MEM[10][15] ),
    .A3(\design_top.MEM[11][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22688_ (.A0(\design_top.MEM[12][15] ),
    .A1(\design_top.MEM[13][15] ),
    .A2(\design_top.MEM[14][15] ),
    .A3(\design_top.MEM[15][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22689_ (.A0(_03574_),
    .A1(_03575_),
    .A2(_03576_),
    .A3(_03577_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22690_ (.A0(\design_top.MEM[16][15] ),
    .A1(\design_top.MEM[17][15] ),
    .A2(\design_top.MEM[18][15] ),
    .A3(\design_top.MEM[19][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22691_ (.A0(\design_top.MEM[20][15] ),
    .A1(\design_top.MEM[21][15] ),
    .A2(\design_top.MEM[22][15] ),
    .A3(\design_top.MEM[23][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22692_ (.A0(\design_top.MEM[24][15] ),
    .A1(\design_top.MEM[25][15] ),
    .A2(\design_top.MEM[26][15] ),
    .A3(\design_top.MEM[27][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22693_ (.A0(\design_top.MEM[28][15] ),
    .A1(\design_top.MEM[29][15] ),
    .A2(\design_top.MEM[30][15] ),
    .A3(\design_top.MEM[31][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22694_ (.A0(_03579_),
    .A1(_03580_),
    .A2(_03581_),
    .A3(_03582_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22695_ (.A0(\design_top.MEM[32][15] ),
    .A1(\design_top.MEM[33][15] ),
    .A2(\design_top.MEM[34][15] ),
    .A3(\design_top.MEM[35][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22696_ (.A0(\design_top.MEM[36][15] ),
    .A1(\design_top.MEM[37][15] ),
    .A2(\design_top.MEM[38][15] ),
    .A3(\design_top.MEM[39][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22697_ (.A0(\design_top.MEM[40][15] ),
    .A1(\design_top.MEM[41][15] ),
    .A2(\design_top.MEM[42][15] ),
    .A3(\design_top.MEM[43][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22698_ (.A0(\design_top.MEM[44][15] ),
    .A1(\design_top.MEM[45][15] ),
    .A2(\design_top.MEM[46][15] ),
    .A3(\design_top.MEM[47][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22699_ (.A0(_03584_),
    .A1(_03585_),
    .A2(_03586_),
    .A3(_03587_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22700_ (.A0(\design_top.MEM[48][15] ),
    .A1(\design_top.MEM[49][15] ),
    .A2(\design_top.MEM[50][15] ),
    .A3(\design_top.MEM[51][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22701_ (.A0(\design_top.MEM[52][15] ),
    .A1(\design_top.MEM[53][15] ),
    .A2(\design_top.MEM[54][15] ),
    .A3(\design_top.MEM[55][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22702_ (.A0(\design_top.MEM[56][15] ),
    .A1(\design_top.MEM[57][15] ),
    .A2(\design_top.MEM[58][15] ),
    .A3(\design_top.MEM[59][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22703_ (.A0(\design_top.MEM[60][15] ),
    .A1(\design_top.MEM[61][15] ),
    .A2(\design_top.MEM[62][15] ),
    .A3(\design_top.MEM[63][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22704_ (.A0(_03589_),
    .A1(_03590_),
    .A2(_03591_),
    .A3(_03592_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22705_ (.A0(_03578_),
    .A1(_03583_),
    .A2(_03588_),
    .A3(_03593_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22706_ (.A0(\design_top.MEM[0][14] ),
    .A1(\design_top.MEM[1][14] ),
    .A2(\design_top.MEM[2][14] ),
    .A3(\design_top.MEM[3][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22707_ (.A0(\design_top.MEM[4][14] ),
    .A1(\design_top.MEM[5][14] ),
    .A2(\design_top.MEM[6][14] ),
    .A3(\design_top.MEM[7][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22708_ (.A0(\design_top.MEM[8][14] ),
    .A1(\design_top.MEM[9][14] ),
    .A2(\design_top.MEM[10][14] ),
    .A3(\design_top.MEM[11][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22709_ (.A0(\design_top.MEM[12][14] ),
    .A1(\design_top.MEM[13][14] ),
    .A2(\design_top.MEM[14][14] ),
    .A3(\design_top.MEM[15][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22710_ (.A0(_03554_),
    .A1(_03555_),
    .A2(_03556_),
    .A3(_03557_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22711_ (.A0(\design_top.MEM[16][14] ),
    .A1(\design_top.MEM[17][14] ),
    .A2(\design_top.MEM[18][14] ),
    .A3(\design_top.MEM[19][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22712_ (.A0(\design_top.MEM[20][14] ),
    .A1(\design_top.MEM[21][14] ),
    .A2(\design_top.MEM[22][14] ),
    .A3(\design_top.MEM[23][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22713_ (.A0(\design_top.MEM[24][14] ),
    .A1(\design_top.MEM[25][14] ),
    .A2(\design_top.MEM[26][14] ),
    .A3(\design_top.MEM[27][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22714_ (.A0(\design_top.MEM[28][14] ),
    .A1(\design_top.MEM[29][14] ),
    .A2(\design_top.MEM[30][14] ),
    .A3(\design_top.MEM[31][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22715_ (.A0(_03559_),
    .A1(_03560_),
    .A2(_03561_),
    .A3(_03562_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22716_ (.A0(\design_top.MEM[32][14] ),
    .A1(\design_top.MEM[33][14] ),
    .A2(\design_top.MEM[34][14] ),
    .A3(\design_top.MEM[35][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22717_ (.A0(\design_top.MEM[36][14] ),
    .A1(\design_top.MEM[37][14] ),
    .A2(\design_top.MEM[38][14] ),
    .A3(\design_top.MEM[39][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22718_ (.A0(\design_top.MEM[40][14] ),
    .A1(\design_top.MEM[41][14] ),
    .A2(\design_top.MEM[42][14] ),
    .A3(\design_top.MEM[43][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22719_ (.A0(\design_top.MEM[44][14] ),
    .A1(\design_top.MEM[45][14] ),
    .A2(\design_top.MEM[46][14] ),
    .A3(\design_top.MEM[47][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22720_ (.A0(_03564_),
    .A1(_03565_),
    .A2(_03566_),
    .A3(_03567_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22721_ (.A0(\design_top.MEM[48][14] ),
    .A1(\design_top.MEM[49][14] ),
    .A2(\design_top.MEM[50][14] ),
    .A3(\design_top.MEM[51][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22722_ (.A0(\design_top.MEM[52][14] ),
    .A1(\design_top.MEM[53][14] ),
    .A2(\design_top.MEM[54][14] ),
    .A3(\design_top.MEM[55][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22723_ (.A0(\design_top.MEM[56][14] ),
    .A1(\design_top.MEM[57][14] ),
    .A2(\design_top.MEM[58][14] ),
    .A3(\design_top.MEM[59][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22724_ (.A0(\design_top.MEM[60][14] ),
    .A1(\design_top.MEM[61][14] ),
    .A2(\design_top.MEM[62][14] ),
    .A3(\design_top.MEM[63][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22725_ (.A0(_03569_),
    .A1(_03570_),
    .A2(_03571_),
    .A3(_03572_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22726_ (.A0(_03558_),
    .A1(_03563_),
    .A2(_03568_),
    .A3(_03573_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22727_ (.A0(\design_top.MEM[0][13] ),
    .A1(\design_top.MEM[1][13] ),
    .A2(\design_top.MEM[2][13] ),
    .A3(\design_top.MEM[3][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22728_ (.A0(\design_top.MEM[4][13] ),
    .A1(\design_top.MEM[5][13] ),
    .A2(\design_top.MEM[6][13] ),
    .A3(\design_top.MEM[7][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22729_ (.A0(\design_top.MEM[8][13] ),
    .A1(\design_top.MEM[9][13] ),
    .A2(\design_top.MEM[10][13] ),
    .A3(\design_top.MEM[11][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22730_ (.A0(\design_top.MEM[12][13] ),
    .A1(\design_top.MEM[13][13] ),
    .A2(\design_top.MEM[14][13] ),
    .A3(\design_top.MEM[15][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22731_ (.A0(_03534_),
    .A1(_03535_),
    .A2(_03536_),
    .A3(_03537_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22732_ (.A0(\design_top.MEM[16][13] ),
    .A1(\design_top.MEM[17][13] ),
    .A2(\design_top.MEM[18][13] ),
    .A3(\design_top.MEM[19][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22733_ (.A0(\design_top.MEM[20][13] ),
    .A1(\design_top.MEM[21][13] ),
    .A2(\design_top.MEM[22][13] ),
    .A3(\design_top.MEM[23][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22734_ (.A0(\design_top.MEM[24][13] ),
    .A1(\design_top.MEM[25][13] ),
    .A2(\design_top.MEM[26][13] ),
    .A3(\design_top.MEM[27][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22735_ (.A0(\design_top.MEM[28][13] ),
    .A1(\design_top.MEM[29][13] ),
    .A2(\design_top.MEM[30][13] ),
    .A3(\design_top.MEM[31][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22736_ (.A0(_03539_),
    .A1(_03540_),
    .A2(_03541_),
    .A3(_03542_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22737_ (.A0(\design_top.MEM[32][13] ),
    .A1(\design_top.MEM[33][13] ),
    .A2(\design_top.MEM[34][13] ),
    .A3(\design_top.MEM[35][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22738_ (.A0(\design_top.MEM[36][13] ),
    .A1(\design_top.MEM[37][13] ),
    .A2(\design_top.MEM[38][13] ),
    .A3(\design_top.MEM[39][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22739_ (.A0(\design_top.MEM[40][13] ),
    .A1(\design_top.MEM[41][13] ),
    .A2(\design_top.MEM[42][13] ),
    .A3(\design_top.MEM[43][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22740_ (.A0(\design_top.MEM[44][13] ),
    .A1(\design_top.MEM[45][13] ),
    .A2(\design_top.MEM[46][13] ),
    .A3(\design_top.MEM[47][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22741_ (.A0(_03544_),
    .A1(_03545_),
    .A2(_03546_),
    .A3(_03547_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22742_ (.A0(\design_top.MEM[48][13] ),
    .A1(\design_top.MEM[49][13] ),
    .A2(\design_top.MEM[50][13] ),
    .A3(\design_top.MEM[51][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22743_ (.A0(\design_top.MEM[52][13] ),
    .A1(\design_top.MEM[53][13] ),
    .A2(\design_top.MEM[54][13] ),
    .A3(\design_top.MEM[55][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22744_ (.A0(\design_top.MEM[56][13] ),
    .A1(\design_top.MEM[57][13] ),
    .A2(\design_top.MEM[58][13] ),
    .A3(\design_top.MEM[59][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22745_ (.A0(\design_top.MEM[60][13] ),
    .A1(\design_top.MEM[61][13] ),
    .A2(\design_top.MEM[62][13] ),
    .A3(\design_top.MEM[63][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22746_ (.A0(_03549_),
    .A1(_03550_),
    .A2(_03551_),
    .A3(_03552_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22747_ (.A0(_03538_),
    .A1(_03543_),
    .A2(_03548_),
    .A3(_03553_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22748_ (.A0(\design_top.MEM[0][12] ),
    .A1(\design_top.MEM[1][12] ),
    .A2(\design_top.MEM[2][12] ),
    .A3(\design_top.MEM[3][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22749_ (.A0(\design_top.MEM[4][12] ),
    .A1(\design_top.MEM[5][12] ),
    .A2(\design_top.MEM[6][12] ),
    .A3(\design_top.MEM[7][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22750_ (.A0(\design_top.MEM[8][12] ),
    .A1(\design_top.MEM[9][12] ),
    .A2(\design_top.MEM[10][12] ),
    .A3(\design_top.MEM[11][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22751_ (.A0(\design_top.MEM[12][12] ),
    .A1(\design_top.MEM[13][12] ),
    .A2(\design_top.MEM[14][12] ),
    .A3(\design_top.MEM[15][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22752_ (.A0(_03514_),
    .A1(_03515_),
    .A2(_03516_),
    .A3(_03517_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22753_ (.A0(\design_top.MEM[16][12] ),
    .A1(\design_top.MEM[17][12] ),
    .A2(\design_top.MEM[18][12] ),
    .A3(\design_top.MEM[19][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22754_ (.A0(\design_top.MEM[20][12] ),
    .A1(\design_top.MEM[21][12] ),
    .A2(\design_top.MEM[22][12] ),
    .A3(\design_top.MEM[23][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22755_ (.A0(\design_top.MEM[24][12] ),
    .A1(\design_top.MEM[25][12] ),
    .A2(\design_top.MEM[26][12] ),
    .A3(\design_top.MEM[27][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22756_ (.A0(\design_top.MEM[28][12] ),
    .A1(\design_top.MEM[29][12] ),
    .A2(\design_top.MEM[30][12] ),
    .A3(\design_top.MEM[31][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22757_ (.A0(_03519_),
    .A1(_03520_),
    .A2(_03521_),
    .A3(_03522_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22758_ (.A0(\design_top.MEM[32][12] ),
    .A1(\design_top.MEM[33][12] ),
    .A2(\design_top.MEM[34][12] ),
    .A3(\design_top.MEM[35][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22759_ (.A0(\design_top.MEM[36][12] ),
    .A1(\design_top.MEM[37][12] ),
    .A2(\design_top.MEM[38][12] ),
    .A3(\design_top.MEM[39][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22760_ (.A0(\design_top.MEM[40][12] ),
    .A1(\design_top.MEM[41][12] ),
    .A2(\design_top.MEM[42][12] ),
    .A3(\design_top.MEM[43][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22761_ (.A0(\design_top.MEM[44][12] ),
    .A1(\design_top.MEM[45][12] ),
    .A2(\design_top.MEM[46][12] ),
    .A3(\design_top.MEM[47][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22762_ (.A0(_03524_),
    .A1(_03525_),
    .A2(_03526_),
    .A3(_03527_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22763_ (.A0(\design_top.MEM[48][12] ),
    .A1(\design_top.MEM[49][12] ),
    .A2(\design_top.MEM[50][12] ),
    .A3(\design_top.MEM[51][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22764_ (.A0(\design_top.MEM[52][12] ),
    .A1(\design_top.MEM[53][12] ),
    .A2(\design_top.MEM[54][12] ),
    .A3(\design_top.MEM[55][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22765_ (.A0(\design_top.MEM[56][12] ),
    .A1(\design_top.MEM[57][12] ),
    .A2(\design_top.MEM[58][12] ),
    .A3(\design_top.MEM[59][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22766_ (.A0(\design_top.MEM[60][12] ),
    .A1(\design_top.MEM[61][12] ),
    .A2(\design_top.MEM[62][12] ),
    .A3(\design_top.MEM[63][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22767_ (.A0(_03529_),
    .A1(_03530_),
    .A2(_03531_),
    .A3(_03532_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22768_ (.A0(_03518_),
    .A1(_03523_),
    .A2(_03528_),
    .A3(_03533_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22769_ (.A0(\design_top.MEM[0][11] ),
    .A1(\design_top.MEM[1][11] ),
    .A2(\design_top.MEM[2][11] ),
    .A3(\design_top.MEM[3][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22770_ (.A0(\design_top.MEM[4][11] ),
    .A1(\design_top.MEM[5][11] ),
    .A2(\design_top.MEM[6][11] ),
    .A3(\design_top.MEM[7][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22771_ (.A0(\design_top.MEM[8][11] ),
    .A1(\design_top.MEM[9][11] ),
    .A2(\design_top.MEM[10][11] ),
    .A3(\design_top.MEM[11][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22772_ (.A0(\design_top.MEM[12][11] ),
    .A1(\design_top.MEM[13][11] ),
    .A2(\design_top.MEM[14][11] ),
    .A3(\design_top.MEM[15][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22773_ (.A0(_03494_),
    .A1(_03495_),
    .A2(_03496_),
    .A3(_03497_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22774_ (.A0(\design_top.MEM[16][11] ),
    .A1(\design_top.MEM[17][11] ),
    .A2(\design_top.MEM[18][11] ),
    .A3(\design_top.MEM[19][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22775_ (.A0(\design_top.MEM[20][11] ),
    .A1(\design_top.MEM[21][11] ),
    .A2(\design_top.MEM[22][11] ),
    .A3(\design_top.MEM[23][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22776_ (.A0(\design_top.MEM[24][11] ),
    .A1(\design_top.MEM[25][11] ),
    .A2(\design_top.MEM[26][11] ),
    .A3(\design_top.MEM[27][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22777_ (.A0(\design_top.MEM[28][11] ),
    .A1(\design_top.MEM[29][11] ),
    .A2(\design_top.MEM[30][11] ),
    .A3(\design_top.MEM[31][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22778_ (.A0(_03499_),
    .A1(_03500_),
    .A2(_03501_),
    .A3(_03502_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22779_ (.A0(\design_top.MEM[32][11] ),
    .A1(\design_top.MEM[33][11] ),
    .A2(\design_top.MEM[34][11] ),
    .A3(\design_top.MEM[35][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22780_ (.A0(\design_top.MEM[36][11] ),
    .A1(\design_top.MEM[37][11] ),
    .A2(\design_top.MEM[38][11] ),
    .A3(\design_top.MEM[39][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22781_ (.A0(\design_top.MEM[40][11] ),
    .A1(\design_top.MEM[41][11] ),
    .A2(\design_top.MEM[42][11] ),
    .A3(\design_top.MEM[43][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22782_ (.A0(\design_top.MEM[44][11] ),
    .A1(\design_top.MEM[45][11] ),
    .A2(\design_top.MEM[46][11] ),
    .A3(\design_top.MEM[47][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22783_ (.A0(_03504_),
    .A1(_03505_),
    .A2(_03506_),
    .A3(_03507_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22784_ (.A0(\design_top.MEM[48][11] ),
    .A1(\design_top.MEM[49][11] ),
    .A2(\design_top.MEM[50][11] ),
    .A3(\design_top.MEM[51][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22785_ (.A0(\design_top.MEM[52][11] ),
    .A1(\design_top.MEM[53][11] ),
    .A2(\design_top.MEM[54][11] ),
    .A3(\design_top.MEM[55][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22786_ (.A0(\design_top.MEM[56][11] ),
    .A1(\design_top.MEM[57][11] ),
    .A2(\design_top.MEM[58][11] ),
    .A3(\design_top.MEM[59][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22787_ (.A0(\design_top.MEM[60][11] ),
    .A1(\design_top.MEM[61][11] ),
    .A2(\design_top.MEM[62][11] ),
    .A3(\design_top.MEM[63][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22788_ (.A0(_03509_),
    .A1(_03510_),
    .A2(_03511_),
    .A3(_03512_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22789_ (.A0(_03498_),
    .A1(_03503_),
    .A2(_03508_),
    .A3(_03513_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22790_ (.A0(\design_top.MEM[0][10] ),
    .A1(\design_top.MEM[1][10] ),
    .A2(\design_top.MEM[2][10] ),
    .A3(\design_top.MEM[3][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22791_ (.A0(\design_top.MEM[4][10] ),
    .A1(\design_top.MEM[5][10] ),
    .A2(\design_top.MEM[6][10] ),
    .A3(\design_top.MEM[7][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22792_ (.A0(\design_top.MEM[8][10] ),
    .A1(\design_top.MEM[9][10] ),
    .A2(\design_top.MEM[10][10] ),
    .A3(\design_top.MEM[11][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22793_ (.A0(\design_top.MEM[12][10] ),
    .A1(\design_top.MEM[13][10] ),
    .A2(\design_top.MEM[14][10] ),
    .A3(\design_top.MEM[15][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22794_ (.A0(_03474_),
    .A1(_03475_),
    .A2(_03476_),
    .A3(_03477_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22795_ (.A0(\design_top.MEM[16][10] ),
    .A1(\design_top.MEM[17][10] ),
    .A2(\design_top.MEM[18][10] ),
    .A3(\design_top.MEM[19][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22796_ (.A0(\design_top.MEM[20][10] ),
    .A1(\design_top.MEM[21][10] ),
    .A2(\design_top.MEM[22][10] ),
    .A3(\design_top.MEM[23][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22797_ (.A0(\design_top.MEM[24][10] ),
    .A1(\design_top.MEM[25][10] ),
    .A2(\design_top.MEM[26][10] ),
    .A3(\design_top.MEM[27][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22798_ (.A0(\design_top.MEM[28][10] ),
    .A1(\design_top.MEM[29][10] ),
    .A2(\design_top.MEM[30][10] ),
    .A3(\design_top.MEM[31][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22799_ (.A0(_03479_),
    .A1(_03480_),
    .A2(_03481_),
    .A3(_03482_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22800_ (.A0(\design_top.MEM[32][10] ),
    .A1(\design_top.MEM[33][10] ),
    .A2(\design_top.MEM[34][10] ),
    .A3(\design_top.MEM[35][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22801_ (.A0(\design_top.MEM[36][10] ),
    .A1(\design_top.MEM[37][10] ),
    .A2(\design_top.MEM[38][10] ),
    .A3(\design_top.MEM[39][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22802_ (.A0(\design_top.MEM[40][10] ),
    .A1(\design_top.MEM[41][10] ),
    .A2(\design_top.MEM[42][10] ),
    .A3(\design_top.MEM[43][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22803_ (.A0(\design_top.MEM[44][10] ),
    .A1(\design_top.MEM[45][10] ),
    .A2(\design_top.MEM[46][10] ),
    .A3(\design_top.MEM[47][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22804_ (.A0(_03484_),
    .A1(_03485_),
    .A2(_03486_),
    .A3(_03487_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22805_ (.A0(\design_top.MEM[48][10] ),
    .A1(\design_top.MEM[49][10] ),
    .A2(\design_top.MEM[50][10] ),
    .A3(\design_top.MEM[51][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22806_ (.A0(\design_top.MEM[52][10] ),
    .A1(\design_top.MEM[53][10] ),
    .A2(\design_top.MEM[54][10] ),
    .A3(\design_top.MEM[55][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22807_ (.A0(\design_top.MEM[56][10] ),
    .A1(\design_top.MEM[57][10] ),
    .A2(\design_top.MEM[58][10] ),
    .A3(\design_top.MEM[59][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22808_ (.A0(\design_top.MEM[60][10] ),
    .A1(\design_top.MEM[61][10] ),
    .A2(\design_top.MEM[62][10] ),
    .A3(\design_top.MEM[63][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22809_ (.A0(_03489_),
    .A1(_03490_),
    .A2(_03491_),
    .A3(_03492_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22810_ (.A0(_03478_),
    .A1(_03483_),
    .A2(_03488_),
    .A3(_03493_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22811_ (.A0(\design_top.MEM[0][9] ),
    .A1(\design_top.MEM[1][9] ),
    .A2(\design_top.MEM[2][9] ),
    .A3(\design_top.MEM[3][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22812_ (.A0(\design_top.MEM[4][9] ),
    .A1(\design_top.MEM[5][9] ),
    .A2(\design_top.MEM[6][9] ),
    .A3(\design_top.MEM[7][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22813_ (.A0(\design_top.MEM[8][9] ),
    .A1(\design_top.MEM[9][9] ),
    .A2(\design_top.MEM[10][9] ),
    .A3(\design_top.MEM[11][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22814_ (.A0(\design_top.MEM[12][9] ),
    .A1(\design_top.MEM[13][9] ),
    .A2(\design_top.MEM[14][9] ),
    .A3(\design_top.MEM[15][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22815_ (.A0(_03454_),
    .A1(_03455_),
    .A2(_03456_),
    .A3(_03457_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22816_ (.A0(\design_top.MEM[16][9] ),
    .A1(\design_top.MEM[17][9] ),
    .A2(\design_top.MEM[18][9] ),
    .A3(\design_top.MEM[19][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22817_ (.A0(\design_top.MEM[20][9] ),
    .A1(\design_top.MEM[21][9] ),
    .A2(\design_top.MEM[22][9] ),
    .A3(\design_top.MEM[23][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22818_ (.A0(\design_top.MEM[24][9] ),
    .A1(\design_top.MEM[25][9] ),
    .A2(\design_top.MEM[26][9] ),
    .A3(\design_top.MEM[27][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22819_ (.A0(\design_top.MEM[28][9] ),
    .A1(\design_top.MEM[29][9] ),
    .A2(\design_top.MEM[30][9] ),
    .A3(\design_top.MEM[31][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22820_ (.A0(_03459_),
    .A1(_03460_),
    .A2(_03461_),
    .A3(_03462_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22821_ (.A0(\design_top.MEM[32][9] ),
    .A1(\design_top.MEM[33][9] ),
    .A2(\design_top.MEM[34][9] ),
    .A3(\design_top.MEM[35][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22822_ (.A0(\design_top.MEM[36][9] ),
    .A1(\design_top.MEM[37][9] ),
    .A2(\design_top.MEM[38][9] ),
    .A3(\design_top.MEM[39][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22823_ (.A0(\design_top.MEM[40][9] ),
    .A1(\design_top.MEM[41][9] ),
    .A2(\design_top.MEM[42][9] ),
    .A3(\design_top.MEM[43][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22824_ (.A0(\design_top.MEM[44][9] ),
    .A1(\design_top.MEM[45][9] ),
    .A2(\design_top.MEM[46][9] ),
    .A3(\design_top.MEM[47][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22825_ (.A0(_03464_),
    .A1(_03465_),
    .A2(_03466_),
    .A3(_03467_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22826_ (.A0(\design_top.MEM[48][9] ),
    .A1(\design_top.MEM[49][9] ),
    .A2(\design_top.MEM[50][9] ),
    .A3(\design_top.MEM[51][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22827_ (.A0(\design_top.MEM[52][9] ),
    .A1(\design_top.MEM[53][9] ),
    .A2(\design_top.MEM[54][9] ),
    .A3(\design_top.MEM[55][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22828_ (.A0(\design_top.MEM[56][9] ),
    .A1(\design_top.MEM[57][9] ),
    .A2(\design_top.MEM[58][9] ),
    .A3(\design_top.MEM[59][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22829_ (.A0(\design_top.MEM[60][9] ),
    .A1(\design_top.MEM[61][9] ),
    .A2(\design_top.MEM[62][9] ),
    .A3(\design_top.MEM[63][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22830_ (.A0(_03469_),
    .A1(_03470_),
    .A2(_03471_),
    .A3(_03472_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22831_ (.A0(_03458_),
    .A1(_03463_),
    .A2(_03468_),
    .A3(_03473_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22832_ (.A0(\design_top.MEM[0][8] ),
    .A1(\design_top.MEM[1][8] ),
    .A2(\design_top.MEM[2][8] ),
    .A3(\design_top.MEM[3][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22833_ (.A0(\design_top.MEM[4][8] ),
    .A1(\design_top.MEM[5][8] ),
    .A2(\design_top.MEM[6][8] ),
    .A3(\design_top.MEM[7][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22834_ (.A0(\design_top.MEM[8][8] ),
    .A1(\design_top.MEM[9][8] ),
    .A2(\design_top.MEM[10][8] ),
    .A3(\design_top.MEM[11][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22835_ (.A0(\design_top.MEM[12][8] ),
    .A1(\design_top.MEM[13][8] ),
    .A2(\design_top.MEM[14][8] ),
    .A3(\design_top.MEM[15][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22836_ (.A0(_03434_),
    .A1(_03435_),
    .A2(_03436_),
    .A3(_03437_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22837_ (.A0(\design_top.MEM[16][8] ),
    .A1(\design_top.MEM[17][8] ),
    .A2(\design_top.MEM[18][8] ),
    .A3(\design_top.MEM[19][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22838_ (.A0(\design_top.MEM[20][8] ),
    .A1(\design_top.MEM[21][8] ),
    .A2(\design_top.MEM[22][8] ),
    .A3(\design_top.MEM[23][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22839_ (.A0(\design_top.MEM[24][8] ),
    .A1(\design_top.MEM[25][8] ),
    .A2(\design_top.MEM[26][8] ),
    .A3(\design_top.MEM[27][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22840_ (.A0(\design_top.MEM[28][8] ),
    .A1(\design_top.MEM[29][8] ),
    .A2(\design_top.MEM[30][8] ),
    .A3(\design_top.MEM[31][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22841_ (.A0(_03439_),
    .A1(_03440_),
    .A2(_03441_),
    .A3(_03442_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22842_ (.A0(\design_top.MEM[32][8] ),
    .A1(\design_top.MEM[33][8] ),
    .A2(\design_top.MEM[34][8] ),
    .A3(\design_top.MEM[35][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22843_ (.A0(\design_top.MEM[36][8] ),
    .A1(\design_top.MEM[37][8] ),
    .A2(\design_top.MEM[38][8] ),
    .A3(\design_top.MEM[39][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22844_ (.A0(\design_top.MEM[40][8] ),
    .A1(\design_top.MEM[41][8] ),
    .A2(\design_top.MEM[42][8] ),
    .A3(\design_top.MEM[43][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22845_ (.A0(\design_top.MEM[44][8] ),
    .A1(\design_top.MEM[45][8] ),
    .A2(\design_top.MEM[46][8] ),
    .A3(\design_top.MEM[47][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22846_ (.A0(_03444_),
    .A1(_03445_),
    .A2(_03446_),
    .A3(_03447_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22847_ (.A0(\design_top.MEM[48][8] ),
    .A1(\design_top.MEM[49][8] ),
    .A2(\design_top.MEM[50][8] ),
    .A3(\design_top.MEM[51][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22848_ (.A0(\design_top.MEM[52][8] ),
    .A1(\design_top.MEM[53][8] ),
    .A2(\design_top.MEM[54][8] ),
    .A3(\design_top.MEM[55][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22849_ (.A0(\design_top.MEM[56][8] ),
    .A1(\design_top.MEM[57][8] ),
    .A2(\design_top.MEM[58][8] ),
    .A3(\design_top.MEM[59][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22850_ (.A0(\design_top.MEM[60][8] ),
    .A1(\design_top.MEM[61][8] ),
    .A2(\design_top.MEM[62][8] ),
    .A3(\design_top.MEM[63][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22851_ (.A0(_03449_),
    .A1(_03450_),
    .A2(_03451_),
    .A3(_03452_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22852_ (.A0(_03438_),
    .A1(_03443_),
    .A2(_03448_),
    .A3(_03453_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22853_ (.A0(\design_top.MEM[0][7] ),
    .A1(\design_top.MEM[1][7] ),
    .A2(\design_top.MEM[2][7] ),
    .A3(\design_top.MEM[3][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22854_ (.A0(\design_top.MEM[4][7] ),
    .A1(\design_top.MEM[5][7] ),
    .A2(\design_top.MEM[6][7] ),
    .A3(\design_top.MEM[7][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22855_ (.A0(\design_top.MEM[8][7] ),
    .A1(\design_top.MEM[9][7] ),
    .A2(\design_top.MEM[10][7] ),
    .A3(\design_top.MEM[11][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22856_ (.A0(\design_top.MEM[12][7] ),
    .A1(\design_top.MEM[13][7] ),
    .A2(\design_top.MEM[14][7] ),
    .A3(\design_top.MEM[15][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22857_ (.A0(_03414_),
    .A1(_03415_),
    .A2(_03416_),
    .A3(_03417_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22858_ (.A0(\design_top.MEM[16][7] ),
    .A1(\design_top.MEM[17][7] ),
    .A2(\design_top.MEM[18][7] ),
    .A3(\design_top.MEM[19][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22859_ (.A0(\design_top.MEM[20][7] ),
    .A1(\design_top.MEM[21][7] ),
    .A2(\design_top.MEM[22][7] ),
    .A3(\design_top.MEM[23][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22860_ (.A0(\design_top.MEM[24][7] ),
    .A1(\design_top.MEM[25][7] ),
    .A2(\design_top.MEM[26][7] ),
    .A3(\design_top.MEM[27][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22861_ (.A0(\design_top.MEM[28][7] ),
    .A1(\design_top.MEM[29][7] ),
    .A2(\design_top.MEM[30][7] ),
    .A3(\design_top.MEM[31][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22862_ (.A0(_03419_),
    .A1(_03420_),
    .A2(_03421_),
    .A3(_03422_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22863_ (.A0(\design_top.MEM[32][7] ),
    .A1(\design_top.MEM[33][7] ),
    .A2(\design_top.MEM[34][7] ),
    .A3(\design_top.MEM[35][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22864_ (.A0(\design_top.MEM[36][7] ),
    .A1(\design_top.MEM[37][7] ),
    .A2(\design_top.MEM[38][7] ),
    .A3(\design_top.MEM[39][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22865_ (.A0(\design_top.MEM[40][7] ),
    .A1(\design_top.MEM[41][7] ),
    .A2(\design_top.MEM[42][7] ),
    .A3(\design_top.MEM[43][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22866_ (.A0(\design_top.MEM[44][7] ),
    .A1(\design_top.MEM[45][7] ),
    .A2(\design_top.MEM[46][7] ),
    .A3(\design_top.MEM[47][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22867_ (.A0(_03424_),
    .A1(_03425_),
    .A2(_03426_),
    .A3(_03427_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22868_ (.A0(\design_top.MEM[48][7] ),
    .A1(\design_top.MEM[49][7] ),
    .A2(\design_top.MEM[50][7] ),
    .A3(\design_top.MEM[51][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22869_ (.A0(\design_top.MEM[52][7] ),
    .A1(\design_top.MEM[53][7] ),
    .A2(\design_top.MEM[54][7] ),
    .A3(\design_top.MEM[55][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22870_ (.A0(\design_top.MEM[56][7] ),
    .A1(\design_top.MEM[57][7] ),
    .A2(\design_top.MEM[58][7] ),
    .A3(\design_top.MEM[59][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22871_ (.A0(\design_top.MEM[60][7] ),
    .A1(\design_top.MEM[61][7] ),
    .A2(\design_top.MEM[62][7] ),
    .A3(\design_top.MEM[63][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22872_ (.A0(_03429_),
    .A1(_03430_),
    .A2(_03431_),
    .A3(_03432_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22873_ (.A0(_03418_),
    .A1(_03423_),
    .A2(_03428_),
    .A3(_03433_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22874_ (.A0(\design_top.MEM[0][6] ),
    .A1(\design_top.MEM[1][6] ),
    .A2(\design_top.MEM[2][6] ),
    .A3(\design_top.MEM[3][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22875_ (.A0(\design_top.MEM[4][6] ),
    .A1(\design_top.MEM[5][6] ),
    .A2(\design_top.MEM[6][6] ),
    .A3(\design_top.MEM[7][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22876_ (.A0(\design_top.MEM[8][6] ),
    .A1(\design_top.MEM[9][6] ),
    .A2(\design_top.MEM[10][6] ),
    .A3(\design_top.MEM[11][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22877_ (.A0(\design_top.MEM[12][6] ),
    .A1(\design_top.MEM[13][6] ),
    .A2(\design_top.MEM[14][6] ),
    .A3(\design_top.MEM[15][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22878_ (.A0(_03394_),
    .A1(_03395_),
    .A2(_03396_),
    .A3(_03397_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22879_ (.A0(\design_top.MEM[16][6] ),
    .A1(\design_top.MEM[17][6] ),
    .A2(\design_top.MEM[18][6] ),
    .A3(\design_top.MEM[19][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22880_ (.A0(\design_top.MEM[20][6] ),
    .A1(\design_top.MEM[21][6] ),
    .A2(\design_top.MEM[22][6] ),
    .A3(\design_top.MEM[23][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22881_ (.A0(\design_top.MEM[24][6] ),
    .A1(\design_top.MEM[25][6] ),
    .A2(\design_top.MEM[26][6] ),
    .A3(\design_top.MEM[27][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22882_ (.A0(\design_top.MEM[28][6] ),
    .A1(\design_top.MEM[29][6] ),
    .A2(\design_top.MEM[30][6] ),
    .A3(\design_top.MEM[31][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22883_ (.A0(_03399_),
    .A1(_03400_),
    .A2(_03401_),
    .A3(_03402_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22884_ (.A0(\design_top.MEM[32][6] ),
    .A1(\design_top.MEM[33][6] ),
    .A2(\design_top.MEM[34][6] ),
    .A3(\design_top.MEM[35][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22885_ (.A0(\design_top.MEM[36][6] ),
    .A1(\design_top.MEM[37][6] ),
    .A2(\design_top.MEM[38][6] ),
    .A3(\design_top.MEM[39][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22886_ (.A0(\design_top.MEM[40][6] ),
    .A1(\design_top.MEM[41][6] ),
    .A2(\design_top.MEM[42][6] ),
    .A3(\design_top.MEM[43][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22887_ (.A0(\design_top.MEM[44][6] ),
    .A1(\design_top.MEM[45][6] ),
    .A2(\design_top.MEM[46][6] ),
    .A3(\design_top.MEM[47][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22888_ (.A0(_03404_),
    .A1(_03405_),
    .A2(_03406_),
    .A3(_03407_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22889_ (.A0(\design_top.MEM[48][6] ),
    .A1(\design_top.MEM[49][6] ),
    .A2(\design_top.MEM[50][6] ),
    .A3(\design_top.MEM[51][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22890_ (.A0(\design_top.MEM[52][6] ),
    .A1(\design_top.MEM[53][6] ),
    .A2(\design_top.MEM[54][6] ),
    .A3(\design_top.MEM[55][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22891_ (.A0(\design_top.MEM[56][6] ),
    .A1(\design_top.MEM[57][6] ),
    .A2(\design_top.MEM[58][6] ),
    .A3(\design_top.MEM[59][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22892_ (.A0(\design_top.MEM[60][6] ),
    .A1(\design_top.MEM[61][6] ),
    .A2(\design_top.MEM[62][6] ),
    .A3(\design_top.MEM[63][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22893_ (.A0(_03409_),
    .A1(_03410_),
    .A2(_03411_),
    .A3(_03412_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22894_ (.A0(_03398_),
    .A1(_03403_),
    .A2(_03408_),
    .A3(_03413_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22895_ (.A0(\design_top.MEM[0][5] ),
    .A1(\design_top.MEM[1][5] ),
    .A2(\design_top.MEM[2][5] ),
    .A3(\design_top.MEM[3][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22896_ (.A0(\design_top.MEM[4][5] ),
    .A1(\design_top.MEM[5][5] ),
    .A2(\design_top.MEM[6][5] ),
    .A3(\design_top.MEM[7][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22897_ (.A0(\design_top.MEM[8][5] ),
    .A1(\design_top.MEM[9][5] ),
    .A2(\design_top.MEM[10][5] ),
    .A3(\design_top.MEM[11][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22898_ (.A0(\design_top.MEM[12][5] ),
    .A1(\design_top.MEM[13][5] ),
    .A2(\design_top.MEM[14][5] ),
    .A3(\design_top.MEM[15][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22899_ (.A0(_03374_),
    .A1(_03375_),
    .A2(_03376_),
    .A3(_03377_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22900_ (.A0(\design_top.MEM[16][5] ),
    .A1(\design_top.MEM[17][5] ),
    .A2(\design_top.MEM[18][5] ),
    .A3(\design_top.MEM[19][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22901_ (.A0(\design_top.MEM[20][5] ),
    .A1(\design_top.MEM[21][5] ),
    .A2(\design_top.MEM[22][5] ),
    .A3(\design_top.MEM[23][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22902_ (.A0(\design_top.MEM[24][5] ),
    .A1(\design_top.MEM[25][5] ),
    .A2(\design_top.MEM[26][5] ),
    .A3(\design_top.MEM[27][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22903_ (.A0(\design_top.MEM[28][5] ),
    .A1(\design_top.MEM[29][5] ),
    .A2(\design_top.MEM[30][5] ),
    .A3(\design_top.MEM[31][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22904_ (.A0(_03379_),
    .A1(_03380_),
    .A2(_03381_),
    .A3(_03382_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22905_ (.A0(\design_top.MEM[32][5] ),
    .A1(\design_top.MEM[33][5] ),
    .A2(\design_top.MEM[34][5] ),
    .A3(\design_top.MEM[35][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22906_ (.A0(\design_top.MEM[36][5] ),
    .A1(\design_top.MEM[37][5] ),
    .A2(\design_top.MEM[38][5] ),
    .A3(\design_top.MEM[39][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22907_ (.A0(\design_top.MEM[40][5] ),
    .A1(\design_top.MEM[41][5] ),
    .A2(\design_top.MEM[42][5] ),
    .A3(\design_top.MEM[43][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22908_ (.A0(\design_top.MEM[44][5] ),
    .A1(\design_top.MEM[45][5] ),
    .A2(\design_top.MEM[46][5] ),
    .A3(\design_top.MEM[47][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22909_ (.A0(_03384_),
    .A1(_03385_),
    .A2(_03386_),
    .A3(_03387_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22910_ (.A0(\design_top.MEM[48][5] ),
    .A1(\design_top.MEM[49][5] ),
    .A2(\design_top.MEM[50][5] ),
    .A3(\design_top.MEM[51][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22911_ (.A0(\design_top.MEM[52][5] ),
    .A1(\design_top.MEM[53][5] ),
    .A2(\design_top.MEM[54][5] ),
    .A3(\design_top.MEM[55][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22912_ (.A0(\design_top.MEM[56][5] ),
    .A1(\design_top.MEM[57][5] ),
    .A2(\design_top.MEM[58][5] ),
    .A3(\design_top.MEM[59][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22913_ (.A0(\design_top.MEM[60][5] ),
    .A1(\design_top.MEM[61][5] ),
    .A2(\design_top.MEM[62][5] ),
    .A3(\design_top.MEM[63][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22914_ (.A0(_03389_),
    .A1(_03390_),
    .A2(_03391_),
    .A3(_03392_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22915_ (.A0(_03378_),
    .A1(_03383_),
    .A2(_03388_),
    .A3(_03393_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22916_ (.A0(\design_top.MEM[0][4] ),
    .A1(\design_top.MEM[1][4] ),
    .A2(\design_top.MEM[2][4] ),
    .A3(\design_top.MEM[3][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22917_ (.A0(\design_top.MEM[4][4] ),
    .A1(\design_top.MEM[5][4] ),
    .A2(\design_top.MEM[6][4] ),
    .A3(\design_top.MEM[7][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22918_ (.A0(\design_top.MEM[8][4] ),
    .A1(\design_top.MEM[9][4] ),
    .A2(\design_top.MEM[10][4] ),
    .A3(\design_top.MEM[11][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22919_ (.A0(\design_top.MEM[12][4] ),
    .A1(\design_top.MEM[13][4] ),
    .A2(\design_top.MEM[14][4] ),
    .A3(\design_top.MEM[15][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22920_ (.A0(_03354_),
    .A1(_03355_),
    .A2(_03356_),
    .A3(_03357_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22921_ (.A0(\design_top.MEM[16][4] ),
    .A1(\design_top.MEM[17][4] ),
    .A2(\design_top.MEM[18][4] ),
    .A3(\design_top.MEM[19][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22922_ (.A0(\design_top.MEM[20][4] ),
    .A1(\design_top.MEM[21][4] ),
    .A2(\design_top.MEM[22][4] ),
    .A3(\design_top.MEM[23][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22923_ (.A0(\design_top.MEM[24][4] ),
    .A1(\design_top.MEM[25][4] ),
    .A2(\design_top.MEM[26][4] ),
    .A3(\design_top.MEM[27][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22924_ (.A0(\design_top.MEM[28][4] ),
    .A1(\design_top.MEM[29][4] ),
    .A2(\design_top.MEM[30][4] ),
    .A3(\design_top.MEM[31][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22925_ (.A0(_03359_),
    .A1(_03360_),
    .A2(_03361_),
    .A3(_03362_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22926_ (.A0(\design_top.MEM[32][4] ),
    .A1(\design_top.MEM[33][4] ),
    .A2(\design_top.MEM[34][4] ),
    .A3(\design_top.MEM[35][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22927_ (.A0(\design_top.MEM[36][4] ),
    .A1(\design_top.MEM[37][4] ),
    .A2(\design_top.MEM[38][4] ),
    .A3(\design_top.MEM[39][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22928_ (.A0(\design_top.MEM[40][4] ),
    .A1(\design_top.MEM[41][4] ),
    .A2(\design_top.MEM[42][4] ),
    .A3(\design_top.MEM[43][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22929_ (.A0(\design_top.MEM[44][4] ),
    .A1(\design_top.MEM[45][4] ),
    .A2(\design_top.MEM[46][4] ),
    .A3(\design_top.MEM[47][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22930_ (.A0(_03364_),
    .A1(_03365_),
    .A2(_03366_),
    .A3(_03367_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22931_ (.A0(\design_top.MEM[48][4] ),
    .A1(\design_top.MEM[49][4] ),
    .A2(\design_top.MEM[50][4] ),
    .A3(\design_top.MEM[51][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22932_ (.A0(\design_top.MEM[52][4] ),
    .A1(\design_top.MEM[53][4] ),
    .A2(\design_top.MEM[54][4] ),
    .A3(\design_top.MEM[55][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22933_ (.A0(\design_top.MEM[56][4] ),
    .A1(\design_top.MEM[57][4] ),
    .A2(\design_top.MEM[58][4] ),
    .A3(\design_top.MEM[59][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22934_ (.A0(\design_top.MEM[60][4] ),
    .A1(\design_top.MEM[61][4] ),
    .A2(\design_top.MEM[62][4] ),
    .A3(\design_top.MEM[63][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22935_ (.A0(_03369_),
    .A1(_03370_),
    .A2(_03371_),
    .A3(_03372_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22936_ (.A0(_03358_),
    .A1(_03363_),
    .A2(_03368_),
    .A3(_03373_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22937_ (.A0(\design_top.MEM[0][3] ),
    .A1(\design_top.MEM[1][3] ),
    .A2(\design_top.MEM[2][3] ),
    .A3(\design_top.MEM[3][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22938_ (.A0(\design_top.MEM[4][3] ),
    .A1(\design_top.MEM[5][3] ),
    .A2(\design_top.MEM[6][3] ),
    .A3(\design_top.MEM[7][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22939_ (.A0(\design_top.MEM[8][3] ),
    .A1(\design_top.MEM[9][3] ),
    .A2(\design_top.MEM[10][3] ),
    .A3(\design_top.MEM[11][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22940_ (.A0(\design_top.MEM[12][3] ),
    .A1(\design_top.MEM[13][3] ),
    .A2(\design_top.MEM[14][3] ),
    .A3(\design_top.MEM[15][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22941_ (.A0(_03334_),
    .A1(_03335_),
    .A2(_03336_),
    .A3(_03337_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22942_ (.A0(\design_top.MEM[16][3] ),
    .A1(\design_top.MEM[17][3] ),
    .A2(\design_top.MEM[18][3] ),
    .A3(\design_top.MEM[19][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22943_ (.A0(\design_top.MEM[20][3] ),
    .A1(\design_top.MEM[21][3] ),
    .A2(\design_top.MEM[22][3] ),
    .A3(\design_top.MEM[23][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22944_ (.A0(\design_top.MEM[24][3] ),
    .A1(\design_top.MEM[25][3] ),
    .A2(\design_top.MEM[26][3] ),
    .A3(\design_top.MEM[27][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22945_ (.A0(\design_top.MEM[28][3] ),
    .A1(\design_top.MEM[29][3] ),
    .A2(\design_top.MEM[30][3] ),
    .A3(\design_top.MEM[31][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22946_ (.A0(_03339_),
    .A1(_03340_),
    .A2(_03341_),
    .A3(_03342_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22947_ (.A0(\design_top.MEM[32][3] ),
    .A1(\design_top.MEM[33][3] ),
    .A2(\design_top.MEM[34][3] ),
    .A3(\design_top.MEM[35][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22948_ (.A0(\design_top.MEM[36][3] ),
    .A1(\design_top.MEM[37][3] ),
    .A2(\design_top.MEM[38][3] ),
    .A3(\design_top.MEM[39][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22949_ (.A0(\design_top.MEM[40][3] ),
    .A1(\design_top.MEM[41][3] ),
    .A2(\design_top.MEM[42][3] ),
    .A3(\design_top.MEM[43][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22950_ (.A0(\design_top.MEM[44][3] ),
    .A1(\design_top.MEM[45][3] ),
    .A2(\design_top.MEM[46][3] ),
    .A3(\design_top.MEM[47][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22951_ (.A0(_03344_),
    .A1(_03345_),
    .A2(_03346_),
    .A3(_03347_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22952_ (.A0(\design_top.MEM[48][3] ),
    .A1(\design_top.MEM[49][3] ),
    .A2(\design_top.MEM[50][3] ),
    .A3(\design_top.MEM[51][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22953_ (.A0(\design_top.MEM[52][3] ),
    .A1(\design_top.MEM[53][3] ),
    .A2(\design_top.MEM[54][3] ),
    .A3(\design_top.MEM[55][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22954_ (.A0(\design_top.MEM[56][3] ),
    .A1(\design_top.MEM[57][3] ),
    .A2(\design_top.MEM[58][3] ),
    .A3(\design_top.MEM[59][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22955_ (.A0(\design_top.MEM[60][3] ),
    .A1(\design_top.MEM[61][3] ),
    .A2(\design_top.MEM[62][3] ),
    .A3(\design_top.MEM[63][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22956_ (.A0(_03349_),
    .A1(_03350_),
    .A2(_03351_),
    .A3(_03352_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22957_ (.A0(_03338_),
    .A1(_03343_),
    .A2(_03348_),
    .A3(_03353_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22958_ (.A0(\design_top.MEM[0][2] ),
    .A1(\design_top.MEM[1][2] ),
    .A2(\design_top.MEM[2][2] ),
    .A3(\design_top.MEM[3][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22959_ (.A0(\design_top.MEM[4][2] ),
    .A1(\design_top.MEM[5][2] ),
    .A2(\design_top.MEM[6][2] ),
    .A3(\design_top.MEM[7][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22960_ (.A0(\design_top.MEM[8][2] ),
    .A1(\design_top.MEM[9][2] ),
    .A2(\design_top.MEM[10][2] ),
    .A3(\design_top.MEM[11][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22961_ (.A0(\design_top.MEM[12][2] ),
    .A1(\design_top.MEM[13][2] ),
    .A2(\design_top.MEM[14][2] ),
    .A3(\design_top.MEM[15][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22962_ (.A0(_03314_),
    .A1(_03315_),
    .A2(_03316_),
    .A3(_03317_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22963_ (.A0(\design_top.MEM[16][2] ),
    .A1(\design_top.MEM[17][2] ),
    .A2(\design_top.MEM[18][2] ),
    .A3(\design_top.MEM[19][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22964_ (.A0(\design_top.MEM[20][2] ),
    .A1(\design_top.MEM[21][2] ),
    .A2(\design_top.MEM[22][2] ),
    .A3(\design_top.MEM[23][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22965_ (.A0(\design_top.MEM[24][2] ),
    .A1(\design_top.MEM[25][2] ),
    .A2(\design_top.MEM[26][2] ),
    .A3(\design_top.MEM[27][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22966_ (.A0(\design_top.MEM[28][2] ),
    .A1(\design_top.MEM[29][2] ),
    .A2(\design_top.MEM[30][2] ),
    .A3(\design_top.MEM[31][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22967_ (.A0(_03319_),
    .A1(_03320_),
    .A2(_03321_),
    .A3(_03322_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22968_ (.A0(\design_top.MEM[32][2] ),
    .A1(\design_top.MEM[33][2] ),
    .A2(\design_top.MEM[34][2] ),
    .A3(\design_top.MEM[35][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22969_ (.A0(\design_top.MEM[36][2] ),
    .A1(\design_top.MEM[37][2] ),
    .A2(\design_top.MEM[38][2] ),
    .A3(\design_top.MEM[39][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22970_ (.A0(\design_top.MEM[40][2] ),
    .A1(\design_top.MEM[41][2] ),
    .A2(\design_top.MEM[42][2] ),
    .A3(\design_top.MEM[43][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22971_ (.A0(\design_top.MEM[44][2] ),
    .A1(\design_top.MEM[45][2] ),
    .A2(\design_top.MEM[46][2] ),
    .A3(\design_top.MEM[47][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22972_ (.A0(_03324_),
    .A1(_03325_),
    .A2(_03326_),
    .A3(_03327_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22973_ (.A0(\design_top.MEM[48][2] ),
    .A1(\design_top.MEM[49][2] ),
    .A2(\design_top.MEM[50][2] ),
    .A3(\design_top.MEM[51][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22974_ (.A0(\design_top.MEM[52][2] ),
    .A1(\design_top.MEM[53][2] ),
    .A2(\design_top.MEM[54][2] ),
    .A3(\design_top.MEM[55][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22975_ (.A0(\design_top.MEM[56][2] ),
    .A1(\design_top.MEM[57][2] ),
    .A2(\design_top.MEM[58][2] ),
    .A3(\design_top.MEM[59][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22976_ (.A0(\design_top.MEM[60][2] ),
    .A1(\design_top.MEM[61][2] ),
    .A2(\design_top.MEM[62][2] ),
    .A3(\design_top.MEM[63][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22977_ (.A0(_03329_),
    .A1(_03330_),
    .A2(_03331_),
    .A3(_03332_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22978_ (.A0(_03318_),
    .A1(_03323_),
    .A2(_03328_),
    .A3(_03333_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22979_ (.A0(\design_top.MEM[0][1] ),
    .A1(\design_top.MEM[1][1] ),
    .A2(\design_top.MEM[2][1] ),
    .A3(\design_top.MEM[3][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22980_ (.A0(\design_top.MEM[4][1] ),
    .A1(\design_top.MEM[5][1] ),
    .A2(\design_top.MEM[6][1] ),
    .A3(\design_top.MEM[7][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22981_ (.A0(\design_top.MEM[8][1] ),
    .A1(\design_top.MEM[9][1] ),
    .A2(\design_top.MEM[10][1] ),
    .A3(\design_top.MEM[11][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22982_ (.A0(\design_top.MEM[12][1] ),
    .A1(\design_top.MEM[13][1] ),
    .A2(\design_top.MEM[14][1] ),
    .A3(\design_top.MEM[15][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22983_ (.A0(_03294_),
    .A1(_03295_),
    .A2(_03296_),
    .A3(_03297_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22984_ (.A0(\design_top.MEM[16][1] ),
    .A1(\design_top.MEM[17][1] ),
    .A2(\design_top.MEM[18][1] ),
    .A3(\design_top.MEM[19][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22985_ (.A0(\design_top.MEM[20][1] ),
    .A1(\design_top.MEM[21][1] ),
    .A2(\design_top.MEM[22][1] ),
    .A3(\design_top.MEM[23][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22986_ (.A0(\design_top.MEM[24][1] ),
    .A1(\design_top.MEM[25][1] ),
    .A2(\design_top.MEM[26][1] ),
    .A3(\design_top.MEM[27][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22987_ (.A0(\design_top.MEM[28][1] ),
    .A1(\design_top.MEM[29][1] ),
    .A2(\design_top.MEM[30][1] ),
    .A3(\design_top.MEM[31][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22988_ (.A0(_03299_),
    .A1(_03300_),
    .A2(_03301_),
    .A3(_03302_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22989_ (.A0(\design_top.MEM[32][1] ),
    .A1(\design_top.MEM[33][1] ),
    .A2(\design_top.MEM[34][1] ),
    .A3(\design_top.MEM[35][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22990_ (.A0(\design_top.MEM[36][1] ),
    .A1(\design_top.MEM[37][1] ),
    .A2(\design_top.MEM[38][1] ),
    .A3(\design_top.MEM[39][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22991_ (.A0(\design_top.MEM[40][1] ),
    .A1(\design_top.MEM[41][1] ),
    .A2(\design_top.MEM[42][1] ),
    .A3(\design_top.MEM[43][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22992_ (.A0(\design_top.MEM[44][1] ),
    .A1(\design_top.MEM[45][1] ),
    .A2(\design_top.MEM[46][1] ),
    .A3(\design_top.MEM[47][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22993_ (.A0(_03304_),
    .A1(_03305_),
    .A2(_03306_),
    .A3(_03307_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22994_ (.A0(\design_top.MEM[48][1] ),
    .A1(\design_top.MEM[49][1] ),
    .A2(\design_top.MEM[50][1] ),
    .A3(\design_top.MEM[51][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22995_ (.A0(\design_top.MEM[52][1] ),
    .A1(\design_top.MEM[53][1] ),
    .A2(\design_top.MEM[54][1] ),
    .A3(\design_top.MEM[55][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22996_ (.A0(\design_top.MEM[56][1] ),
    .A1(\design_top.MEM[57][1] ),
    .A2(\design_top.MEM[58][1] ),
    .A3(\design_top.MEM[59][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22997_ (.A0(\design_top.MEM[60][1] ),
    .A1(\design_top.MEM[61][1] ),
    .A2(\design_top.MEM[62][1] ),
    .A3(\design_top.MEM[63][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22998_ (.A0(_03309_),
    .A1(_03310_),
    .A2(_03311_),
    .A3(_03312_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _22999_ (.A0(_03298_),
    .A1(_03303_),
    .A2(_03308_),
    .A3(_03313_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23000_ (.A0(\design_top.MEM[0][0] ),
    .A1(\design_top.MEM[1][0] ),
    .A2(\design_top.MEM[2][0] ),
    .A3(\design_top.MEM[3][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23001_ (.A0(\design_top.MEM[4][0] ),
    .A1(\design_top.MEM[5][0] ),
    .A2(\design_top.MEM[6][0] ),
    .A3(\design_top.MEM[7][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23002_ (.A0(\design_top.MEM[8][0] ),
    .A1(\design_top.MEM[9][0] ),
    .A2(\design_top.MEM[10][0] ),
    .A3(\design_top.MEM[11][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23003_ (.A0(\design_top.MEM[12][0] ),
    .A1(\design_top.MEM[13][0] ),
    .A2(\design_top.MEM[14][0] ),
    .A3(\design_top.MEM[15][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23004_ (.A0(_03274_),
    .A1(_03275_),
    .A2(_03276_),
    .A3(_03277_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23005_ (.A0(\design_top.MEM[16][0] ),
    .A1(\design_top.MEM[17][0] ),
    .A2(\design_top.MEM[18][0] ),
    .A3(\design_top.MEM[19][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23006_ (.A0(\design_top.MEM[20][0] ),
    .A1(\design_top.MEM[21][0] ),
    .A2(\design_top.MEM[22][0] ),
    .A3(\design_top.MEM[23][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23007_ (.A0(\design_top.MEM[24][0] ),
    .A1(\design_top.MEM[25][0] ),
    .A2(\design_top.MEM[26][0] ),
    .A3(\design_top.MEM[27][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23008_ (.A0(\design_top.MEM[28][0] ),
    .A1(\design_top.MEM[29][0] ),
    .A2(\design_top.MEM[30][0] ),
    .A3(\design_top.MEM[31][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23009_ (.A0(_03279_),
    .A1(_03280_),
    .A2(_03281_),
    .A3(_03282_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23010_ (.A0(\design_top.MEM[32][0] ),
    .A1(\design_top.MEM[33][0] ),
    .A2(\design_top.MEM[34][0] ),
    .A3(\design_top.MEM[35][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23011_ (.A0(\design_top.MEM[36][0] ),
    .A1(\design_top.MEM[37][0] ),
    .A2(\design_top.MEM[38][0] ),
    .A3(\design_top.MEM[39][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23012_ (.A0(\design_top.MEM[40][0] ),
    .A1(\design_top.MEM[41][0] ),
    .A2(\design_top.MEM[42][0] ),
    .A3(\design_top.MEM[43][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23013_ (.A0(\design_top.MEM[44][0] ),
    .A1(\design_top.MEM[45][0] ),
    .A2(\design_top.MEM[46][0] ),
    .A3(\design_top.MEM[47][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23014_ (.A0(_03284_),
    .A1(_03285_),
    .A2(_03286_),
    .A3(_03287_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23015_ (.A0(\design_top.MEM[48][0] ),
    .A1(\design_top.MEM[49][0] ),
    .A2(\design_top.MEM[50][0] ),
    .A3(\design_top.MEM[51][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23016_ (.A0(\design_top.MEM[52][0] ),
    .A1(\design_top.MEM[53][0] ),
    .A2(\design_top.MEM[54][0] ),
    .A3(\design_top.MEM[55][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23017_ (.A0(\design_top.MEM[56][0] ),
    .A1(\design_top.MEM[57][0] ),
    .A2(\design_top.MEM[58][0] ),
    .A3(\design_top.MEM[59][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23018_ (.A0(\design_top.MEM[60][0] ),
    .A1(\design_top.MEM[61][0] ),
    .A2(\design_top.MEM[62][0] ),
    .A3(\design_top.MEM[63][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23019_ (.A0(_03289_),
    .A1(_03290_),
    .A2(_03291_),
    .A3(_03292_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _23020_ (.A0(_03278_),
    .A1(_03283_),
    .A2(_03288_),
    .A3(_03293_),
    .S0(\design_top.IADDR[6] ),
    .S1(\design_top.IADDR[7] ),
    .X(_00141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23021_ (.D(_00141_),
    .Q(\design_top.ROMFF[0] ),
    .CLK(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23022_ (.D(_00152_),
    .Q(\design_top.ROMFF[1] ),
    .CLK(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23023_ (.D(_00163_),
    .Q(\design_top.ROMFF[2] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23024_ (.D(_00166_),
    .Q(\design_top.ROMFF[3] ),
    .CLK(clknet_leaf_408_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23025_ (.D(_00167_),
    .Q(\design_top.ROMFF[4] ),
    .CLK(clknet_leaf_408_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23026_ (.D(_00168_),
    .Q(\design_top.ROMFF[5] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23027_ (.D(_00169_),
    .Q(\design_top.ROMFF[6] ),
    .CLK(clknet_leaf_402_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23028_ (.D(_00170_),
    .Q(\design_top.ROMFF[7] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23029_ (.D(_00171_),
    .Q(\design_top.ROMFF[8] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23030_ (.D(_00172_),
    .Q(\design_top.ROMFF[9] ),
    .CLK(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23031_ (.D(_00142_),
    .Q(\design_top.ROMFF[10] ),
    .CLK(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23032_ (.D(_00143_),
    .Q(\design_top.ROMFF[11] ),
    .CLK(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23033_ (.D(_00144_),
    .Q(\design_top.ROMFF[12] ),
    .CLK(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23034_ (.D(_00145_),
    .Q(\design_top.ROMFF[13] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23035_ (.D(_00146_),
    .Q(\design_top.ROMFF[14] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23036_ (.D(_00147_),
    .Q(\design_top.ROMFF[15] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23037_ (.D(_00148_),
    .Q(\design_top.ROMFF[16] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23038_ (.D(_00149_),
    .Q(\design_top.ROMFF[17] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23039_ (.D(_00150_),
    .Q(\design_top.ROMFF[18] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23040_ (.D(_00151_),
    .Q(\design_top.ROMFF[19] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23041_ (.D(_00153_),
    .Q(\design_top.ROMFF[20] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23042_ (.D(_00154_),
    .Q(\design_top.ROMFF[21] ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23043_ (.D(_00155_),
    .Q(\design_top.ROMFF[22] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23044_ (.D(_00156_),
    .Q(\design_top.ROMFF[23] ),
    .CLK(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23045_ (.D(_00157_),
    .Q(\design_top.ROMFF[24] ),
    .CLK(clknet_leaf_386_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23046_ (.D(_00158_),
    .Q(\design_top.ROMFF[25] ),
    .CLK(clknet_leaf_386_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23047_ (.D(_00159_),
    .Q(\design_top.ROMFF[26] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23048_ (.D(_00160_),
    .Q(\design_top.ROMFF[27] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23049_ (.D(_00161_),
    .Q(\design_top.ROMFF[28] ),
    .CLK(clknet_leaf_384_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23050_ (.D(_00162_),
    .Q(\design_top.ROMFF[29] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23051_ (.D(_00164_),
    .Q(\design_top.ROMFF[30] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23052_ (.D(_00165_),
    .Q(\design_top.ROMFF[31] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23053_ (.D(_00046_),
    .Q(\design_top.core0.XRES ),
    .CLK(clknet_leaf_291_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23054_ (.D(io_in[1]),
    .Q(\design_top.uart0.UART_RXDFF[0] ),
    .CLK(clknet_leaf_351_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23055_ (.D(\design_top.uart0.UART_RXDFF[0] ),
    .Q(\design_top.uart0.UART_RXDFF[1] ),
    .CLK(clknet_leaf_351_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23056_ (.D(\design_top.uart0.UART_RXDFF[1] ),
    .Q(\design_top.uart0.UART_RXDFF[2] ),
    .CLK(clknet_leaf_350_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23057_ (.D(\design_top.XRES_reg ),
    .Q(\design_top.XRES ),
    .CLK(clknet_leaf_337_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23058_ (.D(io_in[0]),
    .Q(\design_top.XRES_reg ),
    .CLK(clknet_leaf_337_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23059_ (.D(\design_top.HLT ),
    .Q(\design_top.HLT2 ),
    .CLK(clknet_leaf_311_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23060_ (.D(\design_top.DADDR[2] ),
    .Q(\design_top.XADDR[2] ),
    .CLK(clknet_leaf_368_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23061_ (.D(\design_top.DADDR[3] ),
    .Q(\design_top.XADDR[3] ),
    .CLK(clknet_leaf_374_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23062_ (.D(\design_top.DADDR[31] ),
    .Q(\design_top.XADDR[31] ),
    .CLK(clknet_leaf_375_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23063_ (.D(_00109_),
    .Q(\design_top.RAMFF[0] ),
    .CLK(clknet_leaf_408_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23064_ (.D(_00120_),
    .Q(\design_top.RAMFF[1] ),
    .CLK(clknet_leaf_433_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23065_ (.D(_00131_),
    .Q(\design_top.RAMFF[2] ),
    .CLK(clknet_leaf_402_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23066_ (.D(_00134_),
    .Q(\design_top.RAMFF[3] ),
    .CLK(clknet_leaf_367_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23067_ (.D(_00135_),
    .Q(\design_top.RAMFF[4] ),
    .CLK(clknet_leaf_369_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23068_ (.D(_00136_),
    .Q(\design_top.RAMFF[5] ),
    .CLK(clknet_leaf_367_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23069_ (.D(_00137_),
    .Q(\design_top.RAMFF[6] ),
    .CLK(clknet_leaf_366_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23070_ (.D(_00138_),
    .Q(\design_top.RAMFF[7] ),
    .CLK(clknet_leaf_366_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23071_ (.D(_00139_),
    .Q(\design_top.RAMFF[8] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23072_ (.D(_00140_),
    .Q(\design_top.RAMFF[9] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23073_ (.D(_00110_),
    .Q(\design_top.RAMFF[10] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23074_ (.D(_00111_),
    .Q(\design_top.RAMFF[11] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23075_ (.D(_00112_),
    .Q(\design_top.RAMFF[12] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23076_ (.D(_00113_),
    .Q(\design_top.RAMFF[13] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23077_ (.D(_00114_),
    .Q(\design_top.RAMFF[14] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23078_ (.D(_00115_),
    .Q(\design_top.RAMFF[15] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23079_ (.D(_00116_),
    .Q(\design_top.RAMFF[16] ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23080_ (.D(_00117_),
    .Q(\design_top.RAMFF[17] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23081_ (.D(_00118_),
    .Q(\design_top.RAMFF[18] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23082_ (.D(_00119_),
    .Q(\design_top.RAMFF[19] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23083_ (.D(_00121_),
    .Q(\design_top.RAMFF[20] ),
    .CLK(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23084_ (.D(_00122_),
    .Q(\design_top.RAMFF[21] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23085_ (.D(_00123_),
    .Q(\design_top.RAMFF[22] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23086_ (.D(_00124_),
    .Q(\design_top.RAMFF[23] ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23087_ (.D(_00125_),
    .Q(\design_top.RAMFF[24] ),
    .CLK(clknet_leaf_374_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23088_ (.D(_00126_),
    .Q(\design_top.RAMFF[25] ),
    .CLK(clknet_leaf_375_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23089_ (.D(_00127_),
    .Q(\design_top.RAMFF[26] ),
    .CLK(clknet_leaf_374_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23090_ (.D(_00128_),
    .Q(\design_top.RAMFF[27] ),
    .CLK(clknet_leaf_370_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23091_ (.D(_00129_),
    .Q(\design_top.RAMFF[28] ),
    .CLK(clknet_leaf_366_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23092_ (.D(_00130_),
    .Q(\design_top.RAMFF[29] ),
    .CLK(clknet_leaf_366_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23093_ (.D(_00132_),
    .Q(\design_top.RAMFF[30] ),
    .CLK(clknet_leaf_373_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23094_ (.D(_00133_),
    .Q(\design_top.RAMFF[31] ),
    .CLK(clknet_leaf_373_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23095_ (.D(_03972_),
    .Q(\design_top.uart0.UART_XFIFO[0] ),
    .CLK(clknet_leaf_368_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23096_ (.D(_03973_),
    .Q(\design_top.uart0.UART_XFIFO[1] ),
    .CLK(clknet_leaf_368_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23097_ (.D(_03974_),
    .Q(\design_top.uart0.UART_XFIFO[2] ),
    .CLK(clknet_leaf_368_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23098_ (.D(_03975_),
    .Q(\design_top.uart0.UART_XFIFO[3] ),
    .CLK(clknet_leaf_368_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23099_ (.D(_03976_),
    .Q(\design_top.uart0.UART_XFIFO[4] ),
    .CLK(clknet_leaf_368_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23100_ (.D(_03977_),
    .Q(\design_top.uart0.UART_XFIFO[5] ),
    .CLK(clknet_leaf_368_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23101_ (.D(_03978_),
    .Q(\design_top.uart0.UART_XFIFO[6] ),
    .CLK(clknet_leaf_347_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23102_ (.D(_03979_),
    .Q(\design_top.uart0.UART_XFIFO[7] ),
    .CLK(clknet_leaf_368_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23103_ (.D(_03980_),
    .Q(\design_top.uart0.UART_XREQ ),
    .CLK(clknet_leaf_345_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23104_ (.D(_03981_),
    .Q(\design_top.uart0.UART_RACK ),
    .CLK(clknet_leaf_352_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23105_ (.D(_03982_),
    .Q(\design_top.core0.REG2[9][0] ),
    .CLK(clknet_leaf_296_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23106_ (.D(_03983_),
    .Q(\design_top.core0.REG2[9][1] ),
    .CLK(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23107_ (.D(_03984_),
    .Q(\design_top.core0.REG2[9][2] ),
    .CLK(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23108_ (.D(_03985_),
    .Q(\design_top.core0.REG2[9][3] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23109_ (.D(_03986_),
    .Q(\design_top.core0.REG2[9][4] ),
    .CLK(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23110_ (.D(_03987_),
    .Q(\design_top.core0.REG2[9][5] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23111_ (.D(_03988_),
    .Q(\design_top.core0.REG2[9][6] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23112_ (.D(_03989_),
    .Q(\design_top.core0.REG2[9][7] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23113_ (.D(_03990_),
    .Q(\design_top.core0.REG2[9][8] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23114_ (.D(_03991_),
    .Q(\design_top.core0.REG2[9][9] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23115_ (.D(_03992_),
    .Q(\design_top.core0.REG2[9][10] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23116_ (.D(_03993_),
    .Q(\design_top.core0.REG2[9][11] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23117_ (.D(_03994_),
    .Q(\design_top.core0.REG2[9][12] ),
    .CLK(clknet_leaf_301_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23118_ (.D(_03995_),
    .Q(\design_top.core0.REG2[9][13] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23119_ (.D(_03996_),
    .Q(\design_top.core0.REG2[9][14] ),
    .CLK(clknet_leaf_301_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23120_ (.D(_03997_),
    .Q(\design_top.core0.REG2[9][15] ),
    .CLK(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23121_ (.D(_03998_),
    .Q(\design_top.core0.REG2[9][16] ),
    .CLK(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23122_ (.D(_03999_),
    .Q(\design_top.core0.REG2[9][17] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23123_ (.D(_04000_),
    .Q(\design_top.core0.REG2[9][18] ),
    .CLK(clknet_leaf_295_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23124_ (.D(_04001_),
    .Q(\design_top.core0.REG2[9][19] ),
    .CLK(clknet_leaf_295_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23125_ (.D(_04002_),
    .Q(\design_top.core0.REG2[9][20] ),
    .CLK(clknet_leaf_295_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23126_ (.D(_04003_),
    .Q(\design_top.core0.REG2[9][21] ),
    .CLK(clknet_leaf_269_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23127_ (.D(_04004_),
    .Q(\design_top.core0.REG2[9][22] ),
    .CLK(clknet_leaf_277_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23128_ (.D(_04005_),
    .Q(\design_top.core0.REG2[9][23] ),
    .CLK(clknet_leaf_278_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23129_ (.D(_04006_),
    .Q(\design_top.core0.REG2[9][24] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23130_ (.D(_04007_),
    .Q(\design_top.core0.REG2[9][25] ),
    .CLK(clknet_leaf_278_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23131_ (.D(_04008_),
    .Q(\design_top.core0.REG2[9][26] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23132_ (.D(_04009_),
    .Q(\design_top.core0.REG2[9][27] ),
    .CLK(clknet_leaf_271_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23133_ (.D(_04010_),
    .Q(\design_top.core0.REG2[9][28] ),
    .CLK(clknet_leaf_260_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23134_ (.D(_04011_),
    .Q(\design_top.core0.REG2[9][29] ),
    .CLK(clknet_leaf_271_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23135_ (.D(_04012_),
    .Q(\design_top.core0.REG2[9][30] ),
    .CLK(clknet_leaf_260_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23136_ (.D(_04013_),
    .Q(\design_top.core0.REG2[9][31] ),
    .CLK(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23137_ (.D(_04014_),
    .Q(\design_top.core0.NXPC[0] ),
    .CLK(clknet_leaf_307_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23138_ (.D(_04015_),
    .Q(\design_top.core0.NXPC[1] ),
    .CLK(clknet_leaf_319_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23139_ (.D(_04016_),
    .Q(\design_top.core0.NXPC[2] ),
    .CLK(clknet_leaf_316_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23140_ (.D(_04017_),
    .Q(\design_top.core0.NXPC[3] ),
    .CLK(clknet_leaf_316_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23141_ (.D(_04018_),
    .Q(\design_top.core0.NXPC[4] ),
    .CLK(clknet_leaf_316_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23142_ (.D(_04019_),
    .Q(\design_top.core0.NXPC[5] ),
    .CLK(clknet_leaf_312_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23143_ (.D(_04020_),
    .Q(\design_top.core0.NXPC[6] ),
    .CLK(clknet_leaf_312_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23144_ (.D(_04021_),
    .Q(\design_top.core0.NXPC[7] ),
    .CLK(clknet_leaf_309_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23145_ (.D(_04022_),
    .Q(\design_top.core0.NXPC[8] ),
    .CLK(clknet_leaf_309_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23146_ (.D(_04023_),
    .Q(\design_top.core0.NXPC[9] ),
    .CLK(clknet_leaf_305_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23147_ (.D(_04024_),
    .Q(\design_top.core0.NXPC[10] ),
    .CLK(clknet_leaf_305_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23148_ (.D(_04025_),
    .Q(\design_top.core0.NXPC[11] ),
    .CLK(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23149_ (.D(_04026_),
    .Q(\design_top.core0.NXPC[12] ),
    .CLK(clknet_leaf_291_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23150_ (.D(_04027_),
    .Q(\design_top.core0.NXPC[13] ),
    .CLK(clknet_leaf_291_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23151_ (.D(_04028_),
    .Q(\design_top.core0.NXPC[14] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23152_ (.D(_04029_),
    .Q(\design_top.core0.NXPC[15] ),
    .CLK(clknet_leaf_288_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23153_ (.D(_04030_),
    .Q(\design_top.core0.NXPC[16] ),
    .CLK(clknet_leaf_288_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23154_ (.D(_04031_),
    .Q(\design_top.core0.NXPC[17] ),
    .CLK(clknet_leaf_288_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23155_ (.D(_04032_),
    .Q(\design_top.core0.NXPC[18] ),
    .CLK(clknet_leaf_289_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23156_ (.D(_04033_),
    .Q(\design_top.core0.NXPC[19] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23157_ (.D(_04034_),
    .Q(\design_top.core0.NXPC[20] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23158_ (.D(_04035_),
    .Q(\design_top.core0.NXPC[21] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23159_ (.D(_04036_),
    .Q(\design_top.core0.NXPC[22] ),
    .CLK(clknet_leaf_284_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23160_ (.D(_04037_),
    .Q(\design_top.core0.NXPC[23] ),
    .CLK(clknet_leaf_283_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23161_ (.D(_04038_),
    .Q(\design_top.core0.NXPC[24] ),
    .CLK(clknet_leaf_282_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23162_ (.D(_04039_),
    .Q(\design_top.core0.NXPC[25] ),
    .CLK(clknet_leaf_282_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23163_ (.D(_04040_),
    .Q(\design_top.core0.NXPC[26] ),
    .CLK(clknet_leaf_282_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23164_ (.D(_04041_),
    .Q(\design_top.core0.NXPC[27] ),
    .CLK(clknet_leaf_331_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23165_ (.D(_04042_),
    .Q(\design_top.core0.NXPC[28] ),
    .CLK(clknet_leaf_330_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23166_ (.D(_04043_),
    .Q(\design_top.core0.NXPC[29] ),
    .CLK(clknet_leaf_330_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23167_ (.D(_04044_),
    .Q(\design_top.core0.NXPC[30] ),
    .CLK(clknet_leaf_330_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23168_ (.D(_04045_),
    .Q(\design_top.core0.NXPC[31] ),
    .CLK(clknet_leaf_329_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23169_ (.D(_04046_),
    .Q(\design_top.core0.PC[0] ),
    .CLK(clknet_leaf_319_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23170_ (.D(_04047_),
    .Q(\design_top.core0.PC[1] ),
    .CLK(clknet_leaf_319_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23171_ (.D(_04048_),
    .Q(\design_top.core0.PC[2] ),
    .CLK(clknet_leaf_316_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23172_ (.D(_04049_),
    .Q(\design_top.core0.PC[3] ),
    .CLK(clknet_leaf_316_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23173_ (.D(_04050_),
    .Q(\design_top.core0.PC[4] ),
    .CLK(clknet_leaf_316_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23174_ (.D(_04051_),
    .Q(\design_top.core0.PC[5] ),
    .CLK(clknet_leaf_312_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23175_ (.D(_04052_),
    .Q(\design_top.core0.PC[6] ),
    .CLK(clknet_leaf_312_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23176_ (.D(_04053_),
    .Q(\design_top.core0.PC[7] ),
    .CLK(clknet_leaf_310_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23177_ (.D(_04054_),
    .Q(\design_top.core0.PC[8] ),
    .CLK(clknet_leaf_307_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23178_ (.D(_04055_),
    .Q(\design_top.core0.PC[9] ),
    .CLK(clknet_leaf_305_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23179_ (.D(_04056_),
    .Q(\design_top.core0.PC[10] ),
    .CLK(clknet_leaf_305_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23180_ (.D(_04057_),
    .Q(\design_top.core0.PC[11] ),
    .CLK(clknet_leaf_291_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23181_ (.D(_04058_),
    .Q(\design_top.core0.PC[12] ),
    .CLK(clknet_leaf_291_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23182_ (.D(_04059_),
    .Q(\design_top.core0.PC[13] ),
    .CLK(clknet_leaf_291_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23183_ (.D(_04060_),
    .Q(\design_top.core0.PC[14] ),
    .CLK(clknet_leaf_290_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23184_ (.D(_04061_),
    .Q(\design_top.core0.PC[15] ),
    .CLK(clknet_leaf_288_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23185_ (.D(_04062_),
    .Q(\design_top.core0.PC[16] ),
    .CLK(clknet_leaf_290_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23186_ (.D(_04063_),
    .Q(\design_top.core0.PC[17] ),
    .CLK(clknet_leaf_288_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23187_ (.D(_04064_),
    .Q(\design_top.core0.PC[18] ),
    .CLK(clknet_leaf_289_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23188_ (.D(_04065_),
    .Q(\design_top.core0.PC[19] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23189_ (.D(_04066_),
    .Q(\design_top.core0.PC[20] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23190_ (.D(_04067_),
    .Q(\design_top.core0.PC[21] ),
    .CLK(clknet_leaf_284_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23191_ (.D(_04068_),
    .Q(\design_top.core0.PC[22] ),
    .CLK(clknet_leaf_283_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23192_ (.D(_04069_),
    .Q(\design_top.core0.PC[23] ),
    .CLK(clknet_leaf_283_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23193_ (.D(_04070_),
    .Q(\design_top.core0.PC[24] ),
    .CLK(clknet_leaf_282_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23194_ (.D(_04071_),
    .Q(\design_top.core0.PC[25] ),
    .CLK(clknet_leaf_283_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23195_ (.D(_04072_),
    .Q(\design_top.core0.PC[26] ),
    .CLK(clknet_leaf_331_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23196_ (.D(_04073_),
    .Q(\design_top.core0.PC[27] ),
    .CLK(clknet_leaf_331_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23197_ (.D(_04074_),
    .Q(\design_top.core0.PC[28] ),
    .CLK(clknet_leaf_331_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23198_ (.D(_04075_),
    .Q(\design_top.core0.PC[29] ),
    .CLK(clknet_leaf_330_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23199_ (.D(_04076_),
    .Q(\design_top.core0.PC[30] ),
    .CLK(clknet_leaf_330_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23200_ (.D(_04077_),
    .Q(\design_top.core0.PC[31] ),
    .CLK(clknet_leaf_329_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23201_ (.D(_04078_),
    .Q(\design_top.uart0.UART_RFIFO[0] ),
    .CLK(clknet_leaf_352_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23202_ (.D(_04079_),
    .Q(\design_top.uart0.UART_RFIFO[1] ),
    .CLK(clknet_leaf_350_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23203_ (.D(_04080_),
    .Q(\design_top.uart0.UART_RFIFO[2] ),
    .CLK(clknet_leaf_352_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23204_ (.D(_04081_),
    .Q(\design_top.uart0.UART_RFIFO[3] ),
    .CLK(clknet_leaf_348_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23205_ (.D(_04082_),
    .Q(\design_top.uart0.UART_RFIFO[4] ),
    .CLK(clknet_leaf_348_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23206_ (.D(_04083_),
    .Q(\design_top.uart0.UART_RFIFO[5] ),
    .CLK(clknet_leaf_348_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23207_ (.D(_04084_),
    .Q(\design_top.uart0.UART_RFIFO[6] ),
    .CLK(clknet_leaf_348_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23208_ (.D(_04085_),
    .Q(\design_top.uart0.UART_RFIFO[7] ),
    .CLK(clknet_leaf_349_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23209_ (.D(_04086_),
    .Q(\design_top.uart0.UART_RREQ ),
    .CLK(clknet_leaf_352_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23210_ (.D(_04087_),
    .Q(\design_top.uart0.UART_XACK ),
    .CLK(clknet_leaf_345_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23211_ (.D(_04088_),
    .Q(\design_top.ROMFF2[0] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23212_ (.D(_04089_),
    .Q(\design_top.ROMFF2[1] ),
    .CLK(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23213_ (.D(_04090_),
    .Q(\design_top.ROMFF2[2] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23214_ (.D(_04091_),
    .Q(\design_top.ROMFF2[3] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23215_ (.D(_04092_),
    .Q(\design_top.ROMFF2[4] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23216_ (.D(_04093_),
    .Q(\design_top.ROMFF2[5] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23217_ (.D(_04094_),
    .Q(\design_top.ROMFF2[6] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23218_ (.D(_04095_),
    .Q(\design_top.ROMFF2[7] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23219_ (.D(_04096_),
    .Q(\design_top.ROMFF2[8] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23220_ (.D(_04097_),
    .Q(\design_top.ROMFF2[9] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23221_ (.D(_04098_),
    .Q(\design_top.ROMFF2[10] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23222_ (.D(_04099_),
    .Q(\design_top.ROMFF2[11] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23223_ (.D(_04100_),
    .Q(\design_top.ROMFF2[12] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23224_ (.D(_04101_),
    .Q(\design_top.ROMFF2[13] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23225_ (.D(_04102_),
    .Q(\design_top.ROMFF2[14] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23226_ (.D(_04103_),
    .Q(\design_top.ROMFF2[15] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23227_ (.D(_04104_),
    .Q(\design_top.ROMFF2[16] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23228_ (.D(_04105_),
    .Q(\design_top.ROMFF2[17] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23229_ (.D(_04106_),
    .Q(\design_top.ROMFF2[18] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23230_ (.D(_04107_),
    .Q(\design_top.ROMFF2[19] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23231_ (.D(_04108_),
    .Q(\design_top.ROMFF2[20] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23232_ (.D(_04109_),
    .Q(\design_top.ROMFF2[21] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23233_ (.D(_04110_),
    .Q(\design_top.ROMFF2[22] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23234_ (.D(_04111_),
    .Q(\design_top.ROMFF2[23] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23235_ (.D(_04112_),
    .Q(\design_top.ROMFF2[24] ),
    .CLK(clknet_leaf_315_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23236_ (.D(_04113_),
    .Q(\design_top.ROMFF2[25] ),
    .CLK(clknet_leaf_314_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23237_ (.D(_04114_),
    .Q(\design_top.ROMFF2[26] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23238_ (.D(_04115_),
    .Q(\design_top.ROMFF2[27] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23239_ (.D(_04116_),
    .Q(\design_top.ROMFF2[28] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23240_ (.D(_04117_),
    .Q(\design_top.ROMFF2[29] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23241_ (.D(_04118_),
    .Q(\design_top.ROMFF2[30] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23242_ (.D(_04119_),
    .Q(\design_top.ROMFF2[31] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23243_ (.D(_04120_),
    .Q(io_out[8]),
    .CLK(clknet_leaf_347_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23244_ (.D(_04121_),
    .Q(io_out[9]),
    .CLK(clknet_leaf_347_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23245_ (.D(_04122_),
    .Q(io_out[10]),
    .CLK(clknet_leaf_347_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23246_ (.D(_04123_),
    .Q(io_out[11]),
    .CLK(clknet_leaf_353_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23247_ (.D(_04124_),
    .Q(\design_top.LEDFF[4] ),
    .CLK(clknet_leaf_347_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23248_ (.D(_04125_),
    .Q(\design_top.LEDFF[5] ),
    .CLK(clknet_leaf_353_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23249_ (.D(_04126_),
    .Q(\design_top.LEDFF[6] ),
    .CLK(clknet_leaf_347_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23250_ (.D(_04127_),
    .Q(\design_top.LEDFF[7] ),
    .CLK(clknet_leaf_347_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23251_ (.D(_04128_),
    .Q(\design_top.LEDFF[8] ),
    .CLK(clknet_leaf_347_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23252_ (.D(_04129_),
    .Q(\design_top.LEDFF[9] ),
    .CLK(clknet_leaf_347_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23253_ (.D(_04130_),
    .Q(\design_top.LEDFF[10] ),
    .CLK(clknet_leaf_347_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23254_ (.D(_04131_),
    .Q(\design_top.LEDFF[11] ),
    .CLK(clknet_leaf_347_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23255_ (.D(_04132_),
    .Q(\design_top.LEDFF[12] ),
    .CLK(clknet_leaf_347_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23256_ (.D(_04133_),
    .Q(\design_top.LEDFF[13] ),
    .CLK(clknet_leaf_347_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23257_ (.D(_04134_),
    .Q(\design_top.LEDFF[14] ),
    .CLK(clknet_leaf_347_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23258_ (.D(_04135_),
    .Q(\design_top.LEDFF[15] ),
    .CLK(clknet_leaf_346_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23259_ (.D(_04136_),
    .Q(io_out[15]),
    .CLK(clknet_leaf_373_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23260_ (.D(_04137_),
    .Q(\design_top.GPIOFF[1] ),
    .CLK(clknet_leaf_373_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23261_ (.D(_04138_),
    .Q(\design_top.GPIOFF[2] ),
    .CLK(clknet_leaf_372_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23262_ (.D(_04139_),
    .Q(\design_top.GPIOFF[3] ),
    .CLK(clknet_leaf_372_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23263_ (.D(_04140_),
    .Q(\design_top.GPIOFF[4] ),
    .CLK(clknet_leaf_372_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23264_ (.D(_04141_),
    .Q(\design_top.GPIOFF[5] ),
    .CLK(clknet_leaf_370_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23265_ (.D(_04142_),
    .Q(\design_top.GPIOFF[6] ),
    .CLK(clknet_leaf_370_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23266_ (.D(_04143_),
    .Q(\design_top.GPIOFF[7] ),
    .CLK(clknet_leaf_373_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23267_ (.D(_04144_),
    .Q(\design_top.GPIOFF[8] ),
    .CLK(clknet_leaf_373_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23268_ (.D(_04145_),
    .Q(\design_top.GPIOFF[9] ),
    .CLK(clknet_leaf_373_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23269_ (.D(_04146_),
    .Q(\design_top.GPIOFF[10] ),
    .CLK(clknet_leaf_370_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23270_ (.D(_04147_),
    .Q(\design_top.GPIOFF[11] ),
    .CLK(clknet_leaf_370_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23271_ (.D(_04148_),
    .Q(\design_top.GPIOFF[12] ),
    .CLK(clknet_leaf_370_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23272_ (.D(_04149_),
    .Q(\design_top.GPIOFF[13] ),
    .CLK(clknet_leaf_370_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23273_ (.D(_04150_),
    .Q(\design_top.GPIOFF[14] ),
    .CLK(clknet_leaf_370_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23274_ (.D(_04151_),
    .Q(\design_top.GPIOFF[15] ),
    .CLK(clknet_leaf_369_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23275_ (.D(_04152_),
    .Q(\design_top.MEM[55][0] ),
    .CLK(clknet_leaf_402_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23276_ (.D(_04153_),
    .Q(\design_top.MEM[55][1] ),
    .CLK(clknet_leaf_405_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23277_ (.D(_04154_),
    .Q(\design_top.MEM[55][2] ),
    .CLK(clknet_leaf_405_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23278_ (.D(_04155_),
    .Q(\design_top.MEM[55][3] ),
    .CLK(clknet_leaf_429_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23279_ (.D(_04156_),
    .Q(\design_top.MEM[55][4] ),
    .CLK(clknet_leaf_429_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23280_ (.D(_04157_),
    .Q(\design_top.MEM[55][5] ),
    .CLK(clknet_leaf_423_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23281_ (.D(_04158_),
    .Q(\design_top.MEM[55][6] ),
    .CLK(clknet_leaf_422_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23282_ (.D(_04159_),
    .Q(\design_top.MEM[55][7] ),
    .CLK(clknet_leaf_422_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23283_ (.D(_04160_),
    .Q(\design_top.MEM[56][0] ),
    .CLK(clknet_leaf_407_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23284_ (.D(_04161_),
    .Q(\design_top.MEM[56][1] ),
    .CLK(clknet_leaf_406_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23285_ (.D(_04162_),
    .Q(\design_top.MEM[56][2] ),
    .CLK(clknet_leaf_407_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23286_ (.D(_04163_),
    .Q(\design_top.MEM[56][3] ),
    .CLK(clknet_leaf_412_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23287_ (.D(_04164_),
    .Q(\design_top.MEM[56][4] ),
    .CLK(clknet_leaf_420_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23288_ (.D(_04165_),
    .Q(\design_top.MEM[56][5] ),
    .CLK(clknet_leaf_419_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23289_ (.D(_04166_),
    .Q(\design_top.MEM[56][6] ),
    .CLK(clknet_leaf_420_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23290_ (.D(_04167_),
    .Q(\design_top.MEM[56][7] ),
    .CLK(clknet_leaf_418_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23291_ (.D(_04168_),
    .Q(\design_top.MEM[57][0] ),
    .CLK(clknet_leaf_408_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23292_ (.D(_04169_),
    .Q(\design_top.MEM[57][1] ),
    .CLK(clknet_leaf_407_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23293_ (.D(_04170_),
    .Q(\design_top.MEM[57][2] ),
    .CLK(clknet_leaf_407_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23294_ (.D(_04171_),
    .Q(\design_top.MEM[57][3] ),
    .CLK(clknet_leaf_413_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23295_ (.D(_04172_),
    .Q(\design_top.MEM[57][4] ),
    .CLK(clknet_leaf_414_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23296_ (.D(_04173_),
    .Q(\design_top.MEM[57][5] ),
    .CLK(clknet_leaf_418_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23297_ (.D(_04174_),
    .Q(\design_top.MEM[57][6] ),
    .CLK(clknet_leaf_418_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23298_ (.D(_04175_),
    .Q(\design_top.MEM[57][7] ),
    .CLK(clknet_leaf_418_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23299_ (.D(_04176_),
    .Q(\design_top.MEM[58][0] ),
    .CLK(clknet_leaf_408_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23300_ (.D(_04177_),
    .Q(\design_top.MEM[58][1] ),
    .CLK(clknet_leaf_412_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23301_ (.D(_04178_),
    .Q(\design_top.MEM[58][2] ),
    .CLK(clknet_leaf_408_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23302_ (.D(_04179_),
    .Q(\design_top.MEM[58][3] ),
    .CLK(clknet_leaf_413_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23303_ (.D(_04180_),
    .Q(\design_top.MEM[58][4] ),
    .CLK(clknet_leaf_420_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23304_ (.D(_04181_),
    .Q(\design_top.MEM[58][5] ),
    .CLK(clknet_leaf_419_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23305_ (.D(_04182_),
    .Q(\design_top.MEM[58][6] ),
    .CLK(clknet_leaf_420_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23306_ (.D(_04183_),
    .Q(\design_top.MEM[58][7] ),
    .CLK(clknet_leaf_419_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23307_ (.D(_04184_),
    .Q(\design_top.MEM[59][0] ),
    .CLK(clknet_leaf_408_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23308_ (.D(_04185_),
    .Q(\design_top.MEM[59][1] ),
    .CLK(clknet_leaf_406_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23309_ (.D(_04186_),
    .Q(\design_top.MEM[59][2] ),
    .CLK(clknet_leaf_407_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23310_ (.D(_04187_),
    .Q(\design_top.MEM[59][3] ),
    .CLK(clknet_leaf_412_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23311_ (.D(_04188_),
    .Q(\design_top.MEM[59][4] ),
    .CLK(clknet_leaf_420_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23312_ (.D(_04189_),
    .Q(\design_top.MEM[59][5] ),
    .CLK(clknet_leaf_419_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23313_ (.D(_04190_),
    .Q(\design_top.MEM[59][6] ),
    .CLK(clknet_leaf_420_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23314_ (.D(_04191_),
    .Q(\design_top.MEM[59][7] ),
    .CLK(clknet_leaf_420_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23315_ (.D(_04192_),
    .Q(\design_top.MEM[5][0] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23316_ (.D(_04193_),
    .Q(\design_top.MEM[5][1] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23317_ (.D(_04194_),
    .Q(\design_top.MEM[5][2] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23318_ (.D(_04195_),
    .Q(\design_top.MEM[5][3] ),
    .CLK(clknet_leaf_400_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23319_ (.D(_04196_),
    .Q(\design_top.MEM[5][4] ),
    .CLK(clknet_leaf_402_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23320_ (.D(_04197_),
    .Q(\design_top.MEM[5][5] ),
    .CLK(clknet_leaf_401_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23321_ (.D(_04198_),
    .Q(\design_top.MEM[5][6] ),
    .CLK(clknet_leaf_400_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23322_ (.D(_04199_),
    .Q(\design_top.MEM[5][7] ),
    .CLK(clknet_leaf_401_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23323_ (.D(_04200_),
    .Q(\design_top.MEM[60][0] ),
    .CLK(clknet_leaf_408_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23324_ (.D(_04201_),
    .Q(\design_top.MEM[60][1] ),
    .CLK(clknet_leaf_406_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23325_ (.D(_04202_),
    .Q(\design_top.MEM[60][2] ),
    .CLK(clknet_leaf_407_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23326_ (.D(_04203_),
    .Q(\design_top.MEM[60][3] ),
    .CLK(clknet_leaf_421_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23327_ (.D(_04204_),
    .Q(\design_top.MEM[60][4] ),
    .CLK(clknet_leaf_421_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23328_ (.D(_04205_),
    .Q(\design_top.MEM[60][5] ),
    .CLK(clknet_leaf_419_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23329_ (.D(_04206_),
    .Q(\design_top.MEM[60][6] ),
    .CLK(clknet_leaf_422_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23330_ (.D(_04207_),
    .Q(\design_top.MEM[60][7] ),
    .CLK(clknet_leaf_423_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23331_ (.D(_04208_),
    .Q(\design_top.core0.REG1[15][0] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23332_ (.D(_04209_),
    .Q(\design_top.core0.REG1[15][1] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23333_ (.D(_04210_),
    .Q(\design_top.core0.REG1[15][2] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23334_ (.D(_04211_),
    .Q(\design_top.core0.REG1[15][3] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23335_ (.D(_04212_),
    .Q(\design_top.core0.REG1[15][4] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23336_ (.D(_04213_),
    .Q(\design_top.core0.REG1[15][5] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23337_ (.D(_04214_),
    .Q(\design_top.core0.REG1[15][6] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23338_ (.D(_04215_),
    .Q(\design_top.core0.REG1[15][7] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23339_ (.D(_04216_),
    .Q(\design_top.core0.REG1[15][8] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23340_ (.D(_04217_),
    .Q(\design_top.core0.REG1[15][9] ),
    .CLK(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23341_ (.D(_04218_),
    .Q(\design_top.core0.REG1[15][10] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23342_ (.D(_04219_),
    .Q(\design_top.core0.REG1[15][11] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23343_ (.D(_04220_),
    .Q(\design_top.core0.REG1[15][12] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23344_ (.D(_04221_),
    .Q(\design_top.core0.REG1[15][13] ),
    .CLK(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23345_ (.D(_04222_),
    .Q(\design_top.core0.REG1[15][14] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23346_ (.D(_04223_),
    .Q(\design_top.core0.REG1[15][15] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23347_ (.D(_04224_),
    .Q(\design_top.core0.REG1[15][16] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23348_ (.D(_04225_),
    .Q(\design_top.core0.REG1[15][17] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23349_ (.D(_04226_),
    .Q(\design_top.core0.REG1[15][18] ),
    .CLK(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23350_ (.D(_04227_),
    .Q(\design_top.core0.REG1[15][19] ),
    .CLK(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23351_ (.D(_04228_),
    .Q(\design_top.core0.REG1[15][20] ),
    .CLK(clknet_leaf_263_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23352_ (.D(_04229_),
    .Q(\design_top.core0.REG1[15][21] ),
    .CLK(clknet_leaf_263_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23353_ (.D(_04230_),
    .Q(\design_top.core0.REG1[15][22] ),
    .CLK(clknet_leaf_264_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23354_ (.D(_04231_),
    .Q(\design_top.core0.REG1[15][23] ),
    .CLK(clknet_leaf_260_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23355_ (.D(_04232_),
    .Q(\design_top.core0.REG1[15][24] ),
    .CLK(clknet_leaf_261_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23356_ (.D(_04233_),
    .Q(\design_top.core0.REG1[15][25] ),
    .CLK(clknet_leaf_260_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23357_ (.D(_04234_),
    .Q(\design_top.core0.REG1[15][26] ),
    .CLK(clknet_leaf_261_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23358_ (.D(_04235_),
    .Q(\design_top.core0.REG1[15][27] ),
    .CLK(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23359_ (.D(_04236_),
    .Q(\design_top.core0.REG1[15][28] ),
    .CLK(clknet_leaf_256_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23360_ (.D(_04237_),
    .Q(\design_top.core0.REG1[15][29] ),
    .CLK(clknet_leaf_259_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23361_ (.D(_04238_),
    .Q(\design_top.core0.REG1[15][30] ),
    .CLK(clknet_leaf_259_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23362_ (.D(_04239_),
    .Q(\design_top.core0.REG1[15][31] ),
    .CLK(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23363_ (.D(_04240_),
    .Q(\design_top.core0.REG1[1][0] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23364_ (.D(_04241_),
    .Q(\design_top.core0.REG1[1][1] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23365_ (.D(_04242_),
    .Q(\design_top.core0.REG1[1][2] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23366_ (.D(_04243_),
    .Q(\design_top.core0.REG1[1][3] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23367_ (.D(_04244_),
    .Q(\design_top.core0.REG1[1][4] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23368_ (.D(_04245_),
    .Q(\design_top.core0.REG1[1][5] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23369_ (.D(_04246_),
    .Q(\design_top.core0.REG1[1][6] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23370_ (.D(_04247_),
    .Q(\design_top.core0.REG1[1][7] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23371_ (.D(_04248_),
    .Q(\design_top.core0.REG1[1][8] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23372_ (.D(_04249_),
    .Q(\design_top.core0.REG1[1][9] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23373_ (.D(_04250_),
    .Q(\design_top.core0.REG1[1][10] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23374_ (.D(_04251_),
    .Q(\design_top.core0.REG1[1][11] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23375_ (.D(_04252_),
    .Q(\design_top.core0.REG1[1][12] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23376_ (.D(_04253_),
    .Q(\design_top.core0.REG1[1][13] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23377_ (.D(_04254_),
    .Q(\design_top.core0.REG1[1][14] ),
    .CLK(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23378_ (.D(_04255_),
    .Q(\design_top.core0.REG1[1][15] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23379_ (.D(_04256_),
    .Q(\design_top.core0.REG1[1][16] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23380_ (.D(_04257_),
    .Q(\design_top.core0.REG1[1][17] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23381_ (.D(_04258_),
    .Q(\design_top.core0.REG1[1][18] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23382_ (.D(_04259_),
    .Q(\design_top.core0.REG1[1][19] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23383_ (.D(_04260_),
    .Q(\design_top.core0.REG1[1][20] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23384_ (.D(_04261_),
    .Q(\design_top.core0.REG1[1][21] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23385_ (.D(_04262_),
    .Q(\design_top.core0.REG1[1][22] ),
    .CLK(clknet_leaf_245_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23386_ (.D(_04263_),
    .Q(\design_top.core0.REG1[1][23] ),
    .CLK(clknet_leaf_244_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23387_ (.D(_04264_),
    .Q(\design_top.core0.REG1[1][24] ),
    .CLK(clknet_leaf_245_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23388_ (.D(_04265_),
    .Q(\design_top.core0.REG1[1][25] ),
    .CLK(clknet_leaf_245_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23389_ (.D(_04266_),
    .Q(\design_top.core0.REG1[1][26] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23390_ (.D(_04267_),
    .Q(\design_top.core0.REG1[1][27] ),
    .CLK(clknet_leaf_251_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23391_ (.D(_04268_),
    .Q(\design_top.core0.REG1[1][28] ),
    .CLK(clknet_leaf_251_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23392_ (.D(_04269_),
    .Q(\design_top.core0.REG1[1][29] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23393_ (.D(_04270_),
    .Q(\design_top.core0.REG1[1][30] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23394_ (.D(_04271_),
    .Q(\design_top.core0.REG1[1][31] ),
    .CLK(clknet_leaf_251_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23395_ (.D(_04272_),
    .Q(\design_top.core0.REG1[2][0] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23396_ (.D(_04273_),
    .Q(\design_top.core0.REG1[2][1] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23397_ (.D(_04274_),
    .Q(\design_top.core0.REG1[2][2] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23398_ (.D(_04275_),
    .Q(\design_top.core0.REG1[2][3] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23399_ (.D(_04276_),
    .Q(\design_top.core0.REG1[2][4] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23400_ (.D(_04277_),
    .Q(\design_top.core0.REG1[2][5] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23401_ (.D(_04278_),
    .Q(\design_top.core0.REG1[2][6] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23402_ (.D(_04279_),
    .Q(\design_top.core0.REG1[2][7] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23403_ (.D(_04280_),
    .Q(\design_top.core0.REG1[2][8] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23404_ (.D(_04281_),
    .Q(\design_top.core0.REG1[2][9] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23405_ (.D(_04282_),
    .Q(\design_top.core0.REG1[2][10] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23406_ (.D(_04283_),
    .Q(\design_top.core0.REG1[2][11] ),
    .CLK(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23407_ (.D(_04284_),
    .Q(\design_top.core0.REG1[2][12] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23408_ (.D(_04285_),
    .Q(\design_top.core0.REG1[2][13] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23409_ (.D(_04286_),
    .Q(\design_top.core0.REG1[2][14] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23410_ (.D(_04287_),
    .Q(\design_top.core0.REG1[2][15] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23411_ (.D(_04288_),
    .Q(\design_top.core0.REG1[2][16] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23412_ (.D(_04289_),
    .Q(\design_top.core0.REG1[2][17] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23413_ (.D(_04290_),
    .Q(\design_top.core0.REG1[2][18] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23414_ (.D(_04291_),
    .Q(\design_top.core0.REG1[2][19] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23415_ (.D(_04292_),
    .Q(\design_top.core0.REG1[2][20] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23416_ (.D(_04293_),
    .Q(\design_top.core0.REG1[2][21] ),
    .CLK(clknet_leaf_244_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23417_ (.D(_04294_),
    .Q(\design_top.core0.REG1[2][22] ),
    .CLK(clknet_leaf_245_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23418_ (.D(_04295_),
    .Q(\design_top.core0.REG1[2][23] ),
    .CLK(clknet_leaf_245_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23419_ (.D(_04296_),
    .Q(\design_top.core0.REG1[2][24] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23420_ (.D(_04297_),
    .Q(\design_top.core0.REG1[2][25] ),
    .CLK(clknet_leaf_245_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23421_ (.D(_04298_),
    .Q(\design_top.core0.REG1[2][26] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23422_ (.D(_04299_),
    .Q(\design_top.core0.REG1[2][27] ),
    .CLK(clknet_leaf_250_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23423_ (.D(_04300_),
    .Q(\design_top.core0.REG1[2][28] ),
    .CLK(clknet_leaf_251_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23424_ (.D(_04301_),
    .Q(\design_top.core0.REG1[2][29] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23425_ (.D(_04302_),
    .Q(\design_top.core0.REG1[2][30] ),
    .CLK(clknet_leaf_251_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23426_ (.D(_04303_),
    .Q(\design_top.core0.REG1[2][31] ),
    .CLK(clknet_leaf_251_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23427_ (.D(_04304_),
    .Q(\design_top.core0.REG1[3][0] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23428_ (.D(_04305_),
    .Q(\design_top.core0.REG1[3][1] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23429_ (.D(_04306_),
    .Q(\design_top.core0.REG1[3][2] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23430_ (.D(_04307_),
    .Q(\design_top.core0.REG1[3][3] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23431_ (.D(_04308_),
    .Q(\design_top.core0.REG1[3][4] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23432_ (.D(_04309_),
    .Q(\design_top.core0.REG1[3][5] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23433_ (.D(_04310_),
    .Q(\design_top.core0.REG1[3][6] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23434_ (.D(_04311_),
    .Q(\design_top.core0.REG1[3][7] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23435_ (.D(_04312_),
    .Q(\design_top.core0.REG1[3][8] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23436_ (.D(_04313_),
    .Q(\design_top.core0.REG1[3][9] ),
    .CLK(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23437_ (.D(_04314_),
    .Q(\design_top.core0.REG1[3][10] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23438_ (.D(_04315_),
    .Q(\design_top.core0.REG1[3][11] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23439_ (.D(_04316_),
    .Q(\design_top.core0.REG1[3][12] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23440_ (.D(_04317_),
    .Q(\design_top.core0.REG1[3][13] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23441_ (.D(_04318_),
    .Q(\design_top.core0.REG1[3][14] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23442_ (.D(_04319_),
    .Q(\design_top.core0.REG1[3][15] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23443_ (.D(_04320_),
    .Q(\design_top.core0.REG1[3][16] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23444_ (.D(_04321_),
    .Q(\design_top.core0.REG1[3][17] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23445_ (.D(_04322_),
    .Q(\design_top.core0.REG1[3][18] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23446_ (.D(_04323_),
    .Q(\design_top.core0.REG1[3][19] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23447_ (.D(_04324_),
    .Q(\design_top.core0.REG1[3][20] ),
    .CLK(clknet_leaf_244_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23448_ (.D(_04325_),
    .Q(\design_top.core0.REG1[3][21] ),
    .CLK(clknet_leaf_244_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23449_ (.D(_04326_),
    .Q(\design_top.core0.REG1[3][22] ),
    .CLK(clknet_leaf_244_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23450_ (.D(_04327_),
    .Q(\design_top.core0.REG1[3][23] ),
    .CLK(clknet_leaf_244_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23451_ (.D(_04328_),
    .Q(\design_top.core0.REG1[3][24] ),
    .CLK(clknet_leaf_245_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23452_ (.D(_04329_),
    .Q(\design_top.core0.REG1[3][25] ),
    .CLK(clknet_leaf_245_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23453_ (.D(_04330_),
    .Q(\design_top.core0.REG1[3][26] ),
    .CLK(clknet_leaf_246_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23454_ (.D(_04331_),
    .Q(\design_top.core0.REG1[3][27] ),
    .CLK(clknet_leaf_250_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23455_ (.D(_04332_),
    .Q(\design_top.core0.REG1[3][28] ),
    .CLK(clknet_leaf_250_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23456_ (.D(_04333_),
    .Q(\design_top.core0.REG1[3][29] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23457_ (.D(_04334_),
    .Q(\design_top.core0.REG1[3][30] ),
    .CLK(clknet_leaf_249_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23458_ (.D(_04335_),
    .Q(\design_top.core0.REG1[3][31] ),
    .CLK(clknet_leaf_250_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23459_ (.D(_04336_),
    .Q(\design_top.core0.REG1[4][0] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23460_ (.D(_04337_),
    .Q(\design_top.core0.REG1[4][1] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23461_ (.D(_04338_),
    .Q(\design_top.core0.REG1[4][2] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23462_ (.D(_04339_),
    .Q(\design_top.core0.REG1[4][3] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23463_ (.D(_04340_),
    .Q(\design_top.core0.REG1[4][4] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23464_ (.D(_04341_),
    .Q(\design_top.core0.REG1[4][5] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23465_ (.D(_04342_),
    .Q(\design_top.core0.REG1[4][6] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23466_ (.D(_04343_),
    .Q(\design_top.core0.REG1[4][7] ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23467_ (.D(_04344_),
    .Q(\design_top.core0.REG1[4][8] ),
    .CLK(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23468_ (.D(_04345_),
    .Q(\design_top.core0.REG1[4][9] ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23469_ (.D(_04346_),
    .Q(\design_top.core0.REG1[4][10] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23470_ (.D(_04347_),
    .Q(\design_top.core0.REG1[4][11] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23471_ (.D(_04348_),
    .Q(\design_top.core0.REG1[4][12] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23472_ (.D(_04349_),
    .Q(\design_top.core0.REG1[4][13] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23473_ (.D(_04350_),
    .Q(\design_top.core0.REG1[4][14] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23474_ (.D(_04351_),
    .Q(\design_top.core0.REG1[4][15] ),
    .CLK(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23475_ (.D(_04352_),
    .Q(\design_top.core0.REG1[4][16] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23476_ (.D(_04353_),
    .Q(\design_top.core0.REG1[4][17] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23477_ (.D(_04354_),
    .Q(\design_top.core0.REG1[4][18] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23478_ (.D(_04355_),
    .Q(\design_top.core0.REG1[4][19] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23479_ (.D(_04356_),
    .Q(\design_top.core0.REG1[4][20] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23480_ (.D(_04357_),
    .Q(\design_top.core0.REG1[4][21] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23481_ (.D(_04358_),
    .Q(\design_top.core0.REG1[4][22] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23482_ (.D(_04359_),
    .Q(\design_top.core0.REG1[4][23] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23483_ (.D(_04360_),
    .Q(\design_top.core0.REG1[4][24] ),
    .CLK(clknet_leaf_247_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23484_ (.D(_04361_),
    .Q(\design_top.core0.REG1[4][25] ),
    .CLK(clknet_leaf_246_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23485_ (.D(_04362_),
    .Q(\design_top.core0.REG1[4][26] ),
    .CLK(clknet_leaf_247_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23486_ (.D(_04363_),
    .Q(\design_top.core0.REG1[4][27] ),
    .CLK(clknet_leaf_249_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23487_ (.D(_04364_),
    .Q(\design_top.core0.REG1[4][28] ),
    .CLK(clknet_leaf_248_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23488_ (.D(_04365_),
    .Q(\design_top.core0.REG1[4][29] ),
    .CLK(clknet_leaf_246_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23489_ (.D(_04366_),
    .Q(\design_top.core0.REG1[4][30] ),
    .CLK(clknet_leaf_248_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23490_ (.D(_04367_),
    .Q(\design_top.core0.REG1[4][31] ),
    .CLK(clknet_leaf_248_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23491_ (.D(_04368_),
    .Q(\design_top.core0.REG1[5][0] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23492_ (.D(_04369_),
    .Q(\design_top.core0.REG1[5][1] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23493_ (.D(_04370_),
    .Q(\design_top.core0.REG1[5][2] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23494_ (.D(_04371_),
    .Q(\design_top.core0.REG1[5][3] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23495_ (.D(_04372_),
    .Q(\design_top.core0.REG1[5][4] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23496_ (.D(_04373_),
    .Q(\design_top.core0.REG1[5][5] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23497_ (.D(_04374_),
    .Q(\design_top.core0.REG1[5][6] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23498_ (.D(_04375_),
    .Q(\design_top.core0.REG1[5][7] ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23499_ (.D(_04376_),
    .Q(\design_top.core0.REG1[5][8] ),
    .CLK(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23500_ (.D(_04377_),
    .Q(\design_top.core0.REG1[5][9] ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23501_ (.D(_04378_),
    .Q(\design_top.core0.REG1[5][10] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23502_ (.D(_04379_),
    .Q(\design_top.core0.REG1[5][11] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23503_ (.D(_04380_),
    .Q(\design_top.core0.REG1[5][12] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23504_ (.D(_04381_),
    .Q(\design_top.core0.REG1[5][13] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23505_ (.D(_04382_),
    .Q(\design_top.core0.REG1[5][14] ),
    .CLK(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23506_ (.D(_04383_),
    .Q(\design_top.core0.REG1[5][15] ),
    .CLK(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23507_ (.D(_04384_),
    .Q(\design_top.core0.REG1[5][16] ),
    .CLK(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23508_ (.D(_04385_),
    .Q(\design_top.core0.REG1[5][17] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23509_ (.D(_04386_),
    .Q(\design_top.core0.REG1[5][18] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23510_ (.D(_04387_),
    .Q(\design_top.core0.REG1[5][19] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23511_ (.D(_04388_),
    .Q(\design_top.core0.REG1[5][20] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23512_ (.D(_04389_),
    .Q(\design_top.core0.REG1[5][21] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23513_ (.D(_04390_),
    .Q(\design_top.core0.REG1[5][22] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23514_ (.D(_04391_),
    .Q(\design_top.core0.REG1[5][23] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23515_ (.D(_04392_),
    .Q(\design_top.core0.REG1[5][24] ),
    .CLK(clknet_leaf_247_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23516_ (.D(_04393_),
    .Q(\design_top.core0.REG1[5][25] ),
    .CLK(clknet_leaf_247_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23517_ (.D(_04394_),
    .Q(\design_top.core0.REG1[5][26] ),
    .CLK(clknet_leaf_247_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23518_ (.D(_04395_),
    .Q(\design_top.core0.REG1[5][27] ),
    .CLK(clknet_leaf_249_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23519_ (.D(_04396_),
    .Q(\design_top.core0.REG1[5][28] ),
    .CLK(clknet_leaf_248_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23520_ (.D(_04397_),
    .Q(\design_top.core0.REG1[5][29] ),
    .CLK(clknet_leaf_246_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23521_ (.D(_04398_),
    .Q(\design_top.core0.REG1[5][30] ),
    .CLK(clknet_leaf_248_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23522_ (.D(_04399_),
    .Q(\design_top.core0.REG1[5][31] ),
    .CLK(clknet_leaf_248_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23523_ (.D(_04400_),
    .Q(\design_top.MEM[61][0] ),
    .CLK(clknet_leaf_408_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23524_ (.D(_04401_),
    .Q(\design_top.MEM[61][1] ),
    .CLK(clknet_leaf_406_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23525_ (.D(_04402_),
    .Q(\design_top.MEM[61][2] ),
    .CLK(clknet_leaf_405_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23526_ (.D(_04403_),
    .Q(\design_top.MEM[61][3] ),
    .CLK(clknet_leaf_413_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23527_ (.D(_04404_),
    .Q(\design_top.MEM[61][4] ),
    .CLK(clknet_leaf_420_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23528_ (.D(_04405_),
    .Q(\design_top.MEM[61][5] ),
    .CLK(clknet_leaf_420_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23529_ (.D(_04406_),
    .Q(\design_top.MEM[61][6] ),
    .CLK(clknet_leaf_420_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23530_ (.D(_04407_),
    .Q(\design_top.MEM[61][7] ),
    .CLK(clknet_leaf_420_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23531_ (.D(_04408_),
    .Q(\design_top.core0.REG1[6][0] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23532_ (.D(_04409_),
    .Q(\design_top.core0.REG1[6][1] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23533_ (.D(_04410_),
    .Q(\design_top.core0.REG1[6][2] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23534_ (.D(_04411_),
    .Q(\design_top.core0.REG1[6][3] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23535_ (.D(_04412_),
    .Q(\design_top.core0.REG1[6][4] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23536_ (.D(_04413_),
    .Q(\design_top.core0.REG1[6][5] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23537_ (.D(_04414_),
    .Q(\design_top.core0.REG1[6][6] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23538_ (.D(_04415_),
    .Q(\design_top.core0.REG1[6][7] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23539_ (.D(_04416_),
    .Q(\design_top.core0.REG1[6][8] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23540_ (.D(_04417_),
    .Q(\design_top.core0.REG1[6][9] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23541_ (.D(_04418_),
    .Q(\design_top.core0.REG1[6][10] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23542_ (.D(_04419_),
    .Q(\design_top.core0.REG1[6][11] ),
    .CLK(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23543_ (.D(_04420_),
    .Q(\design_top.core0.REG1[6][12] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23544_ (.D(_04421_),
    .Q(\design_top.core0.REG1[6][13] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23545_ (.D(_04422_),
    .Q(\design_top.core0.REG1[6][14] ),
    .CLK(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23546_ (.D(_04423_),
    .Q(\design_top.core0.REG1[6][15] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23547_ (.D(_04424_),
    .Q(\design_top.core0.REG1[6][16] ),
    .CLK(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23548_ (.D(_04425_),
    .Q(\design_top.core0.REG1[6][17] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23549_ (.D(_04426_),
    .Q(\design_top.core0.REG1[6][18] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23550_ (.D(_04427_),
    .Q(\design_top.core0.REG1[6][19] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23551_ (.D(_04428_),
    .Q(\design_top.core0.REG1[6][20] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23552_ (.D(_04429_),
    .Q(\design_top.core0.REG1[6][21] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23553_ (.D(_04430_),
    .Q(\design_top.core0.REG1[6][22] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23554_ (.D(_04431_),
    .Q(\design_top.core0.REG1[6][23] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23555_ (.D(_04432_),
    .Q(\design_top.core0.REG1[6][24] ),
    .CLK(clknet_leaf_246_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23556_ (.D(_04433_),
    .Q(\design_top.core0.REG1[6][25] ),
    .CLK(clknet_leaf_247_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23557_ (.D(_04434_),
    .Q(\design_top.core0.REG1[6][26] ),
    .CLK(clknet_leaf_248_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23558_ (.D(_04435_),
    .Q(\design_top.core0.REG1[6][27] ),
    .CLK(clknet_leaf_249_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23559_ (.D(_04436_),
    .Q(\design_top.core0.REG1[6][28] ),
    .CLK(clknet_leaf_249_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23560_ (.D(_04437_),
    .Q(\design_top.core0.REG1[6][29] ),
    .CLK(clknet_leaf_248_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23561_ (.D(_04438_),
    .Q(\design_top.core0.REG1[6][30] ),
    .CLK(clknet_leaf_248_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23562_ (.D(_04439_),
    .Q(\design_top.core0.REG1[6][31] ),
    .CLK(clknet_leaf_248_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23563_ (.D(_04440_),
    .Q(\design_top.core0.REG1[7][0] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23564_ (.D(_04441_),
    .Q(\design_top.core0.REG1[7][1] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23565_ (.D(_04442_),
    .Q(\design_top.core0.REG1[7][2] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23566_ (.D(_04443_),
    .Q(\design_top.core0.REG1[7][3] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23567_ (.D(_04444_),
    .Q(\design_top.core0.REG1[7][4] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23568_ (.D(_04445_),
    .Q(\design_top.core0.REG1[7][5] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23569_ (.D(_04446_),
    .Q(\design_top.core0.REG1[7][6] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23570_ (.D(_04447_),
    .Q(\design_top.core0.REG1[7][7] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23571_ (.D(_04448_),
    .Q(\design_top.core0.REG1[7][8] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23572_ (.D(_04449_),
    .Q(\design_top.core0.REG1[7][9] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23573_ (.D(_04450_),
    .Q(\design_top.core0.REG1[7][10] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23574_ (.D(_04451_),
    .Q(\design_top.core0.REG1[7][11] ),
    .CLK(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23575_ (.D(_04452_),
    .Q(\design_top.core0.REG1[7][12] ),
    .CLK(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23576_ (.D(_04453_),
    .Q(\design_top.core0.REG1[7][13] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23577_ (.D(_04454_),
    .Q(\design_top.core0.REG1[7][14] ),
    .CLK(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23578_ (.D(_04455_),
    .Q(\design_top.core0.REG1[7][15] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23579_ (.D(_04456_),
    .Q(\design_top.core0.REG1[7][16] ),
    .CLK(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23580_ (.D(_04457_),
    .Q(\design_top.core0.REG1[7][17] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23581_ (.D(_04458_),
    .Q(\design_top.core0.REG1[7][18] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23582_ (.D(_04459_),
    .Q(\design_top.core0.REG1[7][19] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23583_ (.D(_04460_),
    .Q(\design_top.core0.REG1[7][20] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23584_ (.D(_04461_),
    .Q(\design_top.core0.REG1[7][21] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23585_ (.D(_04462_),
    .Q(\design_top.core0.REG1[7][22] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23586_ (.D(_04463_),
    .Q(\design_top.core0.REG1[7][23] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23587_ (.D(_04464_),
    .Q(\design_top.core0.REG1[7][24] ),
    .CLK(clknet_leaf_246_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23588_ (.D(_04465_),
    .Q(\design_top.core0.REG1[7][25] ),
    .CLK(clknet_leaf_246_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23589_ (.D(_04466_),
    .Q(\design_top.core0.REG1[7][26] ),
    .CLK(clknet_leaf_247_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23590_ (.D(_04467_),
    .Q(\design_top.core0.REG1[7][27] ),
    .CLK(clknet_leaf_249_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23591_ (.D(_04468_),
    .Q(\design_top.core0.REG1[7][28] ),
    .CLK(clknet_leaf_249_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23592_ (.D(_04469_),
    .Q(\design_top.core0.REG1[7][29] ),
    .CLK(clknet_leaf_246_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23593_ (.D(_04470_),
    .Q(\design_top.core0.REG1[7][30] ),
    .CLK(clknet_leaf_248_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23594_ (.D(_04471_),
    .Q(\design_top.core0.REG1[7][31] ),
    .CLK(clknet_leaf_248_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23595_ (.D(_04472_),
    .Q(\design_top.core0.REG1[8][0] ),
    .CLK(clknet_leaf_235_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23596_ (.D(_04473_),
    .Q(\design_top.core0.REG1[8][1] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23597_ (.D(_04474_),
    .Q(\design_top.core0.REG1[8][2] ),
    .CLK(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23598_ (.D(_04475_),
    .Q(\design_top.core0.REG1[8][3] ),
    .CLK(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23599_ (.D(_04476_),
    .Q(\design_top.core0.REG1[8][4] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23600_ (.D(_04477_),
    .Q(\design_top.core0.REG1[8][5] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23601_ (.D(_04478_),
    .Q(\design_top.core0.REG1[8][6] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23602_ (.D(_04479_),
    .Q(\design_top.core0.REG1[8][7] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23603_ (.D(_04480_),
    .Q(\design_top.core0.REG1[8][8] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23604_ (.D(_04481_),
    .Q(\design_top.core0.REG1[8][9] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23605_ (.D(_04482_),
    .Q(\design_top.core0.REG1[8][10] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23606_ (.D(_04483_),
    .Q(\design_top.core0.REG1[8][11] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23607_ (.D(_04484_),
    .Q(\design_top.core0.REG1[8][12] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23608_ (.D(_04485_),
    .Q(\design_top.core0.REG1[8][13] ),
    .CLK(clknet_leaf_235_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23609_ (.D(_04486_),
    .Q(\design_top.core0.REG1[8][14] ),
    .CLK(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23610_ (.D(_04487_),
    .Q(\design_top.core0.REG1[8][15] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23611_ (.D(_04488_),
    .Q(\design_top.core0.REG1[8][16] ),
    .CLK(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23612_ (.D(_04489_),
    .Q(\design_top.core0.REG1[8][17] ),
    .CLK(clknet_leaf_235_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23613_ (.D(_04490_),
    .Q(\design_top.core0.REG1[8][18] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23614_ (.D(_04491_),
    .Q(\design_top.core0.REG1[8][19] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23615_ (.D(_04492_),
    .Q(\design_top.core0.REG1[8][20] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23616_ (.D(_04493_),
    .Q(\design_top.core0.REG1[8][21] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23617_ (.D(_04494_),
    .Q(\design_top.core0.REG1[8][22] ),
    .CLK(clknet_leaf_262_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23618_ (.D(_04495_),
    .Q(\design_top.core0.REG1[8][23] ),
    .CLK(clknet_leaf_262_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23619_ (.D(_04496_),
    .Q(\design_top.core0.REG1[8][24] ),
    .CLK(clknet_leaf_262_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23620_ (.D(_04497_),
    .Q(\design_top.core0.REG1[8][25] ),
    .CLK(clknet_leaf_262_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23621_ (.D(_04498_),
    .Q(\design_top.core0.REG1[8][26] ),
    .CLK(clknet_leaf_262_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23622_ (.D(_04499_),
    .Q(\design_top.core0.REG1[8][27] ),
    .CLK(clknet_leaf_254_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23623_ (.D(_04500_),
    .Q(\design_top.core0.REG1[8][28] ),
    .CLK(clknet_leaf_255_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23624_ (.D(_04501_),
    .Q(\design_top.core0.REG1[8][29] ),
    .CLK(clknet_leaf_254_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23625_ (.D(_04502_),
    .Q(\design_top.core0.REG1[8][30] ),
    .CLK(clknet_leaf_254_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23626_ (.D(_04503_),
    .Q(\design_top.core0.REG1[8][31] ),
    .CLK(clknet_leaf_255_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23627_ (.D(_04504_),
    .Q(\design_top.core0.REG1[0][0] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23628_ (.D(_04505_),
    .Q(\design_top.core0.REG1[0][1] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23629_ (.D(_04506_),
    .Q(\design_top.core0.REG1[0][2] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23630_ (.D(_04507_),
    .Q(\design_top.core0.REG1[0][3] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23631_ (.D(_04508_),
    .Q(\design_top.core0.REG1[0][4] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23632_ (.D(_04509_),
    .Q(\design_top.core0.REG1[0][5] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23633_ (.D(_04510_),
    .Q(\design_top.core0.REG1[0][6] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23634_ (.D(_04511_),
    .Q(\design_top.core0.REG1[0][7] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23635_ (.D(_04512_),
    .Q(\design_top.core0.REG1[0][8] ),
    .CLK(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23636_ (.D(_04513_),
    .Q(\design_top.core0.REG1[0][9] ),
    .CLK(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23637_ (.D(_04514_),
    .Q(\design_top.core0.REG1[0][10] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23638_ (.D(_04515_),
    .Q(\design_top.core0.REG1[0][11] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23639_ (.D(_04516_),
    .Q(\design_top.core0.REG1[0][12] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23640_ (.D(_04517_),
    .Q(\design_top.core0.REG1[0][13] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23641_ (.D(_04518_),
    .Q(\design_top.core0.REG1[0][14] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23642_ (.D(_04519_),
    .Q(\design_top.core0.REG1[0][15] ),
    .CLK(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23643_ (.D(_04520_),
    .Q(\design_top.core0.REG1[0][16] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23644_ (.D(_04521_),
    .Q(\design_top.core0.REG1[0][17] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23645_ (.D(_04522_),
    .Q(\design_top.core0.REG1[0][18] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23646_ (.D(_04523_),
    .Q(\design_top.core0.REG1[0][19] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23647_ (.D(_04524_),
    .Q(\design_top.core0.REG1[0][20] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23648_ (.D(_04525_),
    .Q(\design_top.core0.REG1[0][21] ),
    .CLK(clknet_leaf_244_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23649_ (.D(_04526_),
    .Q(\design_top.core0.REG1[0][22] ),
    .CLK(clknet_leaf_244_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23650_ (.D(_04527_),
    .Q(\design_top.core0.REG1[0][23] ),
    .CLK(clknet_leaf_244_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23651_ (.D(_04528_),
    .Q(\design_top.core0.REG1[0][24] ),
    .CLK(clknet_leaf_244_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23652_ (.D(_04529_),
    .Q(\design_top.core0.REG1[0][25] ),
    .CLK(clknet_leaf_244_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23653_ (.D(_04530_),
    .Q(\design_top.core0.REG1[0][26] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23654_ (.D(_04531_),
    .Q(\design_top.core0.REG1[0][27] ),
    .CLK(clknet_leaf_250_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23655_ (.D(_04532_),
    .Q(\design_top.core0.REG1[0][28] ),
    .CLK(clknet_leaf_250_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23656_ (.D(_04533_),
    .Q(\design_top.core0.REG1[0][29] ),
    .CLK(clknet_leaf_251_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23657_ (.D(_04534_),
    .Q(\design_top.core0.REG1[0][30] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23658_ (.D(_04535_),
    .Q(\design_top.core0.REG1[0][31] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23659_ (.D(_04536_),
    .Q(\design_top.core0.REG1[10][0] ),
    .CLK(clknet_leaf_235_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23660_ (.D(_04537_),
    .Q(\design_top.core0.REG1[10][1] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23661_ (.D(_04538_),
    .Q(\design_top.core0.REG1[10][2] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23662_ (.D(_04539_),
    .Q(\design_top.core0.REG1[10][3] ),
    .CLK(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23663_ (.D(_04540_),
    .Q(\design_top.core0.REG1[10][4] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23664_ (.D(_04541_),
    .Q(\design_top.core0.REG1[10][5] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23665_ (.D(_04542_),
    .Q(\design_top.core0.REG1[10][6] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23666_ (.D(_04543_),
    .Q(\design_top.core0.REG1[10][7] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23667_ (.D(_04544_),
    .Q(\design_top.core0.REG1[10][8] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23668_ (.D(_04545_),
    .Q(\design_top.core0.REG1[10][9] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23669_ (.D(_04546_),
    .Q(\design_top.core0.REG1[10][10] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23670_ (.D(_04547_),
    .Q(\design_top.core0.REG1[10][11] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23671_ (.D(_04548_),
    .Q(\design_top.core0.REG1[10][12] ),
    .CLK(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23672_ (.D(_04549_),
    .Q(\design_top.core0.REG1[10][13] ),
    .CLK(clknet_leaf_235_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23673_ (.D(_04550_),
    .Q(\design_top.core0.REG1[10][14] ),
    .CLK(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23674_ (.D(_04551_),
    .Q(\design_top.core0.REG1[10][15] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23675_ (.D(_04552_),
    .Q(\design_top.core0.REG1[10][16] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23676_ (.D(_04553_),
    .Q(\design_top.core0.REG1[10][17] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23677_ (.D(_04554_),
    .Q(\design_top.core0.REG1[10][18] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23678_ (.D(_04555_),
    .Q(\design_top.core0.REG1[10][19] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23679_ (.D(_04556_),
    .Q(\design_top.core0.REG1[10][20] ),
    .CLK(clknet_leaf_262_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23680_ (.D(_04557_),
    .Q(\design_top.core0.REG1[10][21] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23681_ (.D(_04558_),
    .Q(\design_top.core0.REG1[10][22] ),
    .CLK(clknet_leaf_262_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23682_ (.D(_04559_),
    .Q(\design_top.core0.REG1[10][23] ),
    .CLK(clknet_leaf_262_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23683_ (.D(_04560_),
    .Q(\design_top.core0.REG1[10][24] ),
    .CLK(clknet_leaf_262_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23684_ (.D(_04561_),
    .Q(\design_top.core0.REG1[10][25] ),
    .CLK(clknet_leaf_253_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23685_ (.D(_04562_),
    .Q(\design_top.core0.REG1[10][26] ),
    .CLK(clknet_leaf_253_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23686_ (.D(_04563_),
    .Q(\design_top.core0.REG1[10][27] ),
    .CLK(clknet_leaf_255_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23687_ (.D(_04564_),
    .Q(\design_top.core0.REG1[10][28] ),
    .CLK(clknet_leaf_255_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23688_ (.D(_04565_),
    .Q(\design_top.core0.REG1[10][29] ),
    .CLK(clknet_leaf_254_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23689_ (.D(_04566_),
    .Q(\design_top.core0.REG1[10][30] ),
    .CLK(clknet_leaf_254_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23690_ (.D(_04567_),
    .Q(\design_top.core0.REG1[10][31] ),
    .CLK(clknet_leaf_255_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23691_ (.D(_04568_),
    .Q(\design_top.core0.REG1[11][0] ),
    .CLK(clknet_leaf_235_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23692_ (.D(_04569_),
    .Q(\design_top.core0.REG1[11][1] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23693_ (.D(_04570_),
    .Q(\design_top.core0.REG1[11][2] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23694_ (.D(_04571_),
    .Q(\design_top.core0.REG1[11][3] ),
    .CLK(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23695_ (.D(_04572_),
    .Q(\design_top.core0.REG1[11][4] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23696_ (.D(_04573_),
    .Q(\design_top.core0.REG1[11][5] ),
    .CLK(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23697_ (.D(_04574_),
    .Q(\design_top.core0.REG1[11][6] ),
    .CLK(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23698_ (.D(_04575_),
    .Q(\design_top.core0.REG1[11][7] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23699_ (.D(_04576_),
    .Q(\design_top.core0.REG1[11][8] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23700_ (.D(_04577_),
    .Q(\design_top.core0.REG1[11][9] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23701_ (.D(_04578_),
    .Q(\design_top.core0.REG1[11][10] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23702_ (.D(_04579_),
    .Q(\design_top.core0.REG1[11][11] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23703_ (.D(_04580_),
    .Q(\design_top.core0.REG1[11][12] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23704_ (.D(_04581_),
    .Q(\design_top.core0.REG1[11][13] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23705_ (.D(_04582_),
    .Q(\design_top.core0.REG1[11][14] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23706_ (.D(_04583_),
    .Q(\design_top.core0.REG1[11][15] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23707_ (.D(_04584_),
    .Q(\design_top.core0.REG1[11][16] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23708_ (.D(_04585_),
    .Q(\design_top.core0.REG1[11][17] ),
    .CLK(clknet_leaf_235_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23709_ (.D(_04586_),
    .Q(\design_top.core0.REG1[11][18] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23710_ (.D(_04587_),
    .Q(\design_top.core0.REG1[11][19] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23711_ (.D(_04588_),
    .Q(\design_top.core0.REG1[11][20] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23712_ (.D(_04589_),
    .Q(\design_top.core0.REG1[11][21] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23713_ (.D(_04590_),
    .Q(\design_top.core0.REG1[11][22] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23714_ (.D(_04591_),
    .Q(\design_top.core0.REG1[11][23] ),
    .CLK(clknet_leaf_262_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23715_ (.D(_04592_),
    .Q(\design_top.core0.REG1[11][24] ),
    .CLK(clknet_leaf_261_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23716_ (.D(_04593_),
    .Q(\design_top.core0.REG1[11][25] ),
    .CLK(clknet_leaf_253_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23717_ (.D(_04594_),
    .Q(\design_top.core0.REG1[11][26] ),
    .CLK(clknet_leaf_253_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23718_ (.D(_04595_),
    .Q(\design_top.core0.REG1[11][27] ),
    .CLK(clknet_leaf_255_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23719_ (.D(_04596_),
    .Q(\design_top.core0.REG1[11][28] ),
    .CLK(clknet_leaf_255_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23720_ (.D(_04597_),
    .Q(\design_top.core0.REG1[11][29] ),
    .CLK(clknet_leaf_254_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23721_ (.D(_04598_),
    .Q(\design_top.core0.REG1[11][30] ),
    .CLK(clknet_leaf_254_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23722_ (.D(_04599_),
    .Q(\design_top.core0.REG1[11][31] ),
    .CLK(clknet_leaf_255_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23723_ (.D(_04600_),
    .Q(\design_top.core0.REG1[12][0] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23724_ (.D(_04601_),
    .Q(\design_top.core0.REG1[12][1] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23725_ (.D(_04602_),
    .Q(\design_top.core0.REG1[12][2] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23726_ (.D(_04603_),
    .Q(\design_top.core0.REG1[12][3] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23727_ (.D(_04604_),
    .Q(\design_top.core0.REG1[12][4] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23728_ (.D(_04605_),
    .Q(\design_top.core0.REG1[12][5] ),
    .CLK(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23729_ (.D(_04606_),
    .Q(\design_top.core0.REG1[12][6] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23730_ (.D(_04607_),
    .Q(\design_top.core0.REG1[12][7] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23731_ (.D(_04608_),
    .Q(\design_top.core0.REG1[12][8] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23732_ (.D(_04609_),
    .Q(\design_top.core0.REG1[12][9] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23733_ (.D(_04610_),
    .Q(\design_top.core0.REG1[12][10] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23734_ (.D(_04611_),
    .Q(\design_top.core0.REG1[12][11] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23735_ (.D(_04612_),
    .Q(\design_top.core0.REG1[12][12] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23736_ (.D(_04613_),
    .Q(\design_top.core0.REG1[12][13] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23737_ (.D(_04614_),
    .Q(\design_top.core0.REG1[12][14] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23738_ (.D(_04615_),
    .Q(\design_top.core0.REG1[12][15] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23739_ (.D(_04616_),
    .Q(\design_top.core0.REG1[12][16] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23740_ (.D(_04617_),
    .Q(\design_top.core0.REG1[12][17] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23741_ (.D(_04618_),
    .Q(\design_top.core0.REG1[12][18] ),
    .CLK(clknet_leaf_263_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23742_ (.D(_04619_),
    .Q(\design_top.core0.REG1[12][19] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23743_ (.D(_04620_),
    .Q(\design_top.core0.REG1[12][20] ),
    .CLK(clknet_leaf_262_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23744_ (.D(_04621_),
    .Q(\design_top.core0.REG1[12][21] ),
    .CLK(clknet_leaf_262_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23745_ (.D(_04622_),
    .Q(\design_top.core0.REG1[12][22] ),
    .CLK(clknet_leaf_264_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23746_ (.D(_04623_),
    .Q(\design_top.core0.REG1[12][23] ),
    .CLK(clknet_leaf_263_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23747_ (.D(_04624_),
    .Q(\design_top.core0.REG1[12][24] ),
    .CLK(clknet_leaf_261_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23748_ (.D(_04625_),
    .Q(\design_top.core0.REG1[12][25] ),
    .CLK(clknet_leaf_260_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23749_ (.D(_04626_),
    .Q(\design_top.core0.REG1[12][26] ),
    .CLK(clknet_leaf_261_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23750_ (.D(_04627_),
    .Q(\design_top.core0.REG1[12][27] ),
    .CLK(clknet_leaf_256_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23751_ (.D(_04628_),
    .Q(\design_top.core0.REG1[12][28] ),
    .CLK(clknet_leaf_256_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23752_ (.D(_04629_),
    .Q(\design_top.core0.REG1[12][29] ),
    .CLK(clknet_leaf_254_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23753_ (.D(_04630_),
    .Q(\design_top.core0.REG1[12][30] ),
    .CLK(clknet_leaf_254_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23754_ (.D(_04631_),
    .Q(\design_top.core0.REG1[12][31] ),
    .CLK(clknet_leaf_256_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23755_ (.D(_04632_),
    .Q(\design_top.core0.REG1[13][0] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23756_ (.D(_04633_),
    .Q(\design_top.core0.REG1[13][1] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23757_ (.D(_04634_),
    .Q(\design_top.core0.REG1[13][2] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23758_ (.D(_04635_),
    .Q(\design_top.core0.REG1[13][3] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23759_ (.D(_04636_),
    .Q(\design_top.core0.REG1[13][4] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23760_ (.D(_04637_),
    .Q(\design_top.core0.REG1[13][5] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23761_ (.D(_04638_),
    .Q(\design_top.core0.REG1[13][6] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23762_ (.D(_04639_),
    .Q(\design_top.core0.REG1[13][7] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23763_ (.D(_04640_),
    .Q(\design_top.core0.REG1[13][8] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23764_ (.D(_04641_),
    .Q(\design_top.core0.REG1[13][9] ),
    .CLK(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23765_ (.D(_04642_),
    .Q(\design_top.core0.REG1[13][10] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23766_ (.D(_04643_),
    .Q(\design_top.core0.REG1[13][11] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23767_ (.D(_04644_),
    .Q(\design_top.core0.REG1[13][12] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23768_ (.D(_04645_),
    .Q(\design_top.core0.REG1[13][13] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23769_ (.D(_04646_),
    .Q(\design_top.core0.REG1[13][14] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23770_ (.D(_04647_),
    .Q(\design_top.core0.REG1[13][15] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23771_ (.D(_04648_),
    .Q(\design_top.core0.REG1[13][16] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23772_ (.D(_04649_),
    .Q(\design_top.core0.REG1[13][17] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23773_ (.D(_04650_),
    .Q(\design_top.core0.REG1[13][18] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23774_ (.D(_04651_),
    .Q(\design_top.core0.REG1[13][19] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23775_ (.D(_04652_),
    .Q(\design_top.core0.REG1[13][20] ),
    .CLK(clknet_leaf_263_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23776_ (.D(_04653_),
    .Q(\design_top.core0.REG1[13][21] ),
    .CLK(clknet_leaf_263_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23777_ (.D(_04654_),
    .Q(\design_top.core0.REG1[13][22] ),
    .CLK(clknet_leaf_263_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23778_ (.D(_04655_),
    .Q(\design_top.core0.REG1[13][23] ),
    .CLK(clknet_leaf_263_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23779_ (.D(_04656_),
    .Q(\design_top.core0.REG1[13][24] ),
    .CLK(clknet_leaf_261_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23780_ (.D(_04657_),
    .Q(\design_top.core0.REG1[13][25] ),
    .CLK(clknet_leaf_260_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23781_ (.D(_04658_),
    .Q(\design_top.core0.REG1[13][26] ),
    .CLK(clknet_leaf_261_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23782_ (.D(_04659_),
    .Q(\design_top.core0.REG1[13][27] ),
    .CLK(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23783_ (.D(_04660_),
    .Q(\design_top.core0.REG1[13][28] ),
    .CLK(clknet_leaf_256_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23784_ (.D(_04661_),
    .Q(\design_top.core0.REG1[13][29] ),
    .CLK(clknet_leaf_256_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23785_ (.D(_04662_),
    .Q(\design_top.core0.REG1[13][30] ),
    .CLK(clknet_leaf_261_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23786_ (.D(_04663_),
    .Q(\design_top.core0.REG1[13][31] ),
    .CLK(clknet_leaf_256_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23787_ (.D(_04664_),
    .Q(\design_top.core0.REG1[14][0] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23788_ (.D(_04665_),
    .Q(\design_top.core0.REG1[14][1] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23789_ (.D(_04666_),
    .Q(\design_top.core0.REG1[14][2] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23790_ (.D(_04667_),
    .Q(\design_top.core0.REG1[14][3] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23791_ (.D(_04668_),
    .Q(\design_top.core0.REG1[14][4] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23792_ (.D(_04669_),
    .Q(\design_top.core0.REG1[14][5] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23793_ (.D(_04670_),
    .Q(\design_top.core0.REG1[14][6] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23794_ (.D(_04671_),
    .Q(\design_top.core0.REG1[14][7] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23795_ (.D(_04672_),
    .Q(\design_top.core0.REG1[14][8] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23796_ (.D(_04673_),
    .Q(\design_top.core0.REG1[14][9] ),
    .CLK(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23797_ (.D(_04674_),
    .Q(\design_top.core0.REG1[14][10] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23798_ (.D(_04675_),
    .Q(\design_top.core0.REG1[14][11] ),
    .CLK(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23799_ (.D(_04676_),
    .Q(\design_top.core0.REG1[14][12] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23800_ (.D(_04677_),
    .Q(\design_top.core0.REG1[14][13] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23801_ (.D(_04678_),
    .Q(\design_top.core0.REG1[14][14] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23802_ (.D(_04679_),
    .Q(\design_top.core0.REG1[14][15] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23803_ (.D(_04680_),
    .Q(\design_top.core0.REG1[14][16] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23804_ (.D(_04681_),
    .Q(\design_top.core0.REG1[14][17] ),
    .CLK(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23805_ (.D(_04682_),
    .Q(\design_top.core0.REG1[14][18] ),
    .CLK(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23806_ (.D(_04683_),
    .Q(\design_top.core0.REG1[14][19] ),
    .CLK(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23807_ (.D(_04684_),
    .Q(\design_top.core0.REG1[14][20] ),
    .CLK(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23808_ (.D(_04685_),
    .Q(\design_top.core0.REG1[14][21] ),
    .CLK(clknet_leaf_263_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23809_ (.D(_04686_),
    .Q(\design_top.core0.REG1[14][22] ),
    .CLK(clknet_leaf_259_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23810_ (.D(_04687_),
    .Q(\design_top.core0.REG1[14][23] ),
    .CLK(clknet_leaf_259_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23811_ (.D(_04688_),
    .Q(\design_top.core0.REG1[14][24] ),
    .CLK(clknet_leaf_259_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23812_ (.D(_04689_),
    .Q(\design_top.core0.REG1[14][25] ),
    .CLK(clknet_leaf_259_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23813_ (.D(_04690_),
    .Q(\design_top.core0.REG1[14][26] ),
    .CLK(clknet_leaf_259_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23814_ (.D(_04691_),
    .Q(\design_top.core0.REG1[14][27] ),
    .CLK(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23815_ (.D(_04692_),
    .Q(\design_top.core0.REG1[14][28] ),
    .CLK(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23816_ (.D(_04693_),
    .Q(\design_top.core0.REG1[14][29] ),
    .CLK(clknet_leaf_259_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23817_ (.D(_04694_),
    .Q(\design_top.core0.REG1[14][30] ),
    .CLK(clknet_leaf_259_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23818_ (.D(_04695_),
    .Q(\design_top.core0.REG1[14][31] ),
    .CLK(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23819_ (.D(_04696_),
    .Q(\design_top.MEM[62][0] ),
    .CLK(clknet_leaf_402_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23820_ (.D(_04697_),
    .Q(\design_top.MEM[62][1] ),
    .CLK(clknet_leaf_405_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23821_ (.D(_04698_),
    .Q(\design_top.MEM[62][2] ),
    .CLK(clknet_leaf_405_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23822_ (.D(_04699_),
    .Q(\design_top.MEM[62][3] ),
    .CLK(clknet_leaf_413_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23823_ (.D(_04700_),
    .Q(\design_top.MEM[62][4] ),
    .CLK(clknet_leaf_412_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23824_ (.D(_04701_),
    .Q(\design_top.MEM[62][5] ),
    .CLK(clknet_leaf_406_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23825_ (.D(_04702_),
    .Q(\design_top.MEM[62][6] ),
    .CLK(clknet_leaf_406_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23826_ (.D(_04703_),
    .Q(\design_top.MEM[62][7] ),
    .CLK(clknet_leaf_429_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23827_ (.D(_04704_),
    .Q(\design_top.MEM[63][0] ),
    .CLK(clknet_leaf_405_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23828_ (.D(_04705_),
    .Q(\design_top.MEM[63][1] ),
    .CLK(clknet_leaf_430_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23829_ (.D(_04706_),
    .Q(\design_top.MEM[63][2] ),
    .CLK(clknet_leaf_405_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23830_ (.D(_04707_),
    .Q(\design_top.MEM[63][3] ),
    .CLK(clknet_leaf_429_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23831_ (.D(_04708_),
    .Q(\design_top.MEM[63][4] ),
    .CLK(clknet_leaf_421_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23832_ (.D(_04709_),
    .Q(\design_top.MEM[63][5] ),
    .CLK(clknet_leaf_422_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23833_ (.D(_04710_),
    .Q(\design_top.MEM[63][6] ),
    .CLK(clknet_leaf_421_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23834_ (.D(_04711_),
    .Q(\design_top.MEM[63][7] ),
    .CLK(clknet_leaf_422_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23835_ (.D(_04712_),
    .Q(\design_top.MEM[6][0] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23836_ (.D(_04713_),
    .Q(\design_top.MEM[6][1] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23837_ (.D(_04714_),
    .Q(\design_top.MEM[6][2] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23838_ (.D(_04715_),
    .Q(\design_top.MEM[6][3] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23839_ (.D(_04716_),
    .Q(\design_top.MEM[6][4] ),
    .CLK(clknet_leaf_403_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23840_ (.D(_04717_),
    .Q(\design_top.MEM[6][5] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23841_ (.D(_04718_),
    .Q(\design_top.MEM[6][6] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23842_ (.D(_04719_),
    .Q(\design_top.MEM[6][7] ),
    .CLK(clknet_leaf_401_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23843_ (.D(_04720_),
    .Q(\design_top.core0.REG2[15][0] ),
    .CLK(clknet_leaf_266_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23844_ (.D(_04721_),
    .Q(\design_top.core0.REG2[15][1] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23845_ (.D(_04722_),
    .Q(\design_top.core0.REG2[15][2] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23846_ (.D(_04723_),
    .Q(\design_top.core0.REG2[15][3] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23847_ (.D(_04724_),
    .Q(\design_top.core0.REG2[15][4] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23848_ (.D(_04725_),
    .Q(\design_top.core0.REG2[15][5] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23849_ (.D(_04726_),
    .Q(\design_top.core0.REG2[15][6] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23850_ (.D(_04727_),
    .Q(\design_top.core0.REG2[15][7] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23851_ (.D(_04728_),
    .Q(\design_top.core0.REG2[15][8] ),
    .CLK(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23852_ (.D(_04729_),
    .Q(\design_top.core0.REG2[15][9] ),
    .CLK(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23853_ (.D(_04730_),
    .Q(\design_top.core0.REG2[15][10] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23854_ (.D(_04731_),
    .Q(\design_top.core0.REG2[15][11] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23855_ (.D(_04732_),
    .Q(\design_top.core0.REG2[15][12] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23856_ (.D(_04733_),
    .Q(\design_top.core0.REG2[15][13] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23857_ (.D(_04734_),
    .Q(\design_top.core0.REG2[15][14] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23858_ (.D(_04735_),
    .Q(\design_top.core0.REG2[15][15] ),
    .CLK(clknet_leaf_298_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23859_ (.D(_04736_),
    .Q(\design_top.core0.REG2[15][16] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23860_ (.D(_04737_),
    .Q(\design_top.core0.REG2[15][17] ),
    .CLK(clknet_leaf_266_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23861_ (.D(_04738_),
    .Q(\design_top.core0.REG2[15][18] ),
    .CLK(clknet_leaf_267_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23862_ (.D(_04739_),
    .Q(\design_top.core0.REG2[15][19] ),
    .CLK(clknet_leaf_267_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23863_ (.D(_04740_),
    .Q(\design_top.core0.REG2[15][20] ),
    .CLK(clknet_leaf_268_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23864_ (.D(_04741_),
    .Q(\design_top.core0.REG2[15][21] ),
    .CLK(clknet_leaf_268_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23865_ (.D(_04742_),
    .Q(\design_top.core0.REG2[15][22] ),
    .CLK(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23866_ (.D(_04743_),
    .Q(\design_top.core0.REG2[15][23] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23867_ (.D(_04744_),
    .Q(\design_top.core0.REG2[15][24] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23868_ (.D(_04745_),
    .Q(\design_top.core0.REG2[15][25] ),
    .CLK(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23869_ (.D(_04746_),
    .Q(\design_top.core0.REG2[15][26] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23870_ (.D(_04747_),
    .Q(\design_top.core0.REG2[15][27] ),
    .CLK(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23871_ (.D(_04748_),
    .Q(\design_top.core0.REG2[15][28] ),
    .CLK(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23872_ (.D(_04749_),
    .Q(\design_top.core0.REG2[15][29] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23873_ (.D(_04750_),
    .Q(\design_top.core0.REG2[15][30] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23874_ (.D(_04751_),
    .Q(\design_top.core0.REG2[15][31] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23875_ (.D(_04752_),
    .Q(\design_top.core0.REG2[1][0] ),
    .CLK(clknet_leaf_266_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23876_ (.D(_04753_),
    .Q(\design_top.core0.REG2[1][1] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23877_ (.D(_04754_),
    .Q(\design_top.core0.REG2[1][2] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23878_ (.D(_04755_),
    .Q(\design_top.core0.REG2[1][3] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23879_ (.D(_04756_),
    .Q(\design_top.core0.REG2[1][4] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23880_ (.D(_04757_),
    .Q(\design_top.core0.REG2[1][5] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23881_ (.D(_04758_),
    .Q(\design_top.core0.REG2[1][6] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23882_ (.D(_04759_),
    .Q(\design_top.core0.REG2[1][7] ),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23883_ (.D(_04760_),
    .Q(\design_top.core0.REG2[1][8] ),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23884_ (.D(_04761_),
    .Q(\design_top.core0.REG2[1][9] ),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23885_ (.D(_04762_),
    .Q(\design_top.core0.REG2[1][10] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23886_ (.D(_04763_),
    .Q(\design_top.core0.REG2[1][11] ),
    .CLK(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23887_ (.D(_04764_),
    .Q(\design_top.core0.REG2[1][12] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23888_ (.D(_04765_),
    .Q(\design_top.core0.REG2[1][13] ),
    .CLK(clknet_leaf_298_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23889_ (.D(_04766_),
    .Q(\design_top.core0.REG2[1][14] ),
    .CLK(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23890_ (.D(_04767_),
    .Q(\design_top.core0.REG2[1][15] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23891_ (.D(_04768_),
    .Q(\design_top.core0.REG2[1][16] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23892_ (.D(_04769_),
    .Q(\design_top.core0.REG2[1][17] ),
    .CLK(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23893_ (.D(_04770_),
    .Q(\design_top.core0.REG2[1][18] ),
    .CLK(clknet_leaf_266_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23894_ (.D(_04771_),
    .Q(\design_top.core0.REG2[1][19] ),
    .CLK(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23895_ (.D(_04772_),
    .Q(\design_top.core0.REG2[1][20] ),
    .CLK(clknet_leaf_268_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23896_ (.D(_04773_),
    .Q(\design_top.core0.REG2[1][21] ),
    .CLK(clknet_leaf_264_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23897_ (.D(_04774_),
    .Q(\design_top.core0.REG2[1][22] ),
    .CLK(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23898_ (.D(_04775_),
    .Q(\design_top.core0.REG2[1][23] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23899_ (.D(_04776_),
    .Q(\design_top.core0.REG2[1][24] ),
    .CLK(clknet_leaf_281_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23900_ (.D(_04777_),
    .Q(\design_top.core0.REG2[1][25] ),
    .CLK(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23901_ (.D(_04778_),
    .Q(\design_top.core0.REG2[1][26] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23902_ (.D(_04779_),
    .Q(\design_top.core0.REG2[1][27] ),
    .CLK(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23903_ (.D(_04780_),
    .Q(\design_top.core0.REG2[1][28] ),
    .CLK(clknet_leaf_258_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23904_ (.D(_04781_),
    .Q(\design_top.core0.REG2[1][29] ),
    .CLK(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23905_ (.D(_04782_),
    .Q(\design_top.core0.REG2[1][30] ),
    .CLK(clknet_leaf_258_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23906_ (.D(_04783_),
    .Q(\design_top.core0.REG2[1][31] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23907_ (.D(_04784_),
    .Q(\design_top.core0.REG2[2][0] ),
    .CLK(clknet_leaf_266_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23908_ (.D(_04785_),
    .Q(\design_top.core0.REG2[2][1] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23909_ (.D(_04786_),
    .Q(\design_top.core0.REG2[2][2] ),
    .CLK(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23910_ (.D(_04787_),
    .Q(\design_top.core0.REG2[2][3] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23911_ (.D(_04788_),
    .Q(\design_top.core0.REG2[2][4] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23912_ (.D(_04789_),
    .Q(\design_top.core0.REG2[2][5] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23913_ (.D(_04790_),
    .Q(\design_top.core0.REG2[2][6] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23914_ (.D(_04791_),
    .Q(\design_top.core0.REG2[2][7] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23915_ (.D(_04792_),
    .Q(\design_top.core0.REG2[2][8] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23916_ (.D(_04793_),
    .Q(\design_top.core0.REG2[2][9] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23917_ (.D(_04794_),
    .Q(\design_top.core0.REG2[2][10] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23918_ (.D(_04795_),
    .Q(\design_top.core0.REG2[2][11] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23919_ (.D(_04796_),
    .Q(\design_top.core0.REG2[2][12] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23920_ (.D(_04797_),
    .Q(\design_top.core0.REG2[2][13] ),
    .CLK(clknet_leaf_267_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23921_ (.D(_04798_),
    .Q(\design_top.core0.REG2[2][14] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23922_ (.D(_04799_),
    .Q(\design_top.core0.REG2[2][15] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23923_ (.D(_04800_),
    .Q(\design_top.core0.REG2[2][16] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23924_ (.D(_04801_),
    .Q(\design_top.core0.REG2[2][17] ),
    .CLK(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23925_ (.D(_04802_),
    .Q(\design_top.core0.REG2[2][18] ),
    .CLK(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23926_ (.D(_04803_),
    .Q(\design_top.core0.REG2[2][19] ),
    .CLK(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23927_ (.D(_04804_),
    .Q(\design_top.core0.REG2[2][20] ),
    .CLK(clknet_leaf_264_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23928_ (.D(_04805_),
    .Q(\design_top.core0.REG2[2][21] ),
    .CLK(clknet_leaf_264_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23929_ (.D(_04806_),
    .Q(\design_top.core0.REG2[2][22] ),
    .CLK(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23930_ (.D(_04807_),
    .Q(\design_top.core0.REG2[2][23] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23931_ (.D(_04808_),
    .Q(\design_top.core0.REG2[2][24] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23932_ (.D(_04809_),
    .Q(\design_top.core0.REG2[2][25] ),
    .CLK(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23933_ (.D(_04810_),
    .Q(\design_top.core0.REG2[2][26] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23934_ (.D(_04811_),
    .Q(\design_top.core0.REG2[2][27] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23935_ (.D(_04812_),
    .Q(\design_top.core0.REG2[2][28] ),
    .CLK(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23936_ (.D(_04813_),
    .Q(\design_top.core0.REG2[2][29] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23937_ (.D(_04814_),
    .Q(\design_top.core0.REG2[2][30] ),
    .CLK(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23938_ (.D(_04815_),
    .Q(\design_top.core0.REG2[2][31] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23939_ (.D(_04816_),
    .Q(\design_top.core0.REG2[3][0] ),
    .CLK(clknet_leaf_266_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23940_ (.D(_04817_),
    .Q(\design_top.core0.REG2[3][1] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23941_ (.D(_04818_),
    .Q(\design_top.core0.REG2[3][2] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23942_ (.D(_04819_),
    .Q(\design_top.core0.REG2[3][3] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23943_ (.D(_04820_),
    .Q(\design_top.core0.REG2[3][4] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23944_ (.D(_04821_),
    .Q(\design_top.core0.REG2[3][5] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23945_ (.D(_04822_),
    .Q(\design_top.core0.REG2[3][6] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23946_ (.D(_04823_),
    .Q(\design_top.core0.REG2[3][7] ),
    .CLK(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23947_ (.D(_04824_),
    .Q(\design_top.core0.REG2[3][8] ),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23948_ (.D(_04825_),
    .Q(\design_top.core0.REG2[3][9] ),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23949_ (.D(_04826_),
    .Q(\design_top.core0.REG2[3][10] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23950_ (.D(_04827_),
    .Q(\design_top.core0.REG2[3][11] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23951_ (.D(_04828_),
    .Q(\design_top.core0.REG2[3][12] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23952_ (.D(_04829_),
    .Q(\design_top.core0.REG2[3][13] ),
    .CLK(clknet_leaf_266_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23953_ (.D(_04830_),
    .Q(\design_top.core0.REG2[3][14] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23954_ (.D(_04831_),
    .Q(\design_top.core0.REG2[3][15] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23955_ (.D(_04832_),
    .Q(\design_top.core0.REG2[3][16] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23956_ (.D(_04833_),
    .Q(\design_top.core0.REG2[3][17] ),
    .CLK(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23957_ (.D(_04834_),
    .Q(\design_top.core0.REG2[3][18] ),
    .CLK(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23958_ (.D(_04835_),
    .Q(\design_top.core0.REG2[3][19] ),
    .CLK(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23959_ (.D(_04836_),
    .Q(\design_top.core0.REG2[3][20] ),
    .CLK(clknet_leaf_264_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23960_ (.D(_04837_),
    .Q(\design_top.core0.REG2[3][21] ),
    .CLK(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23961_ (.D(_04838_),
    .Q(\design_top.core0.REG2[3][22] ),
    .CLK(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23962_ (.D(_04839_),
    .Q(\design_top.core0.REG2[3][23] ),
    .CLK(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23963_ (.D(_04840_),
    .Q(\design_top.core0.REG2[3][24] ),
    .CLK(clknet_leaf_281_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23964_ (.D(_04841_),
    .Q(\design_top.core0.REG2[3][25] ),
    .CLK(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23965_ (.D(_04842_),
    .Q(\design_top.core0.REG2[3][26] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23966_ (.D(_04843_),
    .Q(\design_top.core0.REG2[3][27] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23967_ (.D(_04844_),
    .Q(\design_top.core0.REG2[3][28] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23968_ (.D(_04845_),
    .Q(\design_top.core0.REG2[3][29] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23969_ (.D(_04846_),
    .Q(\design_top.core0.REG2[3][30] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23970_ (.D(_04847_),
    .Q(\design_top.core0.REG2[3][31] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23971_ (.D(_04848_),
    .Q(\design_top.core0.REG2[4][0] ),
    .CLK(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23972_ (.D(_04849_),
    .Q(\design_top.core0.REG2[4][1] ),
    .CLK(clknet_leaf_302_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23973_ (.D(_04850_),
    .Q(\design_top.core0.REG2[4][2] ),
    .CLK(clknet_leaf_309_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23974_ (.D(_04851_),
    .Q(\design_top.core0.REG2[4][3] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23975_ (.D(_04852_),
    .Q(\design_top.core0.REG2[4][4] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23976_ (.D(_04853_),
    .Q(\design_top.core0.REG2[4][5] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23977_ (.D(_04854_),
    .Q(\design_top.core0.REG2[4][6] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23978_ (.D(_04855_),
    .Q(\design_top.core0.REG2[4][7] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23979_ (.D(_04856_),
    .Q(\design_top.core0.REG2[4][8] ),
    .CLK(clknet_leaf_187_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23980_ (.D(_04857_),
    .Q(\design_top.core0.REG2[4][9] ),
    .CLK(clknet_leaf_187_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23981_ (.D(_04858_),
    .Q(\design_top.core0.REG2[4][10] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23982_ (.D(_04859_),
    .Q(\design_top.core0.REG2[4][11] ),
    .CLK(clknet_leaf_302_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23983_ (.D(_04860_),
    .Q(\design_top.core0.REG2[4][12] ),
    .CLK(clknet_leaf_300_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23984_ (.D(_04861_),
    .Q(\design_top.core0.REG2[4][13] ),
    .CLK(clknet_leaf_295_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23985_ (.D(_04862_),
    .Q(\design_top.core0.REG2[4][14] ),
    .CLK(clknet_leaf_302_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23986_ (.D(_04863_),
    .Q(\design_top.core0.REG2[4][15] ),
    .CLK(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23987_ (.D(_04864_),
    .Q(\design_top.core0.REG2[4][16] ),
    .CLK(clknet_leaf_300_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23988_ (.D(_04865_),
    .Q(\design_top.core0.REG2[4][17] ),
    .CLK(clknet_leaf_292_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23989_ (.D(_04866_),
    .Q(\design_top.core0.REG2[4][18] ),
    .CLK(clknet_leaf_292_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23990_ (.D(_04867_),
    .Q(\design_top.core0.REG2[4][19] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23991_ (.D(_04868_),
    .Q(\design_top.core0.REG2[4][20] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23992_ (.D(_04869_),
    .Q(\design_top.core0.REG2[4][21] ),
    .CLK(clknet_leaf_294_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23993_ (.D(_04870_),
    .Q(\design_top.core0.REG2[4][22] ),
    .CLK(clknet_leaf_270_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23994_ (.D(_04871_),
    .Q(\design_top.core0.REG2[4][23] ),
    .CLK(clknet_leaf_287_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23995_ (.D(_04872_),
    .Q(\design_top.core0.REG2[4][24] ),
    .CLK(clknet_leaf_287_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23996_ (.D(_04873_),
    .Q(\design_top.core0.REG2[4][25] ),
    .CLK(clknet_leaf_294_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23997_ (.D(_04874_),
    .Q(\design_top.core0.REG2[4][26] ),
    .CLK(clknet_leaf_287_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23998_ (.D(_04875_),
    .Q(\design_top.core0.REG2[4][27] ),
    .CLK(clknet_leaf_270_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _23999_ (.D(_04876_),
    .Q(\design_top.core0.REG2[4][28] ),
    .CLK(clknet_leaf_268_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24000_ (.D(_04877_),
    .Q(\design_top.core0.REG2[4][29] ),
    .CLK(clknet_leaf_270_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24001_ (.D(_04878_),
    .Q(\design_top.core0.REG2[4][30] ),
    .CLK(clknet_leaf_264_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24002_ (.D(_04879_),
    .Q(\design_top.core0.REG2[4][31] ),
    .CLK(clknet_leaf_272_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24003_ (.D(_04880_),
    .Q(\design_top.MEM[7][0] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24004_ (.D(_04881_),
    .Q(\design_top.MEM[7][1] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24005_ (.D(_04882_),
    .Q(\design_top.MEM[7][2] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24006_ (.D(_04883_),
    .Q(\design_top.MEM[7][3] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24007_ (.D(_04884_),
    .Q(\design_top.MEM[7][4] ),
    .CLK(clknet_leaf_403_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24008_ (.D(_04885_),
    .Q(\design_top.MEM[7][5] ),
    .CLK(clknet_leaf_403_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24009_ (.D(_04886_),
    .Q(\design_top.MEM[7][6] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24010_ (.D(_04887_),
    .Q(\design_top.MEM[7][7] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24011_ (.D(_04888_),
    .Q(\design_top.core0.REG2[5][0] ),
    .CLK(clknet_leaf_296_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24012_ (.D(_04889_),
    .Q(\design_top.core0.REG2[5][1] ),
    .CLK(clknet_leaf_310_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24013_ (.D(_04890_),
    .Q(\design_top.core0.REG2[5][2] ),
    .CLK(clknet_leaf_310_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24014_ (.D(_04891_),
    .Q(\design_top.core0.REG2[5][3] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24015_ (.D(_04892_),
    .Q(\design_top.core0.REG2[5][4] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24016_ (.D(_04893_),
    .Q(\design_top.core0.REG2[5][5] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24017_ (.D(_04894_),
    .Q(\design_top.core0.REG2[5][6] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24018_ (.D(_04895_),
    .Q(\design_top.core0.REG2[5][7] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24019_ (.D(_04896_),
    .Q(\design_top.core0.REG2[5][8] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24020_ (.D(_04897_),
    .Q(\design_top.core0.REG2[5][9] ),
    .CLK(clknet_leaf_187_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24021_ (.D(_04898_),
    .Q(\design_top.core0.REG2[5][10] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24022_ (.D(_04899_),
    .Q(\design_top.core0.REG2[5][11] ),
    .CLK(clknet_leaf_302_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24023_ (.D(_04900_),
    .Q(\design_top.core0.REG2[5][12] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24024_ (.D(_04901_),
    .Q(\design_top.core0.REG2[5][13] ),
    .CLK(clknet_leaf_296_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24025_ (.D(_04902_),
    .Q(\design_top.core0.REG2[5][14] ),
    .CLK(clknet_leaf_302_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24026_ (.D(_04903_),
    .Q(\design_top.core0.REG2[5][15] ),
    .CLK(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24027_ (.D(_04904_),
    .Q(\design_top.core0.REG2[5][16] ),
    .CLK(clknet_leaf_300_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24028_ (.D(_04905_),
    .Q(\design_top.core0.REG2[5][17] ),
    .CLK(clknet_leaf_292_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24029_ (.D(_04906_),
    .Q(\design_top.core0.REG2[5][18] ),
    .CLK(clknet_leaf_295_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24030_ (.D(_04907_),
    .Q(\design_top.core0.REG2[5][19] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24031_ (.D(_04908_),
    .Q(\design_top.core0.REG2[5][20] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24032_ (.D(_04909_),
    .Q(\design_top.core0.REG2[5][21] ),
    .CLK(clknet_leaf_294_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24033_ (.D(_04910_),
    .Q(\design_top.core0.REG2[5][22] ),
    .CLK(clknet_leaf_270_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24034_ (.D(_04911_),
    .Q(\design_top.core0.REG2[5][23] ),
    .CLK(clknet_leaf_287_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24035_ (.D(_04912_),
    .Q(\design_top.core0.REG2[5][24] ),
    .CLK(clknet_leaf_287_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24036_ (.D(_04913_),
    .Q(\design_top.core0.REG2[5][25] ),
    .CLK(clknet_leaf_287_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24037_ (.D(_04914_),
    .Q(\design_top.core0.REG2[5][26] ),
    .CLK(clknet_leaf_287_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24038_ (.D(_04915_),
    .Q(\design_top.core0.REG2[5][27] ),
    .CLK(clknet_leaf_271_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24039_ (.D(_04916_),
    .Q(\design_top.core0.REG2[5][28] ),
    .CLK(clknet_leaf_268_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24040_ (.D(_04917_),
    .Q(\design_top.core0.REG2[5][29] ),
    .CLK(clknet_leaf_270_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24041_ (.D(_04918_),
    .Q(\design_top.core0.REG2[5][30] ),
    .CLK(clknet_leaf_272_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24042_ (.D(_04919_),
    .Q(\design_top.core0.REG2[5][31] ),
    .CLK(clknet_leaf_272_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24043_ (.D(_04920_),
    .Q(\design_top.core0.REG2[6][0] ),
    .CLK(clknet_leaf_292_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24044_ (.D(_04921_),
    .Q(\design_top.core0.REG2[6][1] ),
    .CLK(clknet_leaf_302_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24045_ (.D(_04922_),
    .Q(\design_top.core0.REG2[6][2] ),
    .CLK(clknet_leaf_302_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24046_ (.D(_04923_),
    .Q(\design_top.core0.REG2[6][3] ),
    .CLK(clknet_leaf_309_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24047_ (.D(_04924_),
    .Q(\design_top.core0.REG2[6][4] ),
    .CLK(clknet_leaf_310_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24048_ (.D(_04925_),
    .Q(\design_top.core0.REG2[6][5] ),
    .CLK(clknet_leaf_310_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24049_ (.D(_04926_),
    .Q(\design_top.core0.REG2[6][6] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24050_ (.D(_04927_),
    .Q(\design_top.core0.REG2[6][7] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24051_ (.D(_04928_),
    .Q(\design_top.core0.REG2[6][8] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24052_ (.D(_04929_),
    .Q(\design_top.core0.REG2[6][9] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24053_ (.D(_04930_),
    .Q(\design_top.core0.REG2[6][10] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24054_ (.D(_04931_),
    .Q(\design_top.core0.REG2[6][11] ),
    .CLK(clknet_leaf_301_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24055_ (.D(_04932_),
    .Q(\design_top.core0.REG2[6][12] ),
    .CLK(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24056_ (.D(_04933_),
    .Q(\design_top.core0.REG2[6][13] ),
    .CLK(clknet_leaf_296_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24057_ (.D(_04934_),
    .Q(\design_top.core0.REG2[6][14] ),
    .CLK(clknet_leaf_302_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24058_ (.D(_04935_),
    .Q(\design_top.core0.REG2[6][15] ),
    .CLK(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24059_ (.D(_04936_),
    .Q(\design_top.core0.REG2[6][16] ),
    .CLK(clknet_leaf_300_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24060_ (.D(_04937_),
    .Q(\design_top.core0.REG2[6][17] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24061_ (.D(_04938_),
    .Q(\design_top.core0.REG2[6][18] ),
    .CLK(clknet_leaf_294_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24062_ (.D(_04939_),
    .Q(\design_top.core0.REG2[6][19] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24063_ (.D(_04940_),
    .Q(\design_top.core0.REG2[6][20] ),
    .CLK(clknet_leaf_294_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24064_ (.D(_04941_),
    .Q(\design_top.core0.REG2[6][21] ),
    .CLK(clknet_leaf_294_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24065_ (.D(_04942_),
    .Q(\design_top.core0.REG2[6][22] ),
    .CLK(clknet_leaf_278_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24066_ (.D(_04943_),
    .Q(\design_top.core0.REG2[6][23] ),
    .CLK(clknet_leaf_278_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24067_ (.D(_04944_),
    .Q(\design_top.core0.REG2[6][24] ),
    .CLK(clknet_leaf_286_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24068_ (.D(_04945_),
    .Q(\design_top.core0.REG2[6][25] ),
    .CLK(clknet_leaf_278_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24069_ (.D(_04946_),
    .Q(\design_top.core0.REG2[6][26] ),
    .CLK(clknet_leaf_286_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24070_ (.D(_04947_),
    .Q(\design_top.core0.REG2[6][27] ),
    .CLK(clknet_leaf_271_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24071_ (.D(_04948_),
    .Q(\design_top.core0.REG2[6][28] ),
    .CLK(clknet_leaf_272_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24072_ (.D(_04949_),
    .Q(\design_top.core0.REG2[6][29] ),
    .CLK(clknet_leaf_271_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24073_ (.D(_04950_),
    .Q(\design_top.core0.REG2[6][30] ),
    .CLK(clknet_leaf_260_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24074_ (.D(_04951_),
    .Q(\design_top.core0.REG2[6][31] ),
    .CLK(clknet_leaf_272_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24075_ (.D(_04952_),
    .Q(\design_top.core0.REG2[7][0] ),
    .CLK(clknet_leaf_292_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24076_ (.D(_04953_),
    .Q(\design_top.core0.REG2[7][1] ),
    .CLK(clknet_leaf_302_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24077_ (.D(_04954_),
    .Q(\design_top.core0.REG2[7][2] ),
    .CLK(clknet_leaf_309_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24078_ (.D(_04955_),
    .Q(\design_top.core0.REG2[7][3] ),
    .CLK(clknet_leaf_310_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24079_ (.D(_04956_),
    .Q(\design_top.core0.REG2[7][4] ),
    .CLK(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24080_ (.D(_04957_),
    .Q(\design_top.core0.REG2[7][5] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24081_ (.D(_04958_),
    .Q(\design_top.core0.REG2[7][6] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24082_ (.D(_04959_),
    .Q(\design_top.core0.REG2[7][7] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24083_ (.D(_04960_),
    .Q(\design_top.core0.REG2[7][8] ),
    .CLK(clknet_leaf_187_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24084_ (.D(_04961_),
    .Q(\design_top.core0.REG2[7][9] ),
    .CLK(clknet_leaf_187_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24085_ (.D(_04962_),
    .Q(\design_top.core0.REG2[7][10] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24086_ (.D(_04963_),
    .Q(\design_top.core0.REG2[7][11] ),
    .CLK(clknet_leaf_300_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24087_ (.D(_04964_),
    .Q(\design_top.core0.REG2[7][12] ),
    .CLK(clknet_leaf_300_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24088_ (.D(_04965_),
    .Q(\design_top.core0.REG2[7][13] ),
    .CLK(clknet_leaf_292_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24089_ (.D(_04966_),
    .Q(\design_top.core0.REG2[7][14] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24090_ (.D(_04967_),
    .Q(\design_top.core0.REG2[7][15] ),
    .CLK(clknet_leaf_292_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24091_ (.D(_04968_),
    .Q(\design_top.core0.REG2[7][16] ),
    .CLK(clknet_leaf_300_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24092_ (.D(_04969_),
    .Q(\design_top.core0.REG2[7][17] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24093_ (.D(_04970_),
    .Q(\design_top.core0.REG2[7][18] ),
    .CLK(clknet_leaf_294_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24094_ (.D(_04971_),
    .Q(\design_top.core0.REG2[7][19] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24095_ (.D(_04972_),
    .Q(\design_top.core0.REG2[7][20] ),
    .CLK(clknet_leaf_287_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24096_ (.D(_04973_),
    .Q(\design_top.core0.REG2[7][21] ),
    .CLK(clknet_leaf_294_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24097_ (.D(_04974_),
    .Q(\design_top.core0.REG2[7][22] ),
    .CLK(clknet_leaf_270_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24098_ (.D(_04975_),
    .Q(\design_top.core0.REG2[7][23] ),
    .CLK(clknet_leaf_287_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24099_ (.D(_04976_),
    .Q(\design_top.core0.REG2[7][24] ),
    .CLK(clknet_leaf_286_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24100_ (.D(_04977_),
    .Q(\design_top.core0.REG2[7][25] ),
    .CLK(clknet_leaf_278_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24101_ (.D(_04978_),
    .Q(\design_top.core0.REG2[7][26] ),
    .CLK(clknet_leaf_286_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24102_ (.D(_04979_),
    .Q(\design_top.core0.REG2[7][27] ),
    .CLK(clknet_leaf_271_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24103_ (.D(_04980_),
    .Q(\design_top.core0.REG2[7][28] ),
    .CLK(clknet_leaf_272_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24104_ (.D(_04981_),
    .Q(\design_top.core0.REG2[7][29] ),
    .CLK(clknet_leaf_270_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24105_ (.D(_04982_),
    .Q(\design_top.core0.REG2[7][30] ),
    .CLK(clknet_leaf_260_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24106_ (.D(_04983_),
    .Q(\design_top.core0.REG2[7][31] ),
    .CLK(clknet_leaf_271_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24107_ (.D(_04984_),
    .Q(\design_top.core0.REG2[8][0] ),
    .CLK(clknet_leaf_296_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24108_ (.D(_04985_),
    .Q(\design_top.core0.REG2[8][1] ),
    .CLK(clknet_leaf_302_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24109_ (.D(_04986_),
    .Q(\design_top.core0.REG2[8][2] ),
    .CLK(clknet_leaf_302_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24110_ (.D(_04987_),
    .Q(\design_top.core0.REG2[8][3] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24111_ (.D(_04988_),
    .Q(\design_top.core0.REG2[8][4] ),
    .CLK(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24112_ (.D(_04989_),
    .Q(\design_top.core0.REG2[8][5] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24113_ (.D(_04990_),
    .Q(\design_top.core0.REG2[8][6] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24114_ (.D(_04991_),
    .Q(\design_top.core0.REG2[8][7] ),
    .CLK(clknet_leaf_187_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24115_ (.D(_04992_),
    .Q(\design_top.core0.REG2[8][8] ),
    .CLK(clknet_leaf_187_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24116_ (.D(_04993_),
    .Q(\design_top.core0.REG2[8][9] ),
    .CLK(clknet_leaf_187_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24117_ (.D(_04994_),
    .Q(\design_top.core0.REG2[8][10] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24118_ (.D(_04995_),
    .Q(\design_top.core0.REG2[8][11] ),
    .CLK(clknet_leaf_301_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24119_ (.D(_04996_),
    .Q(\design_top.core0.REG2[8][12] ),
    .CLK(clknet_leaf_300_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24120_ (.D(_04997_),
    .Q(\design_top.core0.REG2[8][13] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24121_ (.D(_04998_),
    .Q(\design_top.core0.REG2[8][14] ),
    .CLK(clknet_leaf_301_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24122_ (.D(_04999_),
    .Q(\design_top.core0.REG2[8][15] ),
    .CLK(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24123_ (.D(_05000_),
    .Q(\design_top.core0.REG2[8][16] ),
    .CLK(clknet_leaf_300_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24124_ (.D(_05001_),
    .Q(\design_top.core0.REG2[8][17] ),
    .CLK(clknet_leaf_295_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24125_ (.D(_05002_),
    .Q(\design_top.core0.REG2[8][18] ),
    .CLK(clknet_leaf_295_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24126_ (.D(_05003_),
    .Q(\design_top.core0.REG2[8][19] ),
    .CLK(clknet_leaf_295_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24127_ (.D(_05004_),
    .Q(\design_top.core0.REG2[8][20] ),
    .CLK(clknet_leaf_294_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24128_ (.D(_05005_),
    .Q(\design_top.core0.REG2[8][21] ),
    .CLK(clknet_leaf_270_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24129_ (.D(_05006_),
    .Q(\design_top.core0.REG2[8][22] ),
    .CLK(clknet_leaf_278_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24130_ (.D(_05007_),
    .Q(\design_top.core0.REG2[8][23] ),
    .CLK(clknet_leaf_278_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24131_ (.D(_05008_),
    .Q(\design_top.core0.REG2[8][24] ),
    .CLK(clknet_leaf_286_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24132_ (.D(_05009_),
    .Q(\design_top.core0.REG2[8][25] ),
    .CLK(clknet_leaf_278_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24133_ (.D(_05010_),
    .Q(\design_top.core0.REG2[8][26] ),
    .CLK(clknet_leaf_286_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24134_ (.D(_05011_),
    .Q(\design_top.core0.REG2[8][27] ),
    .CLK(clknet_leaf_271_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24135_ (.D(_05012_),
    .Q(\design_top.core0.REG2[8][28] ),
    .CLK(clknet_leaf_272_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24136_ (.D(_05013_),
    .Q(\design_top.core0.REG2[8][29] ),
    .CLK(clknet_leaf_271_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24137_ (.D(_05014_),
    .Q(\design_top.core0.REG2[8][30] ),
    .CLK(clknet_leaf_272_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24138_ (.D(_05015_),
    .Q(\design_top.core0.REG2[8][31] ),
    .CLK(clknet_leaf_271_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24139_ (.D(_05016_),
    .Q(\design_top.core0.REG2[0][0] ),
    .CLK(clknet_leaf_298_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24140_ (.D(_05017_),
    .Q(\design_top.core0.REG2[0][1] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24141_ (.D(_05018_),
    .Q(\design_top.core0.REG2[0][2] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24142_ (.D(_05019_),
    .Q(\design_top.core0.REG2[0][3] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24143_ (.D(_05020_),
    .Q(\design_top.core0.REG2[0][4] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24144_ (.D(_05021_),
    .Q(\design_top.core0.REG2[0][5] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24145_ (.D(_05022_),
    .Q(\design_top.core0.REG2[0][6] ),
    .CLK(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24146_ (.D(_05023_),
    .Q(\design_top.core0.REG2[0][7] ),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24147_ (.D(_05024_),
    .Q(\design_top.core0.REG2[0][8] ),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24148_ (.D(_05025_),
    .Q(\design_top.core0.REG2[0][9] ),
    .CLK(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24149_ (.D(_05026_),
    .Q(\design_top.core0.REG2[0][10] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24150_ (.D(_05027_),
    .Q(\design_top.core0.REG2[0][11] ),
    .CLK(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24151_ (.D(_05028_),
    .Q(\design_top.core0.REG2[0][12] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24152_ (.D(_05029_),
    .Q(\design_top.core0.REG2[0][13] ),
    .CLK(clknet_leaf_298_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24153_ (.D(_05030_),
    .Q(\design_top.core0.REG2[0][14] ),
    .CLK(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24154_ (.D(_05031_),
    .Q(\design_top.core0.REG2[0][15] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24155_ (.D(_05032_),
    .Q(\design_top.core0.REG2[0][16] ),
    .CLK(clknet_leaf_266_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24156_ (.D(_05033_),
    .Q(\design_top.core0.REG2[0][17] ),
    .CLK(clknet_leaf_266_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24157_ (.D(_05034_),
    .Q(\design_top.core0.REG2[0][18] ),
    .CLK(clknet_leaf_266_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24158_ (.D(_05035_),
    .Q(\design_top.core0.REG2[0][19] ),
    .CLK(clknet_leaf_266_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24159_ (.D(_05036_),
    .Q(\design_top.core0.REG2[0][20] ),
    .CLK(clknet_leaf_260_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24160_ (.D(_05037_),
    .Q(\design_top.core0.REG2[0][21] ),
    .CLK(clknet_leaf_260_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24161_ (.D(_05038_),
    .Q(\design_top.core0.REG2[0][22] ),
    .CLK(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24162_ (.D(_05039_),
    .Q(\design_top.core0.REG2[0][23] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24163_ (.D(_05040_),
    .Q(\design_top.core0.REG2[0][24] ),
    .CLK(clknet_leaf_281_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24164_ (.D(_05041_),
    .Q(\design_top.core0.REG2[0][25] ),
    .CLK(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24165_ (.D(_05042_),
    .Q(\design_top.core0.REG2[0][26] ),
    .CLK(clknet_leaf_282_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24166_ (.D(_05043_),
    .Q(\design_top.core0.REG2[0][27] ),
    .CLK(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24167_ (.D(_05044_),
    .Q(\design_top.core0.REG2[0][28] ),
    .CLK(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24168_ (.D(_05045_),
    .Q(\design_top.core0.REG2[0][29] ),
    .CLK(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24169_ (.D(_05046_),
    .Q(\design_top.core0.REG2[0][30] ),
    .CLK(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24170_ (.D(_05047_),
    .Q(\design_top.core0.REG2[0][31] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24171_ (.D(_05048_),
    .Q(\design_top.core0.REG2[10][0] ),
    .CLK(clknet_leaf_296_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24172_ (.D(_05049_),
    .Q(\design_top.core0.REG2[10][1] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24173_ (.D(_05050_),
    .Q(\design_top.core0.REG2[10][2] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24174_ (.D(_05051_),
    .Q(\design_top.core0.REG2[10][3] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24175_ (.D(_05052_),
    .Q(\design_top.core0.REG2[10][4] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24176_ (.D(_05053_),
    .Q(\design_top.core0.REG2[10][5] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24177_ (.D(_05054_),
    .Q(\design_top.core0.REG2[10][6] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24178_ (.D(_05055_),
    .Q(\design_top.core0.REG2[10][7] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24179_ (.D(_05056_),
    .Q(\design_top.core0.REG2[10][8] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24180_ (.D(_05057_),
    .Q(\design_top.core0.REG2[10][9] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24181_ (.D(_05058_),
    .Q(\design_top.core0.REG2[10][10] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24182_ (.D(_05059_),
    .Q(\design_top.core0.REG2[10][11] ),
    .CLK(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24183_ (.D(_05060_),
    .Q(\design_top.core0.REG2[10][12] ),
    .CLK(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24184_ (.D(_05061_),
    .Q(\design_top.core0.REG2[10][13] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24185_ (.D(_05062_),
    .Q(\design_top.core0.REG2[10][14] ),
    .CLK(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24186_ (.D(_05063_),
    .Q(\design_top.core0.REG2[10][15] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24187_ (.D(_05064_),
    .Q(\design_top.core0.REG2[10][16] ),
    .CLK(clknet_leaf_298_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24188_ (.D(_05065_),
    .Q(\design_top.core0.REG2[10][17] ),
    .CLK(clknet_leaf_269_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24189_ (.D(_05066_),
    .Q(\design_top.core0.REG2[10][18] ),
    .CLK(clknet_leaf_269_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24190_ (.D(_05067_),
    .Q(\design_top.core0.REG2[10][19] ),
    .CLK(clknet_leaf_269_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24191_ (.D(_05068_),
    .Q(\design_top.core0.REG2[10][20] ),
    .CLK(clknet_leaf_270_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24192_ (.D(_05069_),
    .Q(\design_top.core0.REG2[10][21] ),
    .CLK(clknet_leaf_269_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24193_ (.D(_05070_),
    .Q(\design_top.core0.REG2[10][22] ),
    .CLK(clknet_leaf_277_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24194_ (.D(_05071_),
    .Q(\design_top.core0.REG2[10][23] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24195_ (.D(_05072_),
    .Q(\design_top.core0.REG2[10][24] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24196_ (.D(_05073_),
    .Q(\design_top.core0.REG2[10][25] ),
    .CLK(clknet_leaf_277_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24197_ (.D(_05074_),
    .Q(\design_top.core0.REG2[10][26] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24198_ (.D(_05075_),
    .Q(\design_top.core0.REG2[10][27] ),
    .CLK(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24199_ (.D(_05076_),
    .Q(\design_top.core0.REG2[10][28] ),
    .CLK(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24200_ (.D(_05077_),
    .Q(\design_top.core0.REG2[10][29] ),
    .CLK(clknet_leaf_277_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24201_ (.D(_05078_),
    .Q(\design_top.core0.REG2[10][30] ),
    .CLK(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24202_ (.D(_05079_),
    .Q(\design_top.core0.REG2[10][31] ),
    .CLK(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24203_ (.D(_05080_),
    .Q(\design_top.core0.REG2[11][0] ),
    .CLK(clknet_leaf_296_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24204_ (.D(_05081_),
    .Q(\design_top.core0.REG2[11][1] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24205_ (.D(_05082_),
    .Q(\design_top.core0.REG2[11][2] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24206_ (.D(_05083_),
    .Q(\design_top.core0.REG2[11][3] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24207_ (.D(_05084_),
    .Q(\design_top.core0.REG2[11][4] ),
    .CLK(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24208_ (.D(_05085_),
    .Q(\design_top.core0.REG2[11][5] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24209_ (.D(_05086_),
    .Q(\design_top.core0.REG2[11][6] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24210_ (.D(_05087_),
    .Q(\design_top.core0.REG2[11][7] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24211_ (.D(_05088_),
    .Q(\design_top.core0.REG2[11][8] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24212_ (.D(_05089_),
    .Q(\design_top.core0.REG2[11][9] ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24213_ (.D(_05090_),
    .Q(\design_top.core0.REG2[11][10] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24214_ (.D(_05091_),
    .Q(\design_top.core0.REG2[11][11] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24215_ (.D(_05092_),
    .Q(\design_top.core0.REG2[11][12] ),
    .CLK(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24216_ (.D(_05093_),
    .Q(\design_top.core0.REG2[11][13] ),
    .CLK(clknet_leaf_295_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24217_ (.D(_05094_),
    .Q(\design_top.core0.REG2[11][14] ),
    .CLK(clknet_leaf_301_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24218_ (.D(_05095_),
    .Q(\design_top.core0.REG2[11][15] ),
    .CLK(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24219_ (.D(_05096_),
    .Q(\design_top.core0.REG2[11][16] ),
    .CLK(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24220_ (.D(_05097_),
    .Q(\design_top.core0.REG2[11][17] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24221_ (.D(_05098_),
    .Q(\design_top.core0.REG2[11][18] ),
    .CLK(clknet_leaf_295_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24222_ (.D(_05099_),
    .Q(\design_top.core0.REG2[11][19] ),
    .CLK(clknet_leaf_269_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24223_ (.D(_05100_),
    .Q(\design_top.core0.REG2[11][20] ),
    .CLK(clknet_leaf_269_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24224_ (.D(_05101_),
    .Q(\design_top.core0.REG2[11][21] ),
    .CLK(clknet_leaf_269_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24225_ (.D(_05102_),
    .Q(\design_top.core0.REG2[11][22] ),
    .CLK(clknet_leaf_277_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24226_ (.D(_05103_),
    .Q(\design_top.core0.REG2[11][23] ),
    .CLK(clknet_leaf_278_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24227_ (.D(_05104_),
    .Q(\design_top.core0.REG2[11][24] ),
    .CLK(clknet_leaf_286_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24228_ (.D(_05105_),
    .Q(\design_top.core0.REG2[11][25] ),
    .CLK(clknet_leaf_277_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24229_ (.D(_05106_),
    .Q(\design_top.core0.REG2[11][26] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24230_ (.D(_05107_),
    .Q(\design_top.core0.REG2[11][27] ),
    .CLK(clknet_leaf_271_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24231_ (.D(_05108_),
    .Q(\design_top.core0.REG2[11][28] ),
    .CLK(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24232_ (.D(_05109_),
    .Q(\design_top.core0.REG2[11][29] ),
    .CLK(clknet_leaf_271_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24233_ (.D(_05110_),
    .Q(\design_top.core0.REG2[11][30] ),
    .CLK(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24234_ (.D(_05111_),
    .Q(\design_top.core0.REG2[11][31] ),
    .CLK(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24235_ (.D(_05112_),
    .Q(\design_top.core0.REG2[12][0] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24236_ (.D(_05113_),
    .Q(\design_top.core0.REG2[12][1] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24237_ (.D(_05114_),
    .Q(\design_top.core0.REG2[12][2] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24238_ (.D(_05115_),
    .Q(\design_top.core0.REG2[12][3] ),
    .CLK(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24239_ (.D(_05116_),
    .Q(\design_top.core0.REG2[12][4] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24240_ (.D(_05117_),
    .Q(\design_top.core0.REG2[12][5] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24241_ (.D(_05118_),
    .Q(\design_top.core0.REG2[12][6] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24242_ (.D(_05119_),
    .Q(\design_top.core0.REG2[12][7] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24243_ (.D(_05120_),
    .Q(\design_top.core0.REG2[12][8] ),
    .CLK(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24244_ (.D(_05121_),
    .Q(\design_top.core0.REG2[12][9] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24245_ (.D(_05122_),
    .Q(\design_top.core0.REG2[12][10] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24246_ (.D(_05123_),
    .Q(\design_top.core0.REG2[12][11] ),
    .CLK(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24247_ (.D(_05124_),
    .Q(\design_top.core0.REG2[12][12] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24248_ (.D(_05125_),
    .Q(\design_top.core0.REG2[12][13] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24249_ (.D(_05126_),
    .Q(\design_top.core0.REG2[12][14] ),
    .CLK(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24250_ (.D(_05127_),
    .Q(\design_top.core0.REG2[12][15] ),
    .CLK(clknet_leaf_298_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24251_ (.D(_05128_),
    .Q(\design_top.core0.REG2[12][16] ),
    .CLK(clknet_leaf_298_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24252_ (.D(_05129_),
    .Q(\design_top.core0.REG2[12][17] ),
    .CLK(clknet_leaf_267_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24253_ (.D(_05130_),
    .Q(\design_top.core0.REG2[12][18] ),
    .CLK(clknet_leaf_267_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24254_ (.D(_05131_),
    .Q(\design_top.core0.REG2[12][19] ),
    .CLK(clknet_leaf_268_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24255_ (.D(_05132_),
    .Q(\design_top.core0.REG2[12][20] ),
    .CLK(clknet_leaf_269_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24256_ (.D(_05133_),
    .Q(\design_top.core0.REG2[12][21] ),
    .CLK(clknet_leaf_268_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24257_ (.D(_05134_),
    .Q(\design_top.core0.REG2[12][22] ),
    .CLK(clknet_leaf_277_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24258_ (.D(_05135_),
    .Q(\design_top.core0.REG2[12][23] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24259_ (.D(_05136_),
    .Q(\design_top.core0.REG2[12][24] ),
    .CLK(clknet_leaf_281_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24260_ (.D(_05137_),
    .Q(\design_top.core0.REG2[12][25] ),
    .CLK(clknet_leaf_277_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24261_ (.D(_05138_),
    .Q(\design_top.core0.REG2[12][26] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24262_ (.D(_05139_),
    .Q(\design_top.core0.REG2[12][27] ),
    .CLK(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24263_ (.D(_05140_),
    .Q(\design_top.core0.REG2[12][28] ),
    .CLK(clknet_leaf_258_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24264_ (.D(_05141_),
    .Q(\design_top.core0.REG2[12][29] ),
    .CLK(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24265_ (.D(_05142_),
    .Q(\design_top.core0.REG2[12][30] ),
    .CLK(clknet_leaf_258_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24266_ (.D(_05143_),
    .Q(\design_top.core0.REG2[12][31] ),
    .CLK(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24267_ (.D(_05144_),
    .Q(\design_top.core0.REG2[13][0] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24268_ (.D(_05145_),
    .Q(\design_top.core0.REG2[13][1] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24269_ (.D(_05146_),
    .Q(\design_top.core0.REG2[13][2] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24270_ (.D(_05147_),
    .Q(\design_top.core0.REG2[13][3] ),
    .CLK(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24271_ (.D(_05148_),
    .Q(\design_top.core0.REG2[13][4] ),
    .CLK(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24272_ (.D(_05149_),
    .Q(\design_top.core0.REG2[13][5] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24273_ (.D(_05150_),
    .Q(\design_top.core0.REG2[13][6] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24274_ (.D(_05151_),
    .Q(\design_top.core0.REG2[13][7] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24275_ (.D(_05152_),
    .Q(\design_top.core0.REG2[13][8] ),
    .CLK(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24276_ (.D(_05153_),
    .Q(\design_top.core0.REG2[13][9] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24277_ (.D(_05154_),
    .Q(\design_top.core0.REG2[13][10] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24278_ (.D(_05155_),
    .Q(\design_top.core0.REG2[13][11] ),
    .CLK(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24279_ (.D(_05156_),
    .Q(\design_top.core0.REG2[13][12] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24280_ (.D(_05157_),
    .Q(\design_top.core0.REG2[13][13] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24281_ (.D(_05158_),
    .Q(\design_top.core0.REG2[13][14] ),
    .CLK(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24282_ (.D(_05159_),
    .Q(\design_top.core0.REG2[13][15] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24283_ (.D(_05160_),
    .Q(\design_top.core0.REG2[13][16] ),
    .CLK(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24284_ (.D(_05161_),
    .Q(\design_top.core0.REG2[13][17] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24285_ (.D(_05162_),
    .Q(\design_top.core0.REG2[13][18] ),
    .CLK(clknet_leaf_267_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24286_ (.D(_05163_),
    .Q(\design_top.core0.REG2[13][19] ),
    .CLK(clknet_leaf_267_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24287_ (.D(_05164_),
    .Q(\design_top.core0.REG2[13][20] ),
    .CLK(clknet_leaf_269_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24288_ (.D(_05165_),
    .Q(\design_top.core0.REG2[13][21] ),
    .CLK(clknet_leaf_268_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24289_ (.D(_05166_),
    .Q(\design_top.core0.REG2[13][22] ),
    .CLK(clknet_leaf_277_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24290_ (.D(_05167_),
    .Q(\design_top.core0.REG2[13][23] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24291_ (.D(_05168_),
    .Q(\design_top.core0.REG2[13][24] ),
    .CLK(clknet_leaf_281_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24292_ (.D(_05169_),
    .Q(\design_top.core0.REG2[13][25] ),
    .CLK(clknet_leaf_277_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24293_ (.D(_05170_),
    .Q(\design_top.core0.REG2[13][26] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24294_ (.D(_05171_),
    .Q(\design_top.core0.REG2[13][27] ),
    .CLK(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24295_ (.D(_05172_),
    .Q(\design_top.core0.REG2[13][28] ),
    .CLK(clknet_leaf_258_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24296_ (.D(_05173_),
    .Q(\design_top.core0.REG2[13][29] ),
    .CLK(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24297_ (.D(_05174_),
    .Q(\design_top.core0.REG2[13][30] ),
    .CLK(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24298_ (.D(_05175_),
    .Q(\design_top.core0.REG2[13][31] ),
    .CLK(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24299_ (.D(_05176_),
    .Q(\design_top.core0.REG2[14][0] ),
    .CLK(clknet_leaf_298_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24300_ (.D(_05177_),
    .Q(\design_top.core0.REG2[14][1] ),
    .CLK(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24301_ (.D(_05178_),
    .Q(\design_top.core0.REG2[14][2] ),
    .CLK(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24302_ (.D(_05179_),
    .Q(\design_top.core0.REG2[14][3] ),
    .CLK(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24303_ (.D(_05180_),
    .Q(\design_top.core0.REG2[14][4] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24304_ (.D(_05181_),
    .Q(\design_top.core0.REG2[14][5] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24305_ (.D(_05182_),
    .Q(\design_top.core0.REG2[14][6] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24306_ (.D(_05183_),
    .Q(\design_top.core0.REG2[14][7] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24307_ (.D(_05184_),
    .Q(\design_top.core0.REG2[14][8] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24308_ (.D(_05185_),
    .Q(\design_top.core0.REG2[14][9] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24309_ (.D(_05186_),
    .Q(\design_top.core0.REG2[14][10] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24310_ (.D(_05187_),
    .Q(\design_top.core0.REG2[14][11] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24311_ (.D(_05188_),
    .Q(\design_top.core0.REG2[14][12] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24312_ (.D(_05189_),
    .Q(\design_top.core0.REG2[14][13] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24313_ (.D(_05190_),
    .Q(\design_top.core0.REG2[14][14] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24314_ (.D(_05191_),
    .Q(\design_top.core0.REG2[14][15] ),
    .CLK(clknet_leaf_298_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24315_ (.D(_05192_),
    .Q(\design_top.core0.REG2[14][16] ),
    .CLK(clknet_leaf_298_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24316_ (.D(_05193_),
    .Q(\design_top.core0.REG2[14][17] ),
    .CLK(clknet_leaf_269_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24317_ (.D(_05194_),
    .Q(\design_top.core0.REG2[14][18] ),
    .CLK(clknet_leaf_267_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24318_ (.D(_05195_),
    .Q(\design_top.core0.REG2[14][19] ),
    .CLK(clknet_leaf_267_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24319_ (.D(_05196_),
    .Q(\design_top.core0.REG2[14][20] ),
    .CLK(clknet_leaf_271_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24320_ (.D(_05197_),
    .Q(\design_top.core0.REG2[14][21] ),
    .CLK(clknet_leaf_272_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24321_ (.D(_05198_),
    .Q(\design_top.core0.REG2[14][22] ),
    .CLK(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24322_ (.D(_05199_),
    .Q(\design_top.core0.REG2[14][23] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24323_ (.D(_05200_),
    .Q(\design_top.core0.REG2[14][24] ),
    .CLK(clknet_leaf_281_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24324_ (.D(_05201_),
    .Q(\design_top.core0.REG2[14][25] ),
    .CLK(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24325_ (.D(_05202_),
    .Q(\design_top.core0.REG2[14][26] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24326_ (.D(_05203_),
    .Q(\design_top.core0.REG2[14][27] ),
    .CLK(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24327_ (.D(_05204_),
    .Q(\design_top.core0.REG2[14][28] ),
    .CLK(clknet_leaf_259_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24328_ (.D(_05205_),
    .Q(\design_top.core0.REG2[14][29] ),
    .CLK(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24329_ (.D(_05206_),
    .Q(\design_top.core0.REG2[14][30] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24330_ (.D(_05207_),
    .Q(\design_top.core0.REG2[14][31] ),
    .CLK(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24331_ (.D(_05208_),
    .Q(\design_top.MEM[8][0] ),
    .CLK(clknet_leaf_37_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24332_ (.D(_05209_),
    .Q(\design_top.MEM[8][1] ),
    .CLK(clknet_leaf_37_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24333_ (.D(_05210_),
    .Q(\design_top.MEM[8][2] ),
    .CLK(clknet_leaf_37_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24334_ (.D(_05211_),
    .Q(\design_top.MEM[8][3] ),
    .CLK(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24335_ (.D(_05212_),
    .Q(\design_top.MEM[8][4] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24336_ (.D(_05213_),
    .Q(\design_top.MEM[8][5] ),
    .CLK(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24337_ (.D(_05214_),
    .Q(\design_top.MEM[8][6] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24338_ (.D(_05215_),
    .Q(\design_top.MEM[8][7] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24339_ (.D(_05216_),
    .Q(\design_top.MEM[9][0] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24340_ (.D(_05217_),
    .Q(\design_top.MEM[9][1] ),
    .CLK(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24341_ (.D(_05218_),
    .Q(\design_top.MEM[9][2] ),
    .CLK(clknet_leaf_37_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24342_ (.D(_05219_),
    .Q(\design_top.MEM[9][3] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24343_ (.D(_05220_),
    .Q(\design_top.MEM[9][4] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24344_ (.D(_05221_),
    .Q(\design_top.MEM[9][5] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24345_ (.D(_05222_),
    .Q(\design_top.MEM[9][6] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24346_ (.D(_05223_),
    .Q(\design_top.MEM[9][7] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24347_ (.D(_05224_),
    .Q(\design_top.MEM[26][0] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24348_ (.D(_05225_),
    .Q(\design_top.MEM[26][1] ),
    .CLK(clknet_leaf_435_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24349_ (.D(_05226_),
    .Q(\design_top.MEM[26][2] ),
    .CLK(clknet_leaf_434_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24350_ (.D(_05227_),
    .Q(\design_top.MEM[26][3] ),
    .CLK(clknet_leaf_438_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24351_ (.D(_05228_),
    .Q(\design_top.MEM[26][4] ),
    .CLK(clknet_leaf_438_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24352_ (.D(_05229_),
    .Q(\design_top.MEM[26][5] ),
    .CLK(clknet_leaf_441_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24353_ (.D(_05230_),
    .Q(\design_top.MEM[26][6] ),
    .CLK(clknet_leaf_442_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24354_ (.D(_05231_),
    .Q(\design_top.MEM[26][7] ),
    .CLK(clknet_leaf_442_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24355_ (.D(_05232_),
    .Q(\design_top.MEM[25][0] ),
    .CLK(clknet_leaf_434_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24356_ (.D(_05233_),
    .Q(\design_top.MEM[25][1] ),
    .CLK(clknet_leaf_435_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24357_ (.D(_05234_),
    .Q(\design_top.MEM[25][2] ),
    .CLK(clknet_leaf_434_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24358_ (.D(_05235_),
    .Q(\design_top.MEM[25][3] ),
    .CLK(clknet_leaf_438_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24359_ (.D(_05236_),
    .Q(\design_top.MEM[25][4] ),
    .CLK(clknet_leaf_438_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24360_ (.D(_05237_),
    .Q(\design_top.MEM[25][5] ),
    .CLK(clknet_leaf_441_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24361_ (.D(_05238_),
    .Q(\design_top.MEM[25][6] ),
    .CLK(clknet_leaf_441_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24362_ (.D(_05239_),
    .Q(\design_top.MEM[25][7] ),
    .CLK(clknet_leaf_441_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24363_ (.D(_05240_),
    .Q(\design_top.MEM[38][0] ),
    .CLK(clknet_leaf_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24364_ (.D(_05241_),
    .Q(\design_top.MEM[38][1] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24365_ (.D(_05242_),
    .Q(\design_top.MEM[38][2] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24366_ (.D(_05243_),
    .Q(\design_top.MEM[38][3] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24367_ (.D(_05244_),
    .Q(\design_top.MEM[38][4] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24368_ (.D(_05245_),
    .Q(\design_top.MEM[38][5] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24369_ (.D(_05246_),
    .Q(\design_top.MEM[38][6] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24370_ (.D(_05247_),
    .Q(\design_top.MEM[38][7] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24371_ (.D(_05248_),
    .Q(\design_top.MEM[24][0] ),
    .CLK(clknet_leaf_433_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24372_ (.D(_05249_),
    .Q(\design_top.MEM[24][1] ),
    .CLK(clknet_leaf_435_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24373_ (.D(_05250_),
    .Q(\design_top.MEM[24][2] ),
    .CLK(clknet_leaf_434_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24374_ (.D(_05251_),
    .Q(\design_top.MEM[24][3] ),
    .CLK(clknet_leaf_439_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24375_ (.D(_05252_),
    .Q(\design_top.MEM[24][4] ),
    .CLK(clknet_leaf_439_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24376_ (.D(_05253_),
    .Q(\design_top.MEM[24][5] ),
    .CLK(clknet_leaf_441_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24377_ (.D(_05254_),
    .Q(\design_top.MEM[24][6] ),
    .CLK(clknet_leaf_440_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24378_ (.D(_05255_),
    .Q(\design_top.MEM[24][7] ),
    .CLK(clknet_leaf_425_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24379_ (.D(_05256_),
    .Q(\design_top.MEM[37][0] ),
    .CLK(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24380_ (.D(_05257_),
    .Q(\design_top.MEM[37][1] ),
    .CLK(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24381_ (.D(_05258_),
    .Q(\design_top.MEM[37][2] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24382_ (.D(_05259_),
    .Q(\design_top.MEM[37][3] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24383_ (.D(_05260_),
    .Q(\design_top.MEM[37][4] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24384_ (.D(_05261_),
    .Q(\design_top.MEM[37][5] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24385_ (.D(_05262_),
    .Q(\design_top.MEM[37][6] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24386_ (.D(_05263_),
    .Q(\design_top.MEM[37][7] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24387_ (.D(_05264_),
    .Q(\design_top.MEM[23][0] ),
    .CLK(clknet_leaf_433_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24388_ (.D(_05265_),
    .Q(\design_top.MEM[23][1] ),
    .CLK(clknet_leaf_439_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24389_ (.D(_05266_),
    .Q(\design_top.MEM[23][2] ),
    .CLK(clknet_leaf_432_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24390_ (.D(_05267_),
    .Q(\design_top.MEM[23][3] ),
    .CLK(clknet_leaf_439_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24391_ (.D(_05268_),
    .Q(\design_top.MEM[23][4] ),
    .CLK(clknet_leaf_439_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24392_ (.D(_05269_),
    .Q(\design_top.MEM[23][5] ),
    .CLK(clknet_leaf_425_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24393_ (.D(_05270_),
    .Q(\design_top.MEM[23][6] ),
    .CLK(clknet_leaf_440_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24394_ (.D(_05271_),
    .Q(\design_top.MEM[23][7] ),
    .CLK(clknet_leaf_441_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24395_ (.D(_05272_),
    .Q(\design_top.MEM[45][0] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24396_ (.D(_05273_),
    .Q(\design_top.MEM[45][1] ),
    .CLK(clknet_leaf_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24397_ (.D(_05274_),
    .Q(\design_top.MEM[45][2] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24398_ (.D(_05275_),
    .Q(\design_top.MEM[45][3] ),
    .CLK(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24399_ (.D(_05276_),
    .Q(\design_top.MEM[45][4] ),
    .CLK(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24400_ (.D(_05277_),
    .Q(\design_top.MEM[45][5] ),
    .CLK(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24401_ (.D(_05278_),
    .Q(\design_top.MEM[45][6] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24402_ (.D(_05279_),
    .Q(\design_top.MEM[45][7] ),
    .CLK(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24403_ (.D(_05280_),
    .Q(\design_top.MEM[44][0] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24404_ (.D(_05281_),
    .Q(\design_top.MEM[44][1] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24405_ (.D(_05282_),
    .Q(\design_top.MEM[44][2] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24406_ (.D(_05283_),
    .Q(\design_top.MEM[44][3] ),
    .CLK(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24407_ (.D(_05284_),
    .Q(\design_top.MEM[44][4] ),
    .CLK(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24408_ (.D(_05285_),
    .Q(\design_top.MEM[44][5] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24409_ (.D(_05286_),
    .Q(\design_top.MEM[44][6] ),
    .CLK(clknet_leaf_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24410_ (.D(_05287_),
    .Q(\design_top.MEM[44][7] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24411_ (.D(_05288_),
    .Q(\design_top.MEM[50][0] ),
    .CLK(clknet_leaf_432_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24412_ (.D(_05289_),
    .Q(\design_top.MEM[50][1] ),
    .CLK(clknet_leaf_430_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24413_ (.D(_05290_),
    .Q(\design_top.MEM[50][2] ),
    .CLK(clknet_leaf_432_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24414_ (.D(_05291_),
    .Q(\design_top.MEM[50][3] ),
    .CLK(clknet_leaf_427_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24415_ (.D(_05292_),
    .Q(\design_top.MEM[50][4] ),
    .CLK(clknet_leaf_427_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24416_ (.D(_05293_),
    .Q(\design_top.MEM[50][5] ),
    .CLK(clknet_leaf_424_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24417_ (.D(_05294_),
    .Q(\design_top.MEM[50][6] ),
    .CLK(clknet_leaf_426_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24418_ (.D(_05295_),
    .Q(\design_top.MEM[50][7] ),
    .CLK(clknet_leaf_424_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24419_ (.D(_05296_),
    .Q(\design_top.MEM[43][0] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24420_ (.D(_05297_),
    .Q(\design_top.MEM[43][1] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24421_ (.D(_05298_),
    .Q(\design_top.MEM[43][2] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24422_ (.D(_05299_),
    .Q(\design_top.MEM[43][3] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24423_ (.D(_05300_),
    .Q(\design_top.MEM[43][4] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24424_ (.D(_05301_),
    .Q(\design_top.MEM[43][5] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24425_ (.D(_05302_),
    .Q(\design_top.MEM[43][6] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24426_ (.D(_05303_),
    .Q(\design_top.MEM[43][7] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24427_ (.D(_05304_),
    .Q(\design_top.MEM[4][0] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24428_ (.D(_05305_),
    .Q(\design_top.MEM[4][1] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24429_ (.D(_05306_),
    .Q(\design_top.MEM[4][2] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24430_ (.D(_05307_),
    .Q(\design_top.MEM[4][3] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24431_ (.D(_05308_),
    .Q(\design_top.MEM[4][4] ),
    .CLK(clknet_leaf_402_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24432_ (.D(_05309_),
    .Q(\design_top.MEM[4][5] ),
    .CLK(clknet_leaf_402_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24433_ (.D(_05310_),
    .Q(\design_top.MEM[4][6] ),
    .CLK(clknet_leaf_400_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24434_ (.D(_05311_),
    .Q(\design_top.MEM[4][7] ),
    .CLK(clknet_leaf_401_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24435_ (.D(_05312_),
    .Q(\design_top.MEM[42][0] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24436_ (.D(_05313_),
    .Q(\design_top.MEM[42][1] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24437_ (.D(_05314_),
    .Q(\design_top.MEM[42][2] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24438_ (.D(_05315_),
    .Q(\design_top.MEM[42][3] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24439_ (.D(_05316_),
    .Q(\design_top.MEM[42][4] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24440_ (.D(_05317_),
    .Q(\design_top.MEM[42][5] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24441_ (.D(_05318_),
    .Q(\design_top.MEM[42][6] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24442_ (.D(_05319_),
    .Q(\design_top.MEM[42][7] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24443_ (.D(_05320_),
    .Q(\design_top.MEM[49][0] ),
    .CLK(clknet_leaf_404_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24444_ (.D(_05321_),
    .Q(\design_top.MEM[49][1] ),
    .CLK(clknet_leaf_432_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24445_ (.D(_05322_),
    .Q(\design_top.MEM[49][2] ),
    .CLK(clknet_leaf_432_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24446_ (.D(_05323_),
    .Q(\design_top.MEM[49][3] ),
    .CLK(clknet_leaf_431_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24447_ (.D(_05324_),
    .Q(\design_top.MEM[49][4] ),
    .CLK(clknet_leaf_427_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24448_ (.D(_05325_),
    .Q(\design_top.MEM[49][5] ),
    .CLK(clknet_leaf_426_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24449_ (.D(_05326_),
    .Q(\design_top.MEM[49][6] ),
    .CLK(clknet_leaf_426_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24450_ (.D(_05327_),
    .Q(\design_top.MEM[49][7] ),
    .CLK(clknet_leaf_424_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24451_ (.D(_05328_),
    .Q(\design_top.MEM[41][0] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24452_ (.D(_05329_),
    .Q(\design_top.MEM[41][1] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24453_ (.D(_05330_),
    .Q(\design_top.MEM[41][2] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24454_ (.D(_05331_),
    .Q(\design_top.MEM[41][3] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24455_ (.D(_05332_),
    .Q(\design_top.MEM[41][4] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24456_ (.D(_05333_),
    .Q(\design_top.MEM[41][5] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24457_ (.D(_05334_),
    .Q(\design_top.MEM[41][6] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24458_ (.D(_05335_),
    .Q(\design_top.MEM[41][7] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24459_ (.D(_05336_),
    .Q(\design_top.MEM[48][0] ),
    .CLK(clknet_leaf_404_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24460_ (.D(_05337_),
    .Q(\design_top.MEM[48][1] ),
    .CLK(clknet_leaf_432_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24461_ (.D(_05338_),
    .Q(\design_top.MEM[48][2] ),
    .CLK(clknet_leaf_432_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24462_ (.D(_05339_),
    .Q(\design_top.MEM[48][3] ),
    .CLK(clknet_leaf_430_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24463_ (.D(_05340_),
    .Q(\design_top.MEM[48][4] ),
    .CLK(clknet_leaf_427_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24464_ (.D(_05341_),
    .Q(\design_top.MEM[48][5] ),
    .CLK(clknet_leaf_424_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24465_ (.D(_05342_),
    .Q(\design_top.MEM[48][6] ),
    .CLK(clknet_leaf_426_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24466_ (.D(_05343_),
    .Q(\design_top.MEM[48][7] ),
    .CLK(clknet_leaf_424_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24467_ (.D(_05344_),
    .Q(\design_top.MEM[40][0] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24468_ (.D(_05345_),
    .Q(\design_top.MEM[40][1] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24469_ (.D(_05346_),
    .Q(\design_top.MEM[40][2] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24470_ (.D(_05347_),
    .Q(\design_top.MEM[40][3] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24471_ (.D(_05348_),
    .Q(\design_top.MEM[40][4] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24472_ (.D(_05349_),
    .Q(\design_top.MEM[40][5] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24473_ (.D(_05350_),
    .Q(\design_top.MEM[40][6] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24474_ (.D(_05351_),
    .Q(\design_top.MEM[40][7] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24475_ (.D(_05352_),
    .Q(\design_top.MEM[3][0] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24476_ (.D(_05353_),
    .Q(\design_top.MEM[3][1] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24477_ (.D(_05354_),
    .Q(\design_top.MEM[3][2] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24478_ (.D(_05355_),
    .Q(\design_top.MEM[3][3] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24479_ (.D(_05356_),
    .Q(\design_top.MEM[3][4] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24480_ (.D(_05357_),
    .Q(\design_top.MEM[3][5] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24481_ (.D(_05358_),
    .Q(\design_top.MEM[3][6] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24482_ (.D(_05359_),
    .Q(\design_top.MEM[3][7] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24483_ (.D(_05360_),
    .Q(\design_top.MEM[47][0] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24484_ (.D(_05361_),
    .Q(\design_top.MEM[47][1] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24485_ (.D(_05362_),
    .Q(\design_top.MEM[47][2] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24486_ (.D(_05363_),
    .Q(\design_top.MEM[47][3] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24487_ (.D(_05364_),
    .Q(\design_top.MEM[47][4] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24488_ (.D(_05365_),
    .Q(\design_top.MEM[47][5] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24489_ (.D(_05366_),
    .Q(\design_top.MEM[47][6] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24490_ (.D(_05367_),
    .Q(\design_top.MEM[47][7] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24491_ (.D(_05368_),
    .Q(\design_top.MEM[46][0] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24492_ (.D(_05369_),
    .Q(\design_top.MEM[46][1] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24493_ (.D(_05370_),
    .Q(\design_top.MEM[46][2] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24494_ (.D(_05371_),
    .Q(\design_top.MEM[46][3] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24495_ (.D(_05372_),
    .Q(\design_top.MEM[46][4] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24496_ (.D(_05373_),
    .Q(\design_top.MEM[46][5] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24497_ (.D(_05374_),
    .Q(\design_top.MEM[46][6] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24498_ (.D(_05375_),
    .Q(\design_top.MEM[46][7] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24499_ (.D(_05376_),
    .Q(\design_top.MEM[39][0] ),
    .CLK(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24500_ (.D(_05377_),
    .Q(\design_top.MEM[39][1] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24501_ (.D(_05378_),
    .Q(\design_top.MEM[39][2] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24502_ (.D(_05379_),
    .Q(\design_top.MEM[39][3] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24503_ (.D(_05380_),
    .Q(\design_top.MEM[39][4] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24504_ (.D(_05381_),
    .Q(\design_top.MEM[39][5] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24505_ (.D(_05382_),
    .Q(\design_top.MEM[39][6] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24506_ (.D(_05383_),
    .Q(\design_top.MEM[39][7] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24507_ (.D(_05384_),
    .Q(\design_top.MEM[52][0] ),
    .CLK(clknet_leaf_404_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24508_ (.D(_05385_),
    .Q(\design_top.MEM[52][1] ),
    .CLK(clknet_leaf_405_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24509_ (.D(_05386_),
    .Q(\design_top.MEM[52][2] ),
    .CLK(clknet_leaf_405_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24510_ (.D(_05387_),
    .Q(\design_top.MEM[52][3] ),
    .CLK(clknet_leaf_430_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24511_ (.D(_05388_),
    .Q(\design_top.MEM[52][4] ),
    .CLK(clknet_leaf_428_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24512_ (.D(_05389_),
    .Q(\design_top.MEM[52][5] ),
    .CLK(clknet_leaf_423_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24513_ (.D(_05390_),
    .Q(\design_top.MEM[52][6] ),
    .CLK(clknet_leaf_428_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24514_ (.D(_05391_),
    .Q(\design_top.MEM[52][7] ),
    .CLK(clknet_leaf_423_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24515_ (.D(_05392_),
    .Q(\design_top.MEM[54][0] ),
    .CLK(clknet_leaf_404_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24516_ (.D(_05393_),
    .Q(\design_top.MEM[54][1] ),
    .CLK(clknet_leaf_430_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24517_ (.D(_05394_),
    .Q(\design_top.MEM[54][2] ),
    .CLK(clknet_leaf_404_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24518_ (.D(_05395_),
    .Q(\design_top.MEM[54][3] ),
    .CLK(clknet_leaf_428_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24519_ (.D(_05396_),
    .Q(\design_top.MEM[54][4] ),
    .CLK(clknet_leaf_428_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24520_ (.D(_05397_),
    .Q(\design_top.MEM[54][5] ),
    .CLK(clknet_leaf_423_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24521_ (.D(_05398_),
    .Q(\design_top.MEM[54][6] ),
    .CLK(clknet_leaf_428_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24522_ (.D(_05399_),
    .Q(\design_top.MEM[54][7] ),
    .CLK(clknet_leaf_423_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24523_ (.D(_05400_),
    .Q(\design_top.MEM[51][0] ),
    .CLK(clknet_leaf_404_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24524_ (.D(_05401_),
    .Q(\design_top.MEM[51][1] ),
    .CLK(clknet_leaf_430_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24525_ (.D(_05402_),
    .Q(\design_top.MEM[51][2] ),
    .CLK(clknet_leaf_404_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24526_ (.D(_05403_),
    .Q(\design_top.MEM[51][3] ),
    .CLK(clknet_leaf_427_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24527_ (.D(_05404_),
    .Q(\design_top.MEM[51][4] ),
    .CLK(clknet_leaf_428_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24528_ (.D(_05405_),
    .Q(\design_top.MEM[51][5] ),
    .CLK(clknet_leaf_423_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24529_ (.D(_05406_),
    .Q(\design_top.MEM[51][6] ),
    .CLK(clknet_leaf_426_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24530_ (.D(_05407_),
    .Q(\design_top.MEM[51][7] ),
    .CLK(clknet_leaf_424_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24531_ (.D(_05408_),
    .Q(\design_top.MEM[22][0] ),
    .CLK(clknet_leaf_433_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24532_ (.D(_05409_),
    .Q(\design_top.MEM[22][1] ),
    .CLK(clknet_leaf_431_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24533_ (.D(_05410_),
    .Q(\design_top.MEM[22][2] ),
    .CLK(clknet_leaf_432_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24534_ (.D(_05411_),
    .Q(\design_top.MEM[22][3] ),
    .CLK(clknet_leaf_427_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24535_ (.D(_05412_),
    .Q(\design_top.MEM[22][4] ),
    .CLK(clknet_leaf_426_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24536_ (.D(_05413_),
    .Q(\design_top.MEM[22][5] ),
    .CLK(clknet_leaf_424_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24537_ (.D(_05414_),
    .Q(\design_top.MEM[22][6] ),
    .CLK(clknet_leaf_426_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24538_ (.D(_05415_),
    .Q(\design_top.MEM[22][7] ),
    .CLK(clknet_leaf_425_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24539_ (.D(_05416_),
    .Q(\design_top.MEM[36][0] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24540_ (.D(_05417_),
    .Q(\design_top.MEM[36][1] ),
    .CLK(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24541_ (.D(_05418_),
    .Q(\design_top.MEM[36][2] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24542_ (.D(_05419_),
    .Q(\design_top.MEM[36][3] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24543_ (.D(_05420_),
    .Q(\design_top.MEM[36][4] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24544_ (.D(_05421_),
    .Q(\design_top.MEM[36][5] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24545_ (.D(_05422_),
    .Q(\design_top.MEM[36][6] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24546_ (.D(_05423_),
    .Q(\design_top.MEM[36][7] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24547_ (.D(_05424_),
    .Q(\design_top.MEM[21][0] ),
    .CLK(clknet_leaf_432_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24548_ (.D(_05425_),
    .Q(\design_top.MEM[21][1] ),
    .CLK(clknet_leaf_431_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24549_ (.D(_05426_),
    .Q(\design_top.MEM[21][2] ),
    .CLK(clknet_leaf_435_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24550_ (.D(_05427_),
    .Q(\design_top.MEM[21][3] ),
    .CLK(clknet_leaf_427_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24551_ (.D(_05428_),
    .Q(\design_top.MEM[21][4] ),
    .CLK(clknet_leaf_426_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24552_ (.D(_05429_),
    .Q(\design_top.MEM[21][5] ),
    .CLK(clknet_leaf_425_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24553_ (.D(_05430_),
    .Q(\design_top.MEM[21][6] ),
    .CLK(clknet_leaf_440_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24554_ (.D(_05431_),
    .Q(\design_top.MEM[21][7] ),
    .CLK(clknet_leaf_441_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24555_ (.D(_05432_),
    .Q(\design_top.MEM[20][0] ),
    .CLK(clknet_leaf_432_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24556_ (.D(_05433_),
    .Q(\design_top.MEM[20][1] ),
    .CLK(clknet_leaf_431_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24557_ (.D(_05434_),
    .Q(\design_top.MEM[20][2] ),
    .CLK(clknet_leaf_432_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24558_ (.D(_05435_),
    .Q(\design_top.MEM[20][3] ),
    .CLK(clknet_leaf_427_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24559_ (.D(_05436_),
    .Q(\design_top.MEM[20][4] ),
    .CLK(clknet_leaf_426_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24560_ (.D(_05437_),
    .Q(\design_top.MEM[20][5] ),
    .CLK(clknet_leaf_425_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24561_ (.D(_05438_),
    .Q(\design_top.MEM[20][6] ),
    .CLK(clknet_leaf_426_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24562_ (.D(_05439_),
    .Q(\design_top.MEM[20][7] ),
    .CLK(clknet_leaf_425_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24563_ (.D(_05440_),
    .Q(\design_top.MEM[1][0] ),
    .CLK(clknet_leaf_39_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24564_ (.D(_05441_),
    .Q(\design_top.MEM[1][1] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24565_ (.D(_05442_),
    .Q(\design_top.MEM[1][2] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24566_ (.D(_05443_),
    .Q(\design_top.MEM[1][3] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24567_ (.D(_05444_),
    .Q(\design_top.MEM[1][4] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24568_ (.D(_05445_),
    .Q(\design_top.MEM[1][5] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24569_ (.D(_05446_),
    .Q(\design_top.MEM[1][6] ),
    .CLK(clknet_leaf_39_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24570_ (.D(_05447_),
    .Q(\design_top.MEM[1][7] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24571_ (.D(_05448_),
    .Q(\design_top.MEM[35][0] ),
    .CLK(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24572_ (.D(_05449_),
    .Q(\design_top.MEM[35][1] ),
    .CLK(clknet_leaf_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24573_ (.D(_05450_),
    .Q(\design_top.MEM[35][2] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24574_ (.D(_05451_),
    .Q(\design_top.MEM[35][3] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24575_ (.D(_05452_),
    .Q(\design_top.MEM[35][4] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24576_ (.D(_05453_),
    .Q(\design_top.MEM[35][5] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24577_ (.D(_05454_),
    .Q(\design_top.MEM[35][6] ),
    .CLK(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24578_ (.D(_05455_),
    .Q(\design_top.MEM[35][7] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24579_ (.D(_05456_),
    .Q(\design_top.MEM[53][0] ),
    .CLK(clknet_leaf_404_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24580_ (.D(_05457_),
    .Q(\design_top.MEM[53][1] ),
    .CLK(clknet_leaf_430_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24581_ (.D(_05458_),
    .Q(\design_top.MEM[53][2] ),
    .CLK(clknet_leaf_404_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24582_ (.D(_05459_),
    .Q(\design_top.MEM[53][3] ),
    .CLK(clknet_leaf_430_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24583_ (.D(_05460_),
    .Q(\design_top.MEM[53][4] ),
    .CLK(clknet_leaf_428_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24584_ (.D(_05461_),
    .Q(\design_top.MEM[53][5] ),
    .CLK(clknet_leaf_423_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24585_ (.D(_05462_),
    .Q(\design_top.MEM[53][6] ),
    .CLK(clknet_leaf_422_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24586_ (.D(_05463_),
    .Q(\design_top.MEM[53][7] ),
    .CLK(clknet_leaf_423_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24587_ (.D(_05464_),
    .Q(\design_top.MEM[34][0] ),
    .CLK(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24588_ (.D(_05465_),
    .Q(\design_top.MEM[34][1] ),
    .CLK(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24589_ (.D(_05466_),
    .Q(\design_top.MEM[34][2] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24590_ (.D(_05467_),
    .Q(\design_top.MEM[34][3] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24591_ (.D(_05468_),
    .Q(\design_top.MEM[34][4] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24592_ (.D(_05469_),
    .Q(\design_top.MEM[34][5] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24593_ (.D(_05470_),
    .Q(\design_top.MEM[34][6] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24594_ (.D(_05471_),
    .Q(\design_top.MEM[34][7] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24595_ (.D(_05472_),
    .Q(\design_top.MEM[19][0] ),
    .CLK(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24596_ (.D(_05473_),
    .Q(\design_top.MEM[19][1] ),
    .CLK(clknet_leaf_437_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24597_ (.D(_05474_),
    .Q(\design_top.MEM[19][2] ),
    .CLK(clknet_leaf_437_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24598_ (.D(_05475_),
    .Q(\design_top.MEM[19][3] ),
    .CLK(clknet_leaf_445_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24599_ (.D(_05476_),
    .Q(\design_top.MEM[19][4] ),
    .CLK(clknet_leaf_444_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24600_ (.D(_05477_),
    .Q(\design_top.MEM[19][5] ),
    .CLK(clknet_leaf_444_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24601_ (.D(_05478_),
    .Q(\design_top.MEM[19][6] ),
    .CLK(clknet_leaf_444_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24602_ (.D(_05479_),
    .Q(\design_top.MEM[19][7] ),
    .CLK(clknet_leaf_444_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24603_ (.D(_05480_),
    .Q(\design_top.MEM[18][0] ),
    .CLK(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24604_ (.D(_05481_),
    .Q(\design_top.MEM[18][1] ),
    .CLK(clknet_leaf_445_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24605_ (.D(_05482_),
    .Q(\design_top.MEM[18][2] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24606_ (.D(_05483_),
    .Q(\design_top.MEM[18][3] ),
    .CLK(clknet_leaf_445_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24607_ (.D(_05484_),
    .Q(\design_top.MEM[18][4] ),
    .CLK(clknet_leaf_445_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24608_ (.D(_05485_),
    .Q(\design_top.MEM[18][5] ),
    .CLK(clknet_leaf_443_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24609_ (.D(_05486_),
    .Q(\design_top.MEM[18][6] ),
    .CLK(clknet_leaf_446_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24610_ (.D(_05487_),
    .Q(\design_top.MEM[18][7] ),
    .CLK(clknet_5_0_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24611_ (.D(_05488_),
    .Q(\design_top.MEM[33][0] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24612_ (.D(_05489_),
    .Q(\design_top.MEM[33][1] ),
    .CLK(clknet_leaf_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24613_ (.D(_05490_),
    .Q(\design_top.MEM[33][2] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24614_ (.D(_05491_),
    .Q(\design_top.MEM[33][3] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24615_ (.D(_05492_),
    .Q(\design_top.MEM[33][4] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24616_ (.D(_05493_),
    .Q(\design_top.MEM[33][5] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24617_ (.D(_05494_),
    .Q(\design_top.MEM[33][6] ),
    .CLK(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24618_ (.D(_05495_),
    .Q(\design_top.MEM[33][7] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24619_ (.D(_05496_),
    .Q(\design_top.MEM[32][0] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24620_ (.D(_05497_),
    .Q(\design_top.MEM[32][1] ),
    .CLK(clknet_leaf_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24621_ (.D(_05498_),
    .Q(\design_top.MEM[32][2] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24622_ (.D(_05499_),
    .Q(\design_top.MEM[32][3] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24623_ (.D(_05500_),
    .Q(\design_top.MEM[32][4] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24624_ (.D(_05501_),
    .Q(\design_top.MEM[32][5] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24625_ (.D(_05502_),
    .Q(\design_top.MEM[32][6] ),
    .CLK(clknet_leaf_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24626_ (.D(_05503_),
    .Q(\design_top.MEM[32][7] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24627_ (.D(_05504_),
    .Q(\design_top.MEM[17][0] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24628_ (.D(_05505_),
    .Q(\design_top.MEM[17][1] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24629_ (.D(_05506_),
    .Q(\design_top.MEM[17][2] ),
    .CLK(clknet_leaf_437_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24630_ (.D(_05507_),
    .Q(\design_top.MEM[17][3] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24631_ (.D(_05508_),
    .Q(\design_top.MEM[17][4] ),
    .CLK(clknet_leaf_446_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24632_ (.D(_05509_),
    .Q(\design_top.MEM[17][5] ),
    .CLK(clknet_leaf_446_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24633_ (.D(_05510_),
    .Q(\design_top.MEM[17][6] ),
    .CLK(clknet_leaf_446_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24634_ (.D(_05511_),
    .Q(\design_top.MEM[17][7] ),
    .CLK(clknet_leaf_446_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24635_ (.D(_05512_),
    .Q(\design_top.MEM[16][0] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24636_ (.D(_05513_),
    .Q(\design_top.MEM[16][1] ),
    .CLK(clknet_leaf_437_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24637_ (.D(_05514_),
    .Q(\design_top.MEM[16][2] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24638_ (.D(_05515_),
    .Q(\design_top.MEM[16][3] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24639_ (.D(_05516_),
    .Q(\design_top.MEM[16][4] ),
    .CLK(clknet_leaf_445_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24640_ (.D(_05517_),
    .Q(\design_top.MEM[16][5] ),
    .CLK(clknet_leaf_443_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24641_ (.D(_05518_),
    .Q(\design_top.MEM[16][6] ),
    .CLK(clknet_leaf_446_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24642_ (.D(_05519_),
    .Q(\design_top.MEM[16][7] ),
    .CLK(clknet_leaf_446_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24643_ (.D(_05520_),
    .Q(\design_top.MEM[15][0] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24644_ (.D(_05521_),
    .Q(\design_top.MEM[15][1] ),
    .CLK(clknet_leaf_39_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24645_ (.D(_05522_),
    .Q(\design_top.MEM[15][2] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24646_ (.D(_05523_),
    .Q(\design_top.MEM[15][3] ),
    .CLK(clknet_leaf_37_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24647_ (.D(_05524_),
    .Q(\design_top.MEM[15][4] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24648_ (.D(_05525_),
    .Q(\design_top.MEM[15][5] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24649_ (.D(_05526_),
    .Q(\design_top.MEM[15][6] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24650_ (.D(_05527_),
    .Q(\design_top.MEM[15][7] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24651_ (.D(_05528_),
    .Q(\design_top.MEM[14][0] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24652_ (.D(_05529_),
    .Q(\design_top.MEM[14][1] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24653_ (.D(_05530_),
    .Q(\design_top.MEM[14][2] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24654_ (.D(_05531_),
    .Q(\design_top.MEM[14][3] ),
    .CLK(clknet_leaf_37_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24655_ (.D(_05532_),
    .Q(\design_top.MEM[14][4] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24656_ (.D(_05533_),
    .Q(\design_top.MEM[14][5] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24657_ (.D(_05534_),
    .Q(\design_top.MEM[14][6] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24658_ (.D(_05535_),
    .Q(\design_top.MEM[14][7] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24659_ (.D(_05536_),
    .Q(\design_top.MEM[13][0] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24660_ (.D(_05537_),
    .Q(\design_top.MEM[13][1] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24661_ (.D(_05538_),
    .Q(\design_top.MEM[13][2] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24662_ (.D(_05539_),
    .Q(\design_top.MEM[13][3] ),
    .CLK(clknet_leaf_37_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24663_ (.D(_05540_),
    .Q(\design_top.MEM[13][4] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24664_ (.D(_05541_),
    .Q(\design_top.MEM[13][5] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24665_ (.D(_05542_),
    .Q(\design_top.MEM[13][6] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24666_ (.D(_05543_),
    .Q(\design_top.MEM[13][7] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24667_ (.D(_05544_),
    .Q(\design_top.MEM[12][0] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24668_ (.D(_05545_),
    .Q(\design_top.MEM[12][1] ),
    .CLK(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24669_ (.D(_05546_),
    .Q(\design_top.MEM[12][2] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24670_ (.D(_05547_),
    .Q(\design_top.MEM[12][3] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24671_ (.D(_05548_),
    .Q(\design_top.MEM[12][4] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24672_ (.D(_05549_),
    .Q(\design_top.MEM[12][5] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24673_ (.D(_05550_),
    .Q(\design_top.MEM[12][6] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24674_ (.D(_05551_),
    .Q(\design_top.MEM[12][7] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24675_ (.D(_05552_),
    .Q(\design_top.MEM[11][0] ),
    .CLK(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24676_ (.D(_05553_),
    .Q(\design_top.MEM[11][1] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24677_ (.D(_05554_),
    .Q(\design_top.MEM[11][2] ),
    .CLK(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24678_ (.D(_05555_),
    .Q(\design_top.MEM[11][3] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24679_ (.D(_05556_),
    .Q(\design_top.MEM[11][4] ),
    .CLK(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24680_ (.D(_05557_),
    .Q(\design_top.MEM[11][5] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24681_ (.D(_05558_),
    .Q(\design_top.MEM[11][6] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24682_ (.D(_05559_),
    .Q(\design_top.MEM[11][7] ),
    .CLK(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24683_ (.D(_05560_),
    .Q(\design_top.MEM[10][0] ),
    .CLK(clknet_leaf_29_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24684_ (.D(_05561_),
    .Q(\design_top.MEM[10][1] ),
    .CLK(clknet_leaf_29_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24685_ (.D(_05562_),
    .Q(\design_top.MEM[10][2] ),
    .CLK(clknet_leaf_29_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24686_ (.D(_05563_),
    .Q(\design_top.MEM[10][3] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24687_ (.D(_05564_),
    .Q(\design_top.MEM[10][4] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24688_ (.D(_05565_),
    .Q(\design_top.MEM[10][5] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24689_ (.D(_05566_),
    .Q(\design_top.MEM[10][6] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24690_ (.D(_05567_),
    .Q(\design_top.MEM[10][7] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24691_ (.D(_05568_),
    .Q(\design_top.MEM[0][0] ),
    .CLK(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24692_ (.D(_05569_),
    .Q(\design_top.MEM[0][1] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24693_ (.D(_05570_),
    .Q(\design_top.MEM[0][2] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24694_ (.D(_05571_),
    .Q(\design_top.MEM[0][3] ),
    .CLK(clknet_leaf_39_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24695_ (.D(_05572_),
    .Q(\design_top.MEM[0][4] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24696_ (.D(_05573_),
    .Q(\design_top.MEM[0][5] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24697_ (.D(_05574_),
    .Q(\design_top.MEM[0][6] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24698_ (.D(_05575_),
    .Q(\design_top.MEM[0][7] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24699_ (.D(_05576_),
    .Q(\design_top.core0.REG1[9][0] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24700_ (.D(_05577_),
    .Q(\design_top.core0.REG1[9][1] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24701_ (.D(_05578_),
    .Q(\design_top.core0.REG1[9][2] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24702_ (.D(_05579_),
    .Q(\design_top.core0.REG1[9][3] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24703_ (.D(_05580_),
    .Q(\design_top.core0.REG1[9][4] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24704_ (.D(_05581_),
    .Q(\design_top.core0.REG1[9][5] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24705_ (.D(_05582_),
    .Q(\design_top.core0.REG1[9][6] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24706_ (.D(_05583_),
    .Q(\design_top.core0.REG1[9][7] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24707_ (.D(_05584_),
    .Q(\design_top.core0.REG1[9][8] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24708_ (.D(_05585_),
    .Q(\design_top.core0.REG1[9][9] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24709_ (.D(_05586_),
    .Q(\design_top.core0.REG1[9][10] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24710_ (.D(_05587_),
    .Q(\design_top.core0.REG1[9][11] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24711_ (.D(_05588_),
    .Q(\design_top.core0.REG1[9][12] ),
    .CLK(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24712_ (.D(_05589_),
    .Q(\design_top.core0.REG1[9][13] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24713_ (.D(_05590_),
    .Q(\design_top.core0.REG1[9][14] ),
    .CLK(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24714_ (.D(_05591_),
    .Q(\design_top.core0.REG1[9][15] ),
    .CLK(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24715_ (.D(_05592_),
    .Q(\design_top.core0.REG1[9][16] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24716_ (.D(_05593_),
    .Q(\design_top.core0.REG1[9][17] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24717_ (.D(_05594_),
    .Q(\design_top.core0.REG1[9][18] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24718_ (.D(_05595_),
    .Q(\design_top.core0.REG1[9][19] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24719_ (.D(_05596_),
    .Q(\design_top.core0.REG1[9][20] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24720_ (.D(_05597_),
    .Q(\design_top.core0.REG1[9][21] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24721_ (.D(_05598_),
    .Q(\design_top.core0.REG1[9][22] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24722_ (.D(_05599_),
    .Q(\design_top.core0.REG1[9][23] ),
    .CLK(clknet_leaf_262_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24723_ (.D(_05600_),
    .Q(\design_top.core0.REG1[9][24] ),
    .CLK(clknet_leaf_253_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24724_ (.D(_05601_),
    .Q(\design_top.core0.REG1[9][25] ),
    .CLK(clknet_leaf_253_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24725_ (.D(_05602_),
    .Q(\design_top.core0.REG1[9][26] ),
    .CLK(clknet_leaf_253_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24726_ (.D(_05603_),
    .Q(\design_top.core0.REG1[9][27] ),
    .CLK(clknet_leaf_253_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24727_ (.D(_05604_),
    .Q(\design_top.core0.REG1[9][28] ),
    .CLK(clknet_leaf_255_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24728_ (.D(_05605_),
    .Q(\design_top.core0.REG1[9][29] ),
    .CLK(clknet_leaf_254_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24729_ (.D(_05606_),
    .Q(\design_top.core0.REG1[9][30] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24730_ (.D(_05607_),
    .Q(\design_top.core0.REG1[9][31] ),
    .CLK(clknet_leaf_251_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24731_ (.D(_05608_),
    .Q(\design_top.MEM[31][0] ),
    .CLK(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24732_ (.D(_05609_),
    .Q(\design_top.MEM[31][1] ),
    .CLK(clknet_leaf_437_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24733_ (.D(_05610_),
    .Q(\design_top.MEM[31][2] ),
    .CLK(clknet_leaf_436_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24734_ (.D(_05611_),
    .Q(\design_top.MEM[31][3] ),
    .CLK(clknet_leaf_437_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24735_ (.D(_05612_),
    .Q(\design_top.MEM[31][4] ),
    .CLK(clknet_leaf_444_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24736_ (.D(_05613_),
    .Q(\design_top.MEM[31][5] ),
    .CLK(clknet_leaf_444_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24737_ (.D(_05614_),
    .Q(\design_top.MEM[31][6] ),
    .CLK(clknet_leaf_444_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24738_ (.D(_05615_),
    .Q(\design_top.MEM[31][7] ),
    .CLK(clknet_leaf_444_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24739_ (.D(_05616_),
    .Q(\design_top.MEM[30][0] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24740_ (.D(_05617_),
    .Q(\design_top.MEM[30][1] ),
    .CLK(clknet_leaf_437_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24741_ (.D(_05618_),
    .Q(\design_top.MEM[30][2] ),
    .CLK(clknet_leaf_436_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24742_ (.D(_05619_),
    .Q(\design_top.MEM[30][3] ),
    .CLK(clknet_leaf_437_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24743_ (.D(_05620_),
    .Q(\design_top.MEM[30][4] ),
    .CLK(clknet_leaf_444_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24744_ (.D(_05621_),
    .Q(\design_top.MEM[30][5] ),
    .CLK(clknet_leaf_443_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24745_ (.D(_05622_),
    .Q(\design_top.MEM[30][6] ),
    .CLK(clknet_leaf_444_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24746_ (.D(_05623_),
    .Q(\design_top.MEM[30][7] ),
    .CLK(clknet_leaf_442_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24747_ (.D(_05624_),
    .Q(\design_top.MEM[2][0] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24748_ (.D(_05625_),
    .Q(\design_top.MEM[2][1] ),
    .CLK(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24749_ (.D(_05626_),
    .Q(\design_top.MEM[2][2] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24750_ (.D(_05627_),
    .Q(\design_top.MEM[2][3] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24751_ (.D(_05628_),
    .Q(\design_top.MEM[2][4] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24752_ (.D(_05629_),
    .Q(\design_top.MEM[2][5] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24753_ (.D(_05630_),
    .Q(\design_top.MEM[2][6] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24754_ (.D(_05631_),
    .Q(\design_top.MEM[2][7] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24755_ (.D(_05632_),
    .Q(\design_top.MEM[29][0] ),
    .CLK(clknet_leaf_436_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24756_ (.D(_05633_),
    .Q(\design_top.MEM[29][1] ),
    .CLK(clknet_leaf_436_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24757_ (.D(_05634_),
    .Q(\design_top.MEM[29][2] ),
    .CLK(clknet_leaf_435_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24758_ (.D(_05635_),
    .Q(\design_top.MEM[29][3] ),
    .CLK(clknet_leaf_438_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24759_ (.D(_05636_),
    .Q(\design_top.MEM[29][4] ),
    .CLK(clknet_leaf_438_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24760_ (.D(_05637_),
    .Q(\design_top.MEM[29][5] ),
    .CLK(clknet_leaf_442_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24761_ (.D(_05638_),
    .Q(\design_top.MEM[29][6] ),
    .CLK(clknet_leaf_442_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24762_ (.D(_05639_),
    .Q(\design_top.MEM[29][7] ),
    .CLK(clknet_leaf_441_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24763_ (.D(_05640_),
    .Q(\design_top.MEM[28][0] ),
    .CLK(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24764_ (.D(_05641_),
    .Q(\design_top.MEM[28][1] ),
    .CLK(clknet_leaf_437_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24765_ (.D(_05642_),
    .Q(\design_top.MEM[28][2] ),
    .CLK(clknet_leaf_436_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24766_ (.D(_05643_),
    .Q(\design_top.MEM[28][3] ),
    .CLK(clknet_leaf_444_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24767_ (.D(_05644_),
    .Q(\design_top.MEM[28][4] ),
    .CLK(clknet_leaf_444_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24768_ (.D(_05645_),
    .Q(\design_top.MEM[28][5] ),
    .CLK(clknet_leaf_442_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24769_ (.D(_05646_),
    .Q(\design_top.MEM[28][6] ),
    .CLK(clknet_leaf_444_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24770_ (.D(_05647_),
    .Q(\design_top.MEM[28][7] ),
    .CLK(clknet_leaf_443_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24771_ (.D(_05648_),
    .Q(\design_top.MEM[27][0] ),
    .CLK(clknet_leaf_434_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24772_ (.D(_05649_),
    .Q(\design_top.MEM[27][1] ),
    .CLK(clknet_leaf_435_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24773_ (.D(_05650_),
    .Q(\design_top.MEM[27][2] ),
    .CLK(clknet_leaf_435_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24774_ (.D(_05651_),
    .Q(\design_top.MEM[27][3] ),
    .CLK(clknet_leaf_439_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24775_ (.D(_05652_),
    .Q(\design_top.MEM[27][4] ),
    .CLK(clknet_leaf_438_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24776_ (.D(_05653_),
    .Q(\design_top.MEM[27][5] ),
    .CLK(clknet_leaf_440_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24777_ (.D(_05654_),
    .Q(\design_top.MEM[27][6] ),
    .CLK(clknet_leaf_440_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24778_ (.D(_05655_),
    .Q(\design_top.MEM[27][7] ),
    .CLK(clknet_leaf_440_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24779_ (.D(_05656_),
    .Q(io_out[14]),
    .CLK(clknet_leaf_343_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24780_ (.D(_05657_),
    .Q(\design_top.TIMER[0] ),
    .CLK(clknet_leaf_342_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24781_ (.D(_05658_),
    .Q(\design_top.TIMER[1] ),
    .CLK(clknet_leaf_343_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24782_ (.D(_05659_),
    .Q(\design_top.TIMER[2] ),
    .CLK(clknet_leaf_342_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24783_ (.D(_05660_),
    .Q(\design_top.TIMER[3] ),
    .CLK(clknet_leaf_342_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24784_ (.D(_05661_),
    .Q(\design_top.TIMER[4] ),
    .CLK(clknet_leaf_342_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24785_ (.D(_05662_),
    .Q(\design_top.TIMER[5] ),
    .CLK(clknet_leaf_342_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24786_ (.D(_05663_),
    .Q(\design_top.TIMER[6] ),
    .CLK(clknet_leaf_339_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24787_ (.D(_05664_),
    .Q(\design_top.TIMER[7] ),
    .CLK(clknet_leaf_339_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24788_ (.D(_05665_),
    .Q(\design_top.TIMER[8] ),
    .CLK(clknet_leaf_339_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24789_ (.D(_05666_),
    .Q(\design_top.TIMER[9] ),
    .CLK(clknet_leaf_349_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24790_ (.D(_05667_),
    .Q(\design_top.TIMER[10] ),
    .CLK(clknet_leaf_349_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24791_ (.D(_05668_),
    .Q(\design_top.TIMER[11] ),
    .CLK(clknet_leaf_349_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24792_ (.D(_05669_),
    .Q(\design_top.TIMER[12] ),
    .CLK(clknet_leaf_349_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24793_ (.D(_05670_),
    .Q(\design_top.TIMER[13] ),
    .CLK(clknet_leaf_342_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24794_ (.D(_05671_),
    .Q(\design_top.TIMER[14] ),
    .CLK(clknet_leaf_342_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24795_ (.D(_05672_),
    .Q(\design_top.TIMER[15] ),
    .CLK(clknet_leaf_345_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24796_ (.D(_05673_),
    .Q(\design_top.TIMER[16] ),
    .CLK(clknet_leaf_344_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24797_ (.D(_05674_),
    .Q(\design_top.TIMER[17] ),
    .CLK(clknet_leaf_344_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24798_ (.D(_05675_),
    .Q(\design_top.TIMER[18] ),
    .CLK(clknet_leaf_343_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24799_ (.D(_05676_),
    .Q(\design_top.TIMER[19] ),
    .CLK(clknet_leaf_344_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24800_ (.D(_05677_),
    .Q(\design_top.TIMER[20] ),
    .CLK(clknet_leaf_372_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24801_ (.D(_05678_),
    .Q(\design_top.TIMER[21] ),
    .CLK(clknet_5_14_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24802_ (.D(_05679_),
    .Q(\design_top.TIMER[22] ),
    .CLK(clknet_leaf_332_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24803_ (.D(_05680_),
    .Q(\design_top.TIMER[23] ),
    .CLK(clknet_leaf_344_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24804_ (.D(_05681_),
    .Q(\design_top.TIMER[24] ),
    .CLK(clknet_leaf_332_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24805_ (.D(_05682_),
    .Q(\design_top.TIMER[25] ),
    .CLK(clknet_leaf_332_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24806_ (.D(_05683_),
    .Q(\design_top.TIMER[26] ),
    .CLK(clknet_leaf_332_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24807_ (.D(_05684_),
    .Q(\design_top.TIMER[27] ),
    .CLK(clknet_leaf_333_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24808_ (.D(_05685_),
    .Q(\design_top.TIMER[28] ),
    .CLK(clknet_leaf_343_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24809_ (.D(_05686_),
    .Q(\design_top.TIMER[29] ),
    .CLK(clknet_leaf_343_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24810_ (.D(_05687_),
    .Q(\design_top.TIMER[30] ),
    .CLK(clknet_leaf_343_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24811_ (.D(_05688_),
    .Q(\design_top.TIMER[31] ),
    .CLK(clknet_leaf_343_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24812_ (.D(_05689_),
    .Q(\design_top.uart0.UART_XBAUD[0] ),
    .CLK(clknet_leaf_343_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24813_ (.D(_05690_),
    .Q(\design_top.uart0.UART_XBAUD[1] ),
    .CLK(clknet_leaf_343_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24814_ (.D(_05691_),
    .Q(\design_top.uart0.UART_XBAUD[2] ),
    .CLK(clknet_leaf_341_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24815_ (.D(_05692_),
    .Q(\design_top.uart0.UART_XBAUD[3] ),
    .CLK(clknet_leaf_341_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24816_ (.D(_05693_),
    .Q(\design_top.uart0.UART_XBAUD[4] ),
    .CLK(clknet_leaf_341_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24817_ (.D(_05694_),
    .Q(\design_top.uart0.UART_XBAUD[5] ),
    .CLK(clknet_leaf_334_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24818_ (.D(_05695_),
    .Q(\design_top.uart0.UART_XBAUD[6] ),
    .CLK(clknet_leaf_334_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24819_ (.D(_05696_),
    .Q(\design_top.uart0.UART_XBAUD[7] ),
    .CLK(clknet_leaf_334_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24820_ (.D(_05697_),
    .Q(\design_top.uart0.UART_XBAUD[8] ),
    .CLK(clknet_leaf_334_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24821_ (.D(_05698_),
    .Q(\design_top.uart0.UART_XBAUD[9] ),
    .CLK(clknet_leaf_334_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24822_ (.D(_05699_),
    .Q(\design_top.uart0.UART_XBAUD[10] ),
    .CLK(clknet_leaf_334_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24823_ (.D(_05700_),
    .Q(\design_top.uart0.UART_XBAUD[11] ),
    .CLK(clknet_leaf_333_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24824_ (.D(_05701_),
    .Q(\design_top.uart0.UART_XBAUD[12] ),
    .CLK(clknet_leaf_333_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24825_ (.D(_05702_),
    .Q(\design_top.uart0.UART_XBAUD[13] ),
    .CLK(clknet_leaf_343_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24826_ (.D(_05703_),
    .Q(\design_top.uart0.UART_XBAUD[14] ),
    .CLK(clknet_leaf_341_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24827_ (.D(_05704_),
    .Q(\design_top.uart0.UART_XBAUD[15] ),
    .CLK(clknet_leaf_341_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24828_ (.D(_05705_),
    .Q(\design_top.uart0.UART_RBAUD[0] ),
    .CLK(clknet_leaf_335_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24829_ (.D(_05706_),
    .Q(\design_top.uart0.UART_RBAUD[3] ),
    .CLK(clknet_leaf_338_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24830_ (.D(_05707_),
    .Q(\design_top.uart0.UART_RBAUD[5] ),
    .CLK(clknet_leaf_338_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24831_ (.D(_05708_),
    .Q(\design_top.uart0.UART_RBAUD[8] ),
    .CLK(clknet_leaf_340_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24832_ (.D(_05709_),
    .Q(\design_top.uart0.UART_RBAUD[10] ),
    .CLK(clknet_leaf_335_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24833_ (.D(_05710_),
    .Q(\design_top.uart0.UART_RBAUD[11] ),
    .CLK(clknet_leaf_335_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24834_ (.D(_05711_),
    .Q(\design_top.uart0.UART_RBAUD[12] ),
    .CLK(clknet_leaf_335_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24835_ (.D(_05712_),
    .Q(\design_top.uart0.UART_RBAUD[13] ),
    .CLK(clknet_leaf_335_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24836_ (.D(_05713_),
    .Q(\design_top.uart0.UART_RBAUD[14] ),
    .CLK(clknet_opt_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24837_ (.D(_05714_),
    .Q(\design_top.uart0.UART_RBAUD[15] ),
    .CLK(clknet_leaf_338_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24838_ (.D(_05715_),
    .Q(\design_top.IRES[0] ),
    .CLK(clknet_leaf_353_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24839_ (.D(_05716_),
    .Q(\design_top.IRES[1] ),
    .CLK(clknet_leaf_352_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24840_ (.D(_05717_),
    .Q(\design_top.IRES[2] ),
    .CLK(clknet_leaf_352_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24841_ (.D(_05718_),
    .Q(\design_top.IRES[3] ),
    .CLK(clknet_leaf_352_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24842_ (.D(_05719_),
    .Q(\design_top.IRES[4] ),
    .CLK(clknet_leaf_352_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24843_ (.D(_05720_),
    .Q(\design_top.IRES[5] ),
    .CLK(clknet_leaf_352_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24844_ (.D(_05721_),
    .Q(\design_top.IRES[6] ),
    .CLK(clknet_leaf_352_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24845_ (.D(_05722_),
    .Q(\design_top.IRES[7] ),
    .CLK(clknet_leaf_352_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24846_ (.D(_05723_),
    .Q(\design_top.core0.RESMODE[0] ),
    .CLK(clknet_leaf_292_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24847_ (.D(_05724_),
    .Q(\design_top.core0.RESMODE[1] ),
    .CLK(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24848_ (.D(_05725_),
    .Q(\design_top.core0.RESMODE[2] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24849_ (.D(_05726_),
    .Q(\design_top.core0.RESMODE[3] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24850_ (.D(_05727_),
    .Q(\design_top.uart0.UART_RBAUD[1] ),
    .CLK(clknet_leaf_338_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24851_ (.D(_05728_),
    .Q(\design_top.uart0.UART_RBAUD[2] ),
    .CLK(clknet_leaf_338_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24852_ (.D(_05729_),
    .Q(\design_top.uart0.UART_RBAUD[4] ),
    .CLK(clknet_leaf_338_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24853_ (.D(_05730_),
    .Q(\design_top.uart0.UART_RBAUD[6] ),
    .CLK(clknet_leaf_340_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24854_ (.D(_05731_),
    .Q(\design_top.uart0.UART_RBAUD[7] ),
    .CLK(clknet_leaf_335_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24855_ (.D(_05732_),
    .Q(\design_top.uart0.UART_RBAUD[9] ),
    .CLK(clknet_leaf_335_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24856_ (.D(_05733_),
    .Q(\design_top.uart0.UART_RSTATE[0] ),
    .CLK(clknet_leaf_349_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24857_ (.D(_05734_),
    .Q(\design_top.uart0.UART_RSTATE[1] ),
    .CLK(clknet_leaf_350_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24858_ (.D(_05735_),
    .Q(\design_top.uart0.UART_RSTATE[2] ),
    .CLK(clknet_leaf_350_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24859_ (.D(_05736_),
    .Q(\design_top.uart0.UART_RSTATE[3] ),
    .CLK(clknet_leaf_350_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24860_ (.D(_05737_),
    .Q(\design_top.uart0.UART_XSTATE[0] ),
    .CLK(clknet_leaf_346_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24861_ (.D(_05738_),
    .Q(\design_top.uart0.UART_XSTATE[1] ),
    .CLK(clknet_leaf_346_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24862_ (.D(_05739_),
    .Q(\design_top.uart0.UART_XSTATE[2] ),
    .CLK(clknet_leaf_346_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24863_ (.D(_05740_),
    .Q(\design_top.uart0.UART_XSTATE[3] ),
    .CLK(clknet_leaf_345_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24864_ (.D(_05741_),
    .Q(\design_top.DACK[0] ),
    .CLK(clknet_leaf_368_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24865_ (.D(_05742_),
    .Q(\design_top.DACK[1] ),
    .CLK(clknet_leaf_369_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24866_ (.D(_05743_),
    .Q(_00689_),
    .CLK(clknet_leaf_309_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24867_ (.D(_05744_),
    .Q(_00690_),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24868_ (.D(_05745_),
    .Q(_00691_),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24869_ (.D(_05746_),
    .Q(_00692_),
    .CLK(clknet_leaf_311_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24870_ (.D(_05747_),
    .Q(_00685_),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24871_ (.D(_05748_),
    .Q(_00686_),
    .CLK(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24872_ (.D(_05749_),
    .Q(_00687_),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24873_ (.D(_05750_),
    .Q(_00688_),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24874_ (.D(_05751_),
    .Q(\design_top.MEM[9][24] ),
    .CLK(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24875_ (.D(_05752_),
    .Q(\design_top.MEM[9][25] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24876_ (.D(_05753_),
    .Q(\design_top.MEM[9][26] ),
    .CLK(clknet_leaf_388_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24877_ (.D(_05754_),
    .Q(\design_top.MEM[9][27] ),
    .CLK(clknet_leaf_395_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24878_ (.D(_05755_),
    .Q(\design_top.MEM[9][28] ),
    .CLK(clknet_leaf_395_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24879_ (.D(_05756_),
    .Q(\design_top.MEM[9][29] ),
    .CLK(clknet_leaf_395_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24880_ (.D(_05757_),
    .Q(\design_top.MEM[9][30] ),
    .CLK(clknet_leaf_394_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24881_ (.D(_05758_),
    .Q(\design_top.MEM[9][31] ),
    .CLK(clknet_leaf_393_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24882_ (.D(_05759_),
    .Q(io_out[16]),
    .CLK(clknet_leaf_319_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24883_ (.D(_05760_),
    .Q(io_out[17]),
    .CLK(clknet_leaf_319_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24884_ (.D(_05761_),
    .Q(\design_top.core0.FLUSH[0] ),
    .CLK(clknet_leaf_307_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24885_ (.D(_05762_),
    .Q(\design_top.core0.FLUSH[1] ),
    .CLK(clknet_leaf_307_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24886_ (.D(_05763_),
    .Q(io_out[18]),
    .CLK(clknet_leaf_311_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24887_ (.D(_05764_),
    .Q(io_out[19]),
    .CLK(clknet_leaf_312_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24888_ (.D(_05765_),
    .Q(\design_top.IADDR[4] ),
    .CLK(clknet_leaf_312_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24889_ (.D(_05766_),
    .Q(\design_top.IADDR[5] ),
    .CLK(clknet_leaf_312_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24890_ (.D(_05767_),
    .Q(\design_top.IADDR[6] ),
    .CLK(clknet_leaf_311_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24891_ (.D(_05768_),
    .Q(\design_top.IADDR[7] ),
    .CLK(clknet_leaf_310_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24892_ (.D(_05769_),
    .Q(\design_top.IADDR[8] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24893_ (.D(_05770_),
    .Q(\design_top.IADDR[9] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24894_ (.D(_05771_),
    .Q(\design_top.IADDR[10] ),
    .CLK(clknet_leaf_305_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24895_ (.D(_05772_),
    .Q(\design_top.IADDR[11] ),
    .CLK(clknet_leaf_305_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24896_ (.D(_05773_),
    .Q(\design_top.IADDR[12] ),
    .CLK(clknet_leaf_291_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24897_ (.D(_05774_),
    .Q(\design_top.IADDR[13] ),
    .CLK(clknet_leaf_291_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24898_ (.D(_05775_),
    .Q(\design_top.IADDR[14] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24899_ (.D(_05776_),
    .Q(\design_top.IADDR[15] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24900_ (.D(_05777_),
    .Q(\design_top.IADDR[16] ),
    .CLK(clknet_leaf_288_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24901_ (.D(_05778_),
    .Q(\design_top.IADDR[17] ),
    .CLK(clknet_leaf_288_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24902_ (.D(_05779_),
    .Q(\design_top.IADDR[18] ),
    .CLK(clknet_leaf_288_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24903_ (.D(_05780_),
    .Q(\design_top.IADDR[19] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24904_ (.D(_05781_),
    .Q(\design_top.IADDR[20] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24905_ (.D(_05782_),
    .Q(\design_top.IADDR[21] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24906_ (.D(_05783_),
    .Q(\design_top.IADDR[22] ),
    .CLK(clknet_leaf_284_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24907_ (.D(_05784_),
    .Q(\design_top.IADDR[23] ),
    .CLK(clknet_leaf_282_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24908_ (.D(_05785_),
    .Q(\design_top.IADDR[24] ),
    .CLK(clknet_leaf_282_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24909_ (.D(_05786_),
    .Q(\design_top.IADDR[25] ),
    .CLK(clknet_leaf_282_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24910_ (.D(_05787_),
    .Q(\design_top.IADDR[26] ),
    .CLK(clknet_leaf_283_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24911_ (.D(_05788_),
    .Q(\design_top.IADDR[27] ),
    .CLK(clknet_leaf_283_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24912_ (.D(_05789_),
    .Q(\design_top.IADDR[28] ),
    .CLK(clknet_leaf_330_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24913_ (.D(_05790_),
    .Q(\design_top.IADDR[29] ),
    .CLK(clknet_leaf_283_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24914_ (.D(_05791_),
    .Q(\design_top.IADDR[30] ),
    .CLK(clknet_leaf_283_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24915_ (.D(_05792_),
    .Q(\design_top.IADDR[31] ),
    .CLK(clknet_leaf_329_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24916_ (.D(_05793_),
    .Q(\design_top.core0.XIDATA[7] ),
    .CLK(clknet_leaf_291_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24917_ (.D(_05794_),
    .Q(\design_top.core0.XIDATA[8] ),
    .CLK(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24918_ (.D(_05795_),
    .Q(\design_top.core0.XIDATA[9] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24919_ (.D(_05796_),
    .Q(\design_top.core0.XIDATA[10] ),
    .CLK(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24920_ (.D(_05797_),
    .Q(\design_top.core0.FCT3[0] ),
    .CLK(clknet_leaf_291_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24921_ (.D(_05798_),
    .Q(\design_top.core0.FCT3[1] ),
    .CLK(clknet_leaf_291_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24922_ (.D(_05799_),
    .Q(\design_top.core0.FCT3[2] ),
    .CLK(clknet_leaf_291_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24923_ (.D(_05800_),
    .Q(\design_top.core0.S1PTR[0] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24924_ (.D(_05801_),
    .Q(\design_top.core0.S1PTR[1] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24925_ (.D(_05802_),
    .Q(\design_top.core0.S1PTR[2] ),
    .CLK(clknet_leaf_309_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24926_ (.D(_05803_),
    .Q(\design_top.core0.S1PTR[3] ),
    .CLK(clknet_leaf_309_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24927_ (.D(_05804_),
    .Q(\design_top.core0.S2PTR[0] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24928_ (.D(_05805_),
    .Q(\design_top.core0.S2PTR[1] ),
    .CLK(clknet_leaf_311_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24929_ (.D(_05806_),
    .Q(\design_top.core0.S2PTR[2] ),
    .CLK(clknet_leaf_311_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24930_ (.D(_05807_),
    .Q(\design_top.core0.S2PTR[3] ),
    .CLK(clknet_leaf_312_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24931_ (.D(_05808_),
    .Q(\design_top.core0.FCT7[5] ),
    .CLK(clknet_leaf_320_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24932_ (.D(_05809_),
    .Q(\design_top.core0.XLUI ),
    .CLK(clknet_leaf_308_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24933_ (.D(_05810_),
    .Q(\design_top.core0.XAUIPC ),
    .CLK(clknet_leaf_308_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24934_ (.D(_05811_),
    .Q(\design_top.core0.XJAL ),
    .CLK(clknet_leaf_308_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24935_ (.D(_05812_),
    .Q(\design_top.core0.XJALR ),
    .CLK(clknet_leaf_308_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24936_ (.D(_05813_),
    .Q(\design_top.core0.XBCC ),
    .CLK(clknet_leaf_308_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24937_ (.D(_05814_),
    .Q(\design_top.core0.XLCC ),
    .CLK(clknet_leaf_309_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24938_ (.D(_05815_),
    .Q(\design_top.core0.XSCC ),
    .CLK(clknet_leaf_307_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24939_ (.D(_05816_),
    .Q(\design_top.core0.XMCC ),
    .CLK(clknet_leaf_312_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24940_ (.D(_05817_),
    .Q(\design_top.core0.XRCC ),
    .CLK(clknet_leaf_308_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24941_ (.D(_05818_),
    .Q(\design_top.core0.SIMM[12] ),
    .CLK(clknet_leaf_325_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24942_ (.D(_05819_),
    .Q(\design_top.core0.SIMM[13] ),
    .CLK(clknet_leaf_290_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24943_ (.D(_05820_),
    .Q(\design_top.core0.SIMM[14] ),
    .CLK(clknet_leaf_290_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24944_ (.D(_05821_),
    .Q(\design_top.core0.SIMM[15] ),
    .CLK(clknet_leaf_290_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24945_ (.D(_05822_),
    .Q(\design_top.core0.SIMM[16] ),
    .CLK(clknet_leaf_289_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24946_ (.D(_05823_),
    .Q(\design_top.core0.SIMM[17] ),
    .CLK(clknet_leaf_325_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24947_ (.D(_05824_),
    .Q(\design_top.core0.SIMM[18] ),
    .CLK(clknet_leaf_325_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24948_ (.D(_05825_),
    .Q(\design_top.core0.SIMM[19] ),
    .CLK(clknet_leaf_325_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24949_ (.D(_05826_),
    .Q(\design_top.core0.SIMM[20] ),
    .CLK(clknet_5_26_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24950_ (.D(_05827_),
    .Q(\design_top.core0.SIMM[21] ),
    .CLK(clknet_leaf_329_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24951_ (.D(_05828_),
    .Q(\design_top.core0.SIMM[22] ),
    .CLK(clknet_leaf_329_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24952_ (.D(_05829_),
    .Q(\design_top.core0.SIMM[23] ),
    .CLK(clknet_leaf_329_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24953_ (.D(_05830_),
    .Q(\design_top.core0.SIMM[24] ),
    .CLK(clknet_leaf_331_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24954_ (.D(_05831_),
    .Q(\design_top.core0.SIMM[25] ),
    .CLK(clknet_leaf_331_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24955_ (.D(_05832_),
    .Q(\design_top.core0.SIMM[26] ),
    .CLK(clknet_leaf_325_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24956_ (.D(_05833_),
    .Q(\design_top.core0.SIMM[27] ),
    .CLK(clknet_leaf_327_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24957_ (.D(_05834_),
    .Q(\design_top.core0.SIMM[28] ),
    .CLK(clknet_leaf_328_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24958_ (.D(_05835_),
    .Q(\design_top.core0.SIMM[29] ),
    .CLK(clknet_leaf_328_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24959_ (.D(_05836_),
    .Q(\design_top.core0.SIMM[30] ),
    .CLK(clknet_leaf_327_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24960_ (.D(_05837_),
    .Q(\design_top.core0.SIMM[31] ),
    .CLK(clknet_opt_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24961_ (.D(_05838_),
    .Q(\design_top.core0.SIMM[0] ),
    .CLK(clknet_leaf_321_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24962_ (.D(_05839_),
    .Q(\design_top.core0.SIMM[1] ),
    .CLK(clknet_leaf_322_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24963_ (.D(_05840_),
    .Q(\design_top.core0.SIMM[2] ),
    .CLK(clknet_leaf_318_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24964_ (.D(_05841_),
    .Q(\design_top.core0.SIMM[3] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24965_ (.D(_05842_),
    .Q(\design_top.core0.SIMM[4] ),
    .CLK(clknet_leaf_318_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24966_ (.D(_05843_),
    .Q(\design_top.core0.SIMM[5] ),
    .CLK(clknet_leaf_318_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24967_ (.D(_05844_),
    .Q(\design_top.core0.SIMM[6] ),
    .CLK(clknet_leaf_316_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24968_ (.D(_05845_),
    .Q(\design_top.core0.SIMM[7] ),
    .CLK(clknet_leaf_316_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24969_ (.D(_05846_),
    .Q(\design_top.core0.SIMM[8] ),
    .CLK(clknet_leaf_319_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24970_ (.D(_05847_),
    .Q(\design_top.core0.SIMM[9] ),
    .CLK(clknet_leaf_318_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24971_ (.D(_05848_),
    .Q(\design_top.core0.SIMM[10] ),
    .CLK(clknet_leaf_319_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24972_ (.D(_05849_),
    .Q(\design_top.core0.SIMM[11] ),
    .CLK(clknet_leaf_307_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24973_ (.D(_05850_),
    .Q(\design_top.core0.UIMM[12] ),
    .CLK(clknet_leaf_320_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24974_ (.D(_05851_),
    .Q(\design_top.core0.UIMM[13] ),
    .CLK(clknet_5_24_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24975_ (.D(_05852_),
    .Q(\design_top.core0.UIMM[14] ),
    .CLK(clknet_leaf_321_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24976_ (.D(_05853_),
    .Q(\design_top.core0.UIMM[15] ),
    .CLK(clknet_leaf_320_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24977_ (.D(_05854_),
    .Q(\design_top.core0.UIMM[16] ),
    .CLK(clknet_leaf_321_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24978_ (.D(_05855_),
    .Q(\design_top.core0.UIMM[17] ),
    .CLK(clknet_leaf_321_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24979_ (.D(_05856_),
    .Q(\design_top.core0.UIMM[18] ),
    .CLK(clknet_leaf_321_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24980_ (.D(_05857_),
    .Q(\design_top.core0.UIMM[19] ),
    .CLK(clknet_leaf_321_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24981_ (.D(_05858_),
    .Q(\design_top.core0.UIMM[20] ),
    .CLK(clknet_leaf_321_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24982_ (.D(_05859_),
    .Q(\design_top.core0.UIMM[21] ),
    .CLK(clknet_leaf_320_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24983_ (.D(_05860_),
    .Q(\design_top.core0.UIMM[22] ),
    .CLK(clknet_leaf_320_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24984_ (.D(_05861_),
    .Q(\design_top.core0.UIMM[23] ),
    .CLK(clknet_leaf_321_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24985_ (.D(_05862_),
    .Q(\design_top.core0.UIMM[24] ),
    .CLK(clknet_leaf_321_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24986_ (.D(_05863_),
    .Q(\design_top.core0.UIMM[25] ),
    .CLK(clknet_leaf_322_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24987_ (.D(_05864_),
    .Q(\design_top.core0.UIMM[26] ),
    .CLK(clknet_leaf_322_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24988_ (.D(_05865_),
    .Q(\design_top.core0.UIMM[27] ),
    .CLK(clknet_leaf_318_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24989_ (.D(_05866_),
    .Q(\design_top.core0.UIMM[28] ),
    .CLK(clknet_leaf_318_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24990_ (.D(_05867_),
    .Q(\design_top.core0.UIMM[29] ),
    .CLK(clknet_leaf_318_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24991_ (.D(_05868_),
    .Q(\design_top.core0.UIMM[30] ),
    .CLK(clknet_leaf_322_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24992_ (.D(_05869_),
    .Q(\design_top.core0.UIMM[31] ),
    .CLK(clknet_leaf_322_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24993_ (.D(_05870_),
    .Q(\design_top.IOMUX[3][0] ),
    .CLK(clknet_leaf_346_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24994_ (.D(_05871_),
    .Q(\design_top.IOMUX[3][1] ),
    .CLK(clknet_leaf_346_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24995_ (.D(_05872_),
    .Q(\design_top.IOMUX[3][2] ),
    .CLK(clknet_leaf_345_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24996_ (.D(_05873_),
    .Q(\design_top.IOMUX[3][3] ),
    .CLK(clknet_leaf_345_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24997_ (.D(_05874_),
    .Q(\design_top.IOMUX[3][4] ),
    .CLK(clknet_leaf_345_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24998_ (.D(_05875_),
    .Q(\design_top.IOMUX[3][5] ),
    .CLK(clknet_leaf_369_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _24999_ (.D(_05876_),
    .Q(\design_top.IOMUX[3][6] ),
    .CLK(clknet_leaf_369_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25000_ (.D(_05877_),
    .Q(\design_top.IOMUX[3][7] ),
    .CLK(clknet_leaf_348_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25001_ (.D(_05878_),
    .Q(\design_top.IOMUX[3][8] ),
    .CLK(clknet_leaf_349_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25002_ (.D(_05879_),
    .Q(\design_top.IOMUX[3][9] ),
    .CLK(clknet_leaf_348_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25003_ (.D(_05880_),
    .Q(\design_top.IOMUX[3][10] ),
    .CLK(clknet_leaf_348_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25004_ (.D(_05881_),
    .Q(\design_top.IOMUX[3][11] ),
    .CLK(clknet_leaf_349_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25005_ (.D(_05882_),
    .Q(\design_top.IOMUX[3][12] ),
    .CLK(clknet_leaf_349_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25006_ (.D(_05883_),
    .Q(\design_top.IOMUX[3][13] ),
    .CLK(clknet_leaf_345_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25007_ (.D(_05884_),
    .Q(\design_top.IOMUX[3][14] ),
    .CLK(clknet_leaf_345_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25008_ (.D(_05885_),
    .Q(\design_top.IOMUX[3][15] ),
    .CLK(clknet_leaf_345_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25009_ (.D(_05886_),
    .Q(\design_top.IOMUX[3][16] ),
    .CLK(clknet_leaf_344_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25010_ (.D(_05887_),
    .Q(\design_top.IOMUX[3][17] ),
    .CLK(clknet_leaf_344_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25011_ (.D(_05888_),
    .Q(\design_top.IOMUX[3][18] ),
    .CLK(clknet_leaf_372_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25012_ (.D(_05889_),
    .Q(\design_top.IOMUX[3][19] ),
    .CLK(clknet_leaf_372_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25013_ (.D(_05890_),
    .Q(\design_top.IOMUX[3][20] ),
    .CLK(clknet_leaf_372_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25014_ (.D(_05891_),
    .Q(\design_top.IOMUX[3][21] ),
    .CLK(clknet_leaf_372_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25015_ (.D(_05892_),
    .Q(\design_top.IOMUX[3][22] ),
    .CLK(clknet_leaf_371_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25016_ (.D(_05893_),
    .Q(\design_top.IOMUX[3][23] ),
    .CLK(clknet_leaf_372_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25017_ (.D(_05894_),
    .Q(\design_top.IOMUX[3][24] ),
    .CLK(clknet_leaf_371_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25018_ (.D(_05895_),
    .Q(\design_top.IOMUX[3][25] ),
    .CLK(clknet_leaf_371_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25019_ (.D(_05896_),
    .Q(\design_top.IOMUX[3][26] ),
    .CLK(clknet_leaf_371_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25020_ (.D(_05897_),
    .Q(\design_top.IOMUX[3][27] ),
    .CLK(clknet_leaf_371_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25021_ (.D(_05898_),
    .Q(\design_top.IOMUX[3][28] ),
    .CLK(clknet_leaf_371_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25022_ (.D(_05899_),
    .Q(\design_top.IOMUX[3][29] ),
    .CLK(clknet_leaf_371_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25023_ (.D(_05900_),
    .Q(\design_top.IOMUX[3][30] ),
    .CLK(clknet_leaf_371_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25024_ (.D(_05901_),
    .Q(\design_top.IOMUX[3][31] ),
    .CLK(clknet_leaf_371_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25025_ (.D(_05902_),
    .Q(\design_top.MEM[55][8] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25026_ (.D(_05903_),
    .Q(\design_top.MEM[55][9] ),
    .CLK(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25027_ (.D(_05904_),
    .Q(\design_top.MEM[55][10] ),
    .CLK(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25028_ (.D(_05905_),
    .Q(\design_top.MEM[55][11] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25029_ (.D(_05906_),
    .Q(\design_top.MEM[55][12] ),
    .CLK(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25030_ (.D(_05907_),
    .Q(\design_top.MEM[55][13] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25031_ (.D(_05908_),
    .Q(\design_top.MEM[55][14] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25032_ (.D(_05909_),
    .Q(\design_top.MEM[55][15] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25033_ (.D(_05910_),
    .Q(\design_top.MEM[56][24] ),
    .CLK(clknet_leaf_387_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25034_ (.D(_05911_),
    .Q(\design_top.MEM[56][25] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25035_ (.D(_05912_),
    .Q(\design_top.MEM[56][26] ),
    .CLK(clknet_leaf_314_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25036_ (.D(_05913_),
    .Q(\design_top.MEM[56][27] ),
    .CLK(clknet_leaf_382_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25037_ (.D(_05914_),
    .Q(\design_top.MEM[56][28] ),
    .CLK(clknet_leaf_378_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25038_ (.D(_05915_),
    .Q(\design_top.MEM[56][29] ),
    .CLK(clknet_leaf_378_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25039_ (.D(_05916_),
    .Q(\design_top.MEM[56][30] ),
    .CLK(clknet_leaf_378_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25040_ (.D(_05917_),
    .Q(\design_top.MEM[56][31] ),
    .CLK(clknet_leaf_381_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25041_ (.D(_05918_),
    .Q(\design_top.MEM[56][16] ),
    .CLK(clknet_leaf_155_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25042_ (.D(_05919_),
    .Q(\design_top.MEM[56][17] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25043_ (.D(_05920_),
    .Q(\design_top.MEM[56][18] ),
    .CLK(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25044_ (.D(_05921_),
    .Q(\design_top.MEM[56][19] ),
    .CLK(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25045_ (.D(_05922_),
    .Q(\design_top.MEM[56][20] ),
    .CLK(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25046_ (.D(_05923_),
    .Q(\design_top.MEM[56][21] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25047_ (.D(_05924_),
    .Q(\design_top.MEM[56][22] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25048_ (.D(_05925_),
    .Q(\design_top.MEM[56][23] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25049_ (.D(_05926_),
    .Q(\design_top.MEM[56][8] ),
    .CLK(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25050_ (.D(_05927_),
    .Q(\design_top.MEM[56][9] ),
    .CLK(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25051_ (.D(_05928_),
    .Q(\design_top.MEM[56][10] ),
    .CLK(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25052_ (.D(_05929_),
    .Q(\design_top.MEM[56][11] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25053_ (.D(_05930_),
    .Q(\design_top.MEM[56][12] ),
    .CLK(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25054_ (.D(_05931_),
    .Q(\design_top.MEM[56][13] ),
    .CLK(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25055_ (.D(_05932_),
    .Q(\design_top.MEM[56][14] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25056_ (.D(_05933_),
    .Q(\design_top.MEM[56][15] ),
    .CLK(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25057_ (.D(_05934_),
    .Q(\design_top.MEM[57][24] ),
    .CLK(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25058_ (.D(_05935_),
    .Q(\design_top.MEM[57][25] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25059_ (.D(_05936_),
    .Q(\design_top.MEM[57][26] ),
    .CLK(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25060_ (.D(_05937_),
    .Q(\design_top.MEM[57][27] ),
    .CLK(clknet_leaf_380_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25061_ (.D(_05938_),
    .Q(\design_top.MEM[57][28] ),
    .CLK(clknet_leaf_378_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25062_ (.D(_05939_),
    .Q(\design_top.MEM[57][29] ),
    .CLK(clknet_leaf_378_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25063_ (.D(_05940_),
    .Q(\design_top.MEM[57][30] ),
    .CLK(clknet_leaf_378_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25064_ (.D(_05941_),
    .Q(\design_top.MEM[57][31] ),
    .CLK(clknet_leaf_382_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25065_ (.D(_05942_),
    .Q(\design_top.MEM[57][16] ),
    .CLK(clknet_leaf_155_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25066_ (.D(_05943_),
    .Q(\design_top.MEM[57][17] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25067_ (.D(_05944_),
    .Q(\design_top.MEM[57][18] ),
    .CLK(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25068_ (.D(_05945_),
    .Q(\design_top.MEM[57][19] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25069_ (.D(_05946_),
    .Q(\design_top.MEM[57][20] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25070_ (.D(_05947_),
    .Q(\design_top.MEM[57][21] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25071_ (.D(_05948_),
    .Q(\design_top.MEM[57][22] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25072_ (.D(_05949_),
    .Q(\design_top.MEM[57][23] ),
    .CLK(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25073_ (.D(_05950_),
    .Q(\design_top.MEM[57][8] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25074_ (.D(_05951_),
    .Q(\design_top.MEM[57][9] ),
    .CLK(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25075_ (.D(_05952_),
    .Q(\design_top.MEM[57][10] ),
    .CLK(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25076_ (.D(_05953_),
    .Q(\design_top.MEM[57][11] ),
    .CLK(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25077_ (.D(_05954_),
    .Q(\design_top.MEM[57][12] ),
    .CLK(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25078_ (.D(_05955_),
    .Q(\design_top.MEM[57][13] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25079_ (.D(_05956_),
    .Q(\design_top.MEM[57][14] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25080_ (.D(_05957_),
    .Q(\design_top.MEM[57][15] ),
    .CLK(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25081_ (.D(_05958_),
    .Q(\design_top.MEM[58][24] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25082_ (.D(_05959_),
    .Q(\design_top.MEM[58][25] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25083_ (.D(_05960_),
    .Q(\design_top.MEM[58][26] ),
    .CLK(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25084_ (.D(_05961_),
    .Q(\design_top.MEM[58][27] ),
    .CLK(clknet_leaf_376_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25085_ (.D(_05962_),
    .Q(\design_top.MEM[58][28] ),
    .CLK(clknet_leaf_378_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25086_ (.D(_05963_),
    .Q(\design_top.MEM[58][29] ),
    .CLK(clknet_leaf_378_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25087_ (.D(_05964_),
    .Q(\design_top.MEM[58][30] ),
    .CLK(clknet_leaf_378_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25088_ (.D(_05965_),
    .Q(\design_top.MEM[58][31] ),
    .CLK(clknet_leaf_382_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25089_ (.D(_05966_),
    .Q(\design_top.MEM[58][16] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25090_ (.D(_05967_),
    .Q(\design_top.MEM[58][17] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25091_ (.D(_05968_),
    .Q(\design_top.MEM[58][18] ),
    .CLK(clknet_leaf_155_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25092_ (.D(_05969_),
    .Q(\design_top.MEM[58][19] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25093_ (.D(_05970_),
    .Q(\design_top.MEM[58][20] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25094_ (.D(_05971_),
    .Q(\design_top.MEM[58][21] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25095_ (.D(_05972_),
    .Q(\design_top.MEM[58][22] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25096_ (.D(_05973_),
    .Q(\design_top.MEM[58][23] ),
    .CLK(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25097_ (.D(_05974_),
    .Q(\design_top.MEM[58][8] ),
    .CLK(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25098_ (.D(_05975_),
    .Q(\design_top.MEM[58][9] ),
    .CLK(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25099_ (.D(_05976_),
    .Q(\design_top.MEM[58][10] ),
    .CLK(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25100_ (.D(_05977_),
    .Q(\design_top.MEM[58][11] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25101_ (.D(_05978_),
    .Q(\design_top.MEM[58][12] ),
    .CLK(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25102_ (.D(_05979_),
    .Q(\design_top.MEM[58][13] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25103_ (.D(_05980_),
    .Q(\design_top.MEM[58][14] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25104_ (.D(_05981_),
    .Q(\design_top.MEM[58][15] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25105_ (.D(_05982_),
    .Q(\design_top.MEM[59][24] ),
    .CLK(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25106_ (.D(_05983_),
    .Q(\design_top.MEM[59][25] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25107_ (.D(_05984_),
    .Q(\design_top.MEM[59][26] ),
    .CLK(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25108_ (.D(_05985_),
    .Q(\design_top.MEM[59][27] ),
    .CLK(clknet_leaf_375_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25109_ (.D(_05986_),
    .Q(\design_top.MEM[59][28] ),
    .CLK(clknet_leaf_380_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25110_ (.D(_05987_),
    .Q(\design_top.MEM[59][29] ),
    .CLK(clknet_leaf_378_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25111_ (.D(_05988_),
    .Q(\design_top.MEM[59][30] ),
    .CLK(clknet_leaf_376_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25112_ (.D(_05989_),
    .Q(\design_top.MEM[59][31] ),
    .CLK(clknet_leaf_381_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25113_ (.D(_05990_),
    .Q(\design_top.MEM[59][16] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25114_ (.D(_05991_),
    .Q(\design_top.MEM[59][17] ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25115_ (.D(_05992_),
    .Q(\design_top.MEM[59][18] ),
    .CLK(clknet_leaf_155_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25116_ (.D(_05993_),
    .Q(\design_top.MEM[59][19] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25117_ (.D(_05994_),
    .Q(\design_top.MEM[59][20] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25118_ (.D(_05995_),
    .Q(\design_top.MEM[59][21] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25119_ (.D(_05996_),
    .Q(\design_top.MEM[59][22] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25120_ (.D(_05997_),
    .Q(\design_top.MEM[59][23] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25121_ (.D(_05998_),
    .Q(\design_top.MEM[59][8] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25122_ (.D(_05999_),
    .Q(\design_top.MEM[59][9] ),
    .CLK(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25123_ (.D(_06000_),
    .Q(\design_top.MEM[59][10] ),
    .CLK(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25124_ (.D(_06001_),
    .Q(\design_top.MEM[59][11] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25125_ (.D(_06002_),
    .Q(\design_top.MEM[59][12] ),
    .CLK(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25126_ (.D(_06003_),
    .Q(\design_top.MEM[59][13] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25127_ (.D(_06004_),
    .Q(\design_top.MEM[59][14] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25128_ (.D(_06005_),
    .Q(\design_top.MEM[59][15] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25129_ (.D(_06006_),
    .Q(\design_top.MEM[5][8] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25130_ (.D(_06007_),
    .Q(\design_top.MEM[5][9] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25131_ (.D(_06008_),
    .Q(\design_top.MEM[5][10] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25132_ (.D(_06009_),
    .Q(\design_top.MEM[5][11] ),
    .CLK(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25133_ (.D(_06010_),
    .Q(\design_top.MEM[5][12] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25134_ (.D(_06011_),
    .Q(\design_top.MEM[5][13] ),
    .CLK(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25135_ (.D(_06012_),
    .Q(\design_top.MEM[5][14] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25136_ (.D(_06013_),
    .Q(\design_top.MEM[5][15] ),
    .CLK(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25137_ (.D(_06014_),
    .Q(\design_top.MEM[5][16] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25138_ (.D(_06015_),
    .Q(\design_top.MEM[5][17] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25139_ (.D(_06016_),
    .Q(\design_top.MEM[5][18] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25140_ (.D(_06017_),
    .Q(\design_top.MEM[5][19] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25141_ (.D(_06018_),
    .Q(\design_top.MEM[5][20] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25142_ (.D(_06019_),
    .Q(\design_top.MEM[5][21] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25143_ (.D(_06020_),
    .Q(\design_top.MEM[5][22] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25144_ (.D(_06021_),
    .Q(\design_top.MEM[5][23] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25145_ (.D(_06022_),
    .Q(\design_top.MEM[5][24] ),
    .CLK(clknet_leaf_387_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25146_ (.D(_06023_),
    .Q(\design_top.MEM[5][25] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25147_ (.D(_06024_),
    .Q(\design_top.MEM[5][26] ),
    .CLK(clknet_leaf_386_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25148_ (.D(_06025_),
    .Q(\design_top.MEM[5][27] ),
    .CLK(clknet_leaf_381_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25149_ (.D(_06026_),
    .Q(\design_top.MEM[5][28] ),
    .CLK(clknet_leaf_381_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25150_ (.D(_06027_),
    .Q(\design_top.MEM[5][29] ),
    .CLK(clknet_leaf_380_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25151_ (.D(_06028_),
    .Q(\design_top.MEM[5][30] ),
    .CLK(clknet_leaf_380_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25152_ (.D(_06029_),
    .Q(\design_top.MEM[5][31] ),
    .CLK(clknet_leaf_380_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25153_ (.D(_06030_),
    .Q(\design_top.MEM[60][24] ),
    .CLK(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25154_ (.D(_06031_),
    .Q(\design_top.MEM[60][25] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25155_ (.D(_06032_),
    .Q(\design_top.MEM[60][26] ),
    .CLK(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25156_ (.D(_06033_),
    .Q(\design_top.MEM[60][27] ),
    .CLK(clknet_leaf_384_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25157_ (.D(_06034_),
    .Q(\design_top.MEM[60][28] ),
    .CLK(clknet_leaf_381_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25158_ (.D(_06035_),
    .Q(\design_top.MEM[60][29] ),
    .CLK(clknet_leaf_382_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25159_ (.D(_06036_),
    .Q(\design_top.MEM[60][30] ),
    .CLK(clknet_leaf_382_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25160_ (.D(_06037_),
    .Q(\design_top.MEM[60][31] ),
    .CLK(clknet_leaf_384_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25161_ (.D(_06038_),
    .Q(\design_top.MEM[60][16] ),
    .CLK(clknet_leaf_172_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25162_ (.D(_06039_),
    .Q(\design_top.MEM[60][17] ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25163_ (.D(_06040_),
    .Q(\design_top.MEM[60][18] ),
    .CLK(clknet_leaf_155_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25164_ (.D(_06041_),
    .Q(\design_top.MEM[60][19] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25165_ (.D(_06042_),
    .Q(\design_top.MEM[60][20] ),
    .CLK(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25166_ (.D(_06043_),
    .Q(\design_top.MEM[60][21] ),
    .CLK(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25167_ (.D(_06044_),
    .Q(\design_top.MEM[60][22] ),
    .CLK(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25168_ (.D(_06045_),
    .Q(\design_top.MEM[60][23] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25169_ (.D(_06046_),
    .Q(\design_top.MEM[60][8] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25170_ (.D(_06047_),
    .Q(\design_top.MEM[60][9] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25171_ (.D(_06048_),
    .Q(\design_top.MEM[60][10] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25172_ (.D(_06049_),
    .Q(\design_top.MEM[60][11] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25173_ (.D(_06050_),
    .Q(\design_top.MEM[60][12] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25174_ (.D(_06051_),
    .Q(\design_top.MEM[60][13] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25175_ (.D(_06052_),
    .Q(\design_top.MEM[60][14] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25176_ (.D(_06053_),
    .Q(\design_top.MEM[60][15] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25177_ (.D(_06054_),
    .Q(\design_top.MEM[61][24] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25178_ (.D(_06055_),
    .Q(\design_top.MEM[61][25] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25179_ (.D(_06056_),
    .Q(\design_top.MEM[61][26] ),
    .CLK(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25180_ (.D(_06057_),
    .Q(\design_top.MEM[61][27] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25181_ (.D(_06058_),
    .Q(\design_top.MEM[61][28] ),
    .CLK(clknet_leaf_384_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25182_ (.D(_06059_),
    .Q(\design_top.MEM[61][29] ),
    .CLK(clknet_leaf_383_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25183_ (.D(_06060_),
    .Q(\design_top.MEM[61][30] ),
    .CLK(clknet_leaf_383_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25184_ (.D(_06061_),
    .Q(\design_top.MEM[61][31] ),
    .CLK(clknet_leaf_384_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25185_ (.D(_06062_),
    .Q(\design_top.MEM[61][16] ),
    .CLK(clknet_leaf_172_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25186_ (.D(_06063_),
    .Q(\design_top.MEM[61][17] ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25187_ (.D(_06064_),
    .Q(\design_top.MEM[61][18] ),
    .CLK(clknet_leaf_155_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25188_ (.D(_06065_),
    .Q(\design_top.MEM[61][19] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25189_ (.D(_06066_),
    .Q(\design_top.MEM[61][20] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25190_ (.D(_06067_),
    .Q(\design_top.MEM[61][21] ),
    .CLK(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25191_ (.D(_06068_),
    .Q(\design_top.MEM[61][22] ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25192_ (.D(_06069_),
    .Q(\design_top.MEM[61][23] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25193_ (.D(_06070_),
    .Q(\design_top.MEM[61][8] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25194_ (.D(_06071_),
    .Q(\design_top.MEM[61][9] ),
    .CLK(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25195_ (.D(_06072_),
    .Q(\design_top.MEM[61][10] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25196_ (.D(_06073_),
    .Q(\design_top.MEM[61][11] ),
    .CLK(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25197_ (.D(_06074_),
    .Q(\design_top.MEM[61][12] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25198_ (.D(_06075_),
    .Q(\design_top.MEM[61][13] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25199_ (.D(_06076_),
    .Q(\design_top.MEM[61][14] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25200_ (.D(_06077_),
    .Q(\design_top.MEM[61][15] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25201_ (.D(_06078_),
    .Q(\design_top.MEM[62][24] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25202_ (.D(_06079_),
    .Q(\design_top.MEM[62][25] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25203_ (.D(_06080_),
    .Q(\design_top.MEM[62][26] ),
    .CLK(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25204_ (.D(_06081_),
    .Q(\design_top.MEM[62][27] ),
    .CLK(clknet_leaf_383_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25205_ (.D(_06082_),
    .Q(\design_top.MEM[62][28] ),
    .CLK(clknet_leaf_385_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25206_ (.D(_06083_),
    .Q(\design_top.MEM[62][29] ),
    .CLK(clknet_leaf_383_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25207_ (.D(_06084_),
    .Q(\design_top.MEM[62][30] ),
    .CLK(clknet_leaf_383_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25208_ (.D(_06085_),
    .Q(\design_top.MEM[62][31] ),
    .CLK(clknet_leaf_384_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25209_ (.D(_06086_),
    .Q(\design_top.MEM[62][16] ),
    .CLK(clknet_leaf_172_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25210_ (.D(_06087_),
    .Q(\design_top.MEM[62][17] ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25211_ (.D(_06088_),
    .Q(\design_top.MEM[62][18] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25212_ (.D(_06089_),
    .Q(\design_top.MEM[62][19] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25213_ (.D(_06090_),
    .Q(\design_top.MEM[62][20] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25214_ (.D(_06091_),
    .Q(\design_top.MEM[62][21] ),
    .CLK(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25215_ (.D(_06092_),
    .Q(\design_top.MEM[62][22] ),
    .CLK(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25216_ (.D(_06093_),
    .Q(\design_top.MEM[62][23] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25217_ (.D(_06094_),
    .Q(\design_top.MEM[62][8] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25218_ (.D(_06095_),
    .Q(\design_top.MEM[62][9] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25219_ (.D(_06096_),
    .Q(\design_top.MEM[62][10] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25220_ (.D(_06097_),
    .Q(\design_top.MEM[62][11] ),
    .CLK(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25221_ (.D(_06098_),
    .Q(\design_top.MEM[62][12] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25222_ (.D(_06099_),
    .Q(\design_top.MEM[62][13] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25223_ (.D(_06100_),
    .Q(\design_top.MEM[62][14] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25224_ (.D(_06101_),
    .Q(\design_top.MEM[62][15] ),
    .CLK(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25225_ (.D(_06102_),
    .Q(\design_top.MEM[63][24] ),
    .CLK(clknet_leaf_314_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25226_ (.D(_06103_),
    .Q(\design_top.MEM[63][25] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25227_ (.D(_06104_),
    .Q(\design_top.MEM[63][26] ),
    .CLK(clknet_leaf_386_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25228_ (.D(_06105_),
    .Q(\design_top.MEM[63][27] ),
    .CLK(clknet_leaf_385_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25229_ (.D(_06106_),
    .Q(\design_top.MEM[63][28] ),
    .CLK(clknet_leaf_381_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25230_ (.D(_06107_),
    .Q(\design_top.MEM[63][29] ),
    .CLK(clknet_leaf_381_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25231_ (.D(_06108_),
    .Q(\design_top.MEM[63][30] ),
    .CLK(clknet_leaf_385_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25232_ (.D(_06109_),
    .Q(\design_top.MEM[63][31] ),
    .CLK(clknet_leaf_385_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25233_ (.D(_06110_),
    .Q(\design_top.MEM[63][16] ),
    .CLK(clknet_leaf_172_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25234_ (.D(_06111_),
    .Q(\design_top.MEM[63][17] ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25235_ (.D(_06112_),
    .Q(\design_top.MEM[63][18] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25236_ (.D(_06113_),
    .Q(\design_top.MEM[63][19] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25237_ (.D(_06114_),
    .Q(\design_top.MEM[63][20] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25238_ (.D(_06115_),
    .Q(\design_top.MEM[63][21] ),
    .CLK(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25239_ (.D(_06116_),
    .Q(\design_top.MEM[63][22] ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25240_ (.D(_06117_),
    .Q(\design_top.MEM[63][23] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25241_ (.D(_06118_),
    .Q(\design_top.MEM[63][8] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25242_ (.D(_06119_),
    .Q(\design_top.MEM[63][9] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25243_ (.D(_06120_),
    .Q(\design_top.MEM[63][10] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25244_ (.D(_06121_),
    .Q(\design_top.MEM[63][11] ),
    .CLK(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25245_ (.D(_06122_),
    .Q(\design_top.MEM[63][12] ),
    .CLK(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25246_ (.D(_06123_),
    .Q(\design_top.MEM[63][13] ),
    .CLK(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25247_ (.D(_06124_),
    .Q(\design_top.MEM[63][14] ),
    .CLK(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25248_ (.D(_06125_),
    .Q(\design_top.MEM[63][15] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25249_ (.D(_06126_),
    .Q(\design_top.MEM[6][8] ),
    .CLK(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25250_ (.D(_06127_),
    .Q(\design_top.MEM[6][9] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25251_ (.D(_06128_),
    .Q(\design_top.MEM[6][10] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25252_ (.D(_06129_),
    .Q(\design_top.MEM[6][11] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25253_ (.D(_06130_),
    .Q(\design_top.MEM[6][12] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25254_ (.D(_06131_),
    .Q(\design_top.MEM[6][13] ),
    .CLK(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25255_ (.D(_06132_),
    .Q(\design_top.MEM[6][14] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25256_ (.D(_06133_),
    .Q(\design_top.MEM[6][15] ),
    .CLK(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25257_ (.D(_06134_),
    .Q(\design_top.MEM[6][16] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25258_ (.D(_06135_),
    .Q(\design_top.MEM[6][17] ),
    .CLK(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25259_ (.D(_06136_),
    .Q(\design_top.MEM[6][18] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25260_ (.D(_06137_),
    .Q(\design_top.MEM[6][19] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25261_ (.D(_06138_),
    .Q(\design_top.MEM[6][20] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25262_ (.D(_06139_),
    .Q(\design_top.MEM[6][21] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25263_ (.D(_06140_),
    .Q(\design_top.MEM[6][22] ),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25264_ (.D(_06141_),
    .Q(\design_top.MEM[6][23] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25265_ (.D(_06142_),
    .Q(\design_top.MEM[6][24] ),
    .CLK(clknet_leaf_387_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25266_ (.D(_06143_),
    .Q(\design_top.MEM[6][25] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25267_ (.D(_06144_),
    .Q(\design_top.MEM[6][26] ),
    .CLK(clknet_leaf_387_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25268_ (.D(_06145_),
    .Q(\design_top.MEM[6][27] ),
    .CLK(clknet_leaf_385_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25269_ (.D(_06146_),
    .Q(\design_top.MEM[6][28] ),
    .CLK(clknet_leaf_393_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25270_ (.D(_06147_),
    .Q(\design_top.MEM[6][29] ),
    .CLK(clknet_leaf_381_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25271_ (.D(_06148_),
    .Q(\design_top.MEM[6][30] ),
    .CLK(clknet_leaf_381_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25272_ (.D(_06149_),
    .Q(\design_top.MEM[6][31] ),
    .CLK(clknet_leaf_389_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25273_ (.D(_06150_),
    .Q(\design_top.MEM[7][8] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25274_ (.D(_06151_),
    .Q(\design_top.MEM[7][9] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25275_ (.D(_06152_),
    .Q(\design_top.MEM[7][10] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25276_ (.D(_06153_),
    .Q(\design_top.MEM[7][11] ),
    .CLK(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25277_ (.D(_06154_),
    .Q(\design_top.MEM[7][12] ),
    .CLK(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25278_ (.D(_06155_),
    .Q(\design_top.MEM[7][13] ),
    .CLK(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25279_ (.D(_06156_),
    .Q(\design_top.MEM[7][14] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25280_ (.D(_06157_),
    .Q(\design_top.MEM[7][15] ),
    .CLK(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25281_ (.D(_06158_),
    .Q(\design_top.MEM[7][16] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25282_ (.D(_06159_),
    .Q(\design_top.MEM[7][17] ),
    .CLK(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25283_ (.D(_06160_),
    .Q(\design_top.MEM[7][18] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25284_ (.D(_06161_),
    .Q(\design_top.MEM[7][19] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25285_ (.D(_06162_),
    .Q(\design_top.MEM[7][20] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25286_ (.D(_06163_),
    .Q(\design_top.MEM[7][21] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25287_ (.D(_06164_),
    .Q(\design_top.MEM[7][22] ),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25288_ (.D(_06165_),
    .Q(\design_top.MEM[7][23] ),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25289_ (.D(_06166_),
    .Q(\design_top.MEM[7][24] ),
    .CLK(clknet_leaf_387_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25290_ (.D(_06167_),
    .Q(\design_top.MEM[7][25] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25291_ (.D(_06168_),
    .Q(\design_top.MEM[7][26] ),
    .CLK(clknet_leaf_387_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25292_ (.D(_06169_),
    .Q(\design_top.MEM[7][27] ),
    .CLK(clknet_leaf_381_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25293_ (.D(_06170_),
    .Q(\design_top.MEM[7][28] ),
    .CLK(clknet_leaf_393_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25294_ (.D(_06171_),
    .Q(\design_top.MEM[7][29] ),
    .CLK(clknet_leaf_381_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25295_ (.D(_06172_),
    .Q(\design_top.MEM[7][30] ),
    .CLK(clknet_leaf_380_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25296_ (.D(_06173_),
    .Q(\design_top.MEM[7][31] ),
    .CLK(clknet_leaf_393_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25297_ (.D(_06174_),
    .Q(\design_top.MEM[8][8] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25298_ (.D(_06175_),
    .Q(\design_top.MEM[8][9] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25299_ (.D(_06176_),
    .Q(\design_top.MEM[8][10] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25300_ (.D(_06177_),
    .Q(\design_top.MEM[8][11] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25301_ (.D(_06178_),
    .Q(\design_top.MEM[8][12] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25302_ (.D(_06179_),
    .Q(\design_top.MEM[8][13] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25303_ (.D(_06180_),
    .Q(\design_top.MEM[8][14] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25304_ (.D(_06181_),
    .Q(\design_top.MEM[8][15] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25305_ (.D(_06182_),
    .Q(\design_top.MEM[8][16] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25306_ (.D(_06183_),
    .Q(\design_top.MEM[8][17] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25307_ (.D(_06184_),
    .Q(\design_top.MEM[8][18] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25308_ (.D(_06185_),
    .Q(\design_top.MEM[8][19] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25309_ (.D(_06186_),
    .Q(\design_top.MEM[8][20] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25310_ (.D(_06187_),
    .Q(\design_top.MEM[8][21] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25311_ (.D(_06188_),
    .Q(\design_top.MEM[8][22] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25312_ (.D(_06189_),
    .Q(\design_top.MEM[8][23] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25313_ (.D(_06190_),
    .Q(\design_top.MEM[8][24] ),
    .CLK(clknet_leaf_388_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25314_ (.D(_06191_),
    .Q(\design_top.MEM[8][25] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25315_ (.D(_06192_),
    .Q(\design_top.MEM[8][26] ),
    .CLK(clknet_leaf_388_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25316_ (.D(_06193_),
    .Q(\design_top.MEM[8][27] ),
    .CLK(clknet_leaf_379_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25317_ (.D(_06194_),
    .Q(\design_top.MEM[8][28] ),
    .CLK(clknet_leaf_395_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25318_ (.D(_06195_),
    .Q(\design_top.MEM[8][29] ),
    .CLK(clknet_leaf_379_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25319_ (.D(_06196_),
    .Q(\design_top.MEM[8][30] ),
    .CLK(clknet_leaf_379_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25320_ (.D(_06197_),
    .Q(\design_top.MEM[8][31] ),
    .CLK(clknet_leaf_393_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25321_ (.D(_06198_),
    .Q(\design_top.MEM[9][8] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25322_ (.D(_06199_),
    .Q(\design_top.MEM[9][9] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25323_ (.D(_06200_),
    .Q(\design_top.MEM[9][10] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25324_ (.D(_06201_),
    .Q(\design_top.MEM[9][11] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25325_ (.D(_06202_),
    .Q(\design_top.MEM[9][12] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25326_ (.D(_06203_),
    .Q(\design_top.MEM[9][13] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25327_ (.D(_06204_),
    .Q(\design_top.MEM[9][14] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25328_ (.D(_06205_),
    .Q(\design_top.MEM[9][15] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25329_ (.D(_06206_),
    .Q(\design_top.MEM[9][16] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25330_ (.D(_06207_),
    .Q(\design_top.MEM[9][17] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25331_ (.D(_06208_),
    .Q(\design_top.MEM[9][18] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25332_ (.D(_06209_),
    .Q(\design_top.MEM[9][19] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25333_ (.D(_06210_),
    .Q(\design_top.MEM[9][20] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25334_ (.D(_06211_),
    .Q(\design_top.MEM[9][21] ),
    .CLK(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25335_ (.D(_06212_),
    .Q(\design_top.MEM[9][22] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25336_ (.D(_06213_),
    .Q(\design_top.MEM[9][23] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25337_ (.D(_06214_),
    .Q(\design_top.MEM[27][8] ),
    .CLK(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25338_ (.D(_06215_),
    .Q(\design_top.MEM[27][9] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25339_ (.D(_06216_),
    .Q(\design_top.MEM[27][10] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25340_ (.D(_06217_),
    .Q(\design_top.MEM[27][11] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25341_ (.D(_06218_),
    .Q(\design_top.MEM[27][12] ),
    .CLK(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25342_ (.D(_06219_),
    .Q(\design_top.MEM[27][13] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25343_ (.D(_06220_),
    .Q(\design_top.MEM[27][14] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25344_ (.D(_06221_),
    .Q(\design_top.MEM[27][15] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25345_ (.D(_06222_),
    .Q(\design_top.MEM[26][24] ),
    .CLK(clknet_leaf_396_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25346_ (.D(_06223_),
    .Q(\design_top.MEM[26][25] ),
    .CLK(clknet_leaf_398_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25347_ (.D(_06224_),
    .Q(\design_top.MEM[26][26] ),
    .CLK(clknet_leaf_389_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25348_ (.D(_06225_),
    .Q(\design_top.MEM[26][27] ),
    .CLK(clknet_leaf_410_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25349_ (.D(_06226_),
    .Q(\design_top.MEM[26][28] ),
    .CLK(clknet_leaf_410_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25350_ (.D(_06227_),
    .Q(\design_top.MEM[26][29] ),
    .CLK(clknet_leaf_411_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25351_ (.D(_06228_),
    .Q(\design_top.MEM[26][30] ),
    .CLK(clknet_leaf_409_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25352_ (.D(_06229_),
    .Q(\design_top.MEM[26][31] ),
    .CLK(clknet_leaf_409_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25353_ (.D(_06230_),
    .Q(\design_top.MEM[26][16] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25354_ (.D(_06231_),
    .Q(\design_top.MEM[26][17] ),
    .CLK(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25355_ (.D(_06232_),
    .Q(\design_top.MEM[26][18] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25356_ (.D(_06233_),
    .Q(\design_top.MEM[26][19] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25357_ (.D(_06234_),
    .Q(\design_top.MEM[26][20] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25358_ (.D(_06235_),
    .Q(\design_top.MEM[26][21] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25359_ (.D(_06236_),
    .Q(\design_top.MEM[26][22] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25360_ (.D(_06237_),
    .Q(\design_top.MEM[26][23] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25361_ (.D(_06238_),
    .Q(\design_top.MEM[26][8] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25362_ (.D(_06239_),
    .Q(\design_top.MEM[26][9] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25363_ (.D(_06240_),
    .Q(\design_top.MEM[26][10] ),
    .CLK(clknet_leaf_48_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25364_ (.D(_06241_),
    .Q(\design_top.MEM[26][11] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25365_ (.D(_06242_),
    .Q(\design_top.MEM[26][12] ),
    .CLK(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25366_ (.D(_06243_),
    .Q(\design_top.MEM[26][13] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25367_ (.D(_06244_),
    .Q(\design_top.MEM[26][14] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25368_ (.D(_06245_),
    .Q(\design_top.MEM[26][15] ),
    .CLK(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25369_ (.D(_06246_),
    .Q(\design_top.MEM[25][24] ),
    .CLK(clknet_leaf_398_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25370_ (.D(_06247_),
    .Q(\design_top.MEM[25][25] ),
    .CLK(clknet_leaf_401_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25371_ (.D(_06248_),
    .Q(\design_top.MEM[25][26] ),
    .CLK(clknet_leaf_392_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25372_ (.D(_06249_),
    .Q(\design_top.MEM[25][27] ),
    .CLK(clknet_leaf_411_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25373_ (.D(_06250_),
    .Q(\design_top.MEM[25][28] ),
    .CLK(clknet_leaf_414_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25374_ (.D(_06251_),
    .Q(\design_top.MEM[25][29] ),
    .CLK(clknet_leaf_414_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25375_ (.D(_06252_),
    .Q(\design_top.MEM[25][30] ),
    .CLK(clknet_leaf_411_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25376_ (.D(_06253_),
    .Q(\design_top.MEM[25][31] ),
    .CLK(clknet_leaf_410_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25377_ (.D(_06254_),
    .Q(\design_top.MEM[25][16] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25378_ (.D(_06255_),
    .Q(\design_top.MEM[25][17] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25379_ (.D(_06256_),
    .Q(\design_top.MEM[25][18] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25380_ (.D(_06257_),
    .Q(\design_top.MEM[25][19] ),
    .CLK(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25381_ (.D(_06258_),
    .Q(\design_top.MEM[25][20] ),
    .CLK(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25382_ (.D(_06259_),
    .Q(\design_top.MEM[25][21] ),
    .CLK(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25383_ (.D(_06260_),
    .Q(\design_top.MEM[25][22] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25384_ (.D(_06261_),
    .Q(\design_top.MEM[25][23] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25385_ (.D(_06262_),
    .Q(\design_top.MEM[20][24] ),
    .CLK(clknet_leaf_398_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25386_ (.D(_06263_),
    .Q(\design_top.MEM[20][25] ),
    .CLK(clknet_leaf_401_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25387_ (.D(_06264_),
    .Q(\design_top.MEM[20][26] ),
    .CLK(clknet_leaf_392_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25388_ (.D(_06265_),
    .Q(\design_top.MEM[20][27] ),
    .CLK(clknet_leaf_411_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25389_ (.D(_06266_),
    .Q(\design_top.MEM[20][28] ),
    .CLK(clknet_leaf_415_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25390_ (.D(_06267_),
    .Q(\design_top.MEM[20][29] ),
    .CLK(clknet_leaf_414_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25391_ (.D(_06268_),
    .Q(\design_top.MEM[20][30] ),
    .CLK(clknet_leaf_411_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25392_ (.D(_06269_),
    .Q(\design_top.MEM[20][31] ),
    .CLK(clknet_leaf_410_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25393_ (.D(_06270_),
    .Q(\design_top.MEM[38][16] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25394_ (.D(_06271_),
    .Q(\design_top.MEM[38][17] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25395_ (.D(_06272_),
    .Q(\design_top.MEM[38][18] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25396_ (.D(_06273_),
    .Q(\design_top.MEM[38][19] ),
    .CLK(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25397_ (.D(_06274_),
    .Q(\design_top.MEM[38][20] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25398_ (.D(_06275_),
    .Q(\design_top.MEM[38][21] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25399_ (.D(_06276_),
    .Q(\design_top.MEM[38][22] ),
    .CLK(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25400_ (.D(_06277_),
    .Q(\design_top.MEM[38][23] ),
    .CLK(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25401_ (.D(_06278_),
    .Q(\design_top.MEM[25][8] ),
    .CLK(clknet_leaf_48_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25402_ (.D(_06279_),
    .Q(\design_top.MEM[25][9] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25403_ (.D(_06280_),
    .Q(\design_top.MEM[25][10] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25404_ (.D(_06281_),
    .Q(\design_top.MEM[25][11] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25405_ (.D(_06282_),
    .Q(\design_top.MEM[25][12] ),
    .CLK(clknet_leaf_29_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25406_ (.D(_06283_),
    .Q(\design_top.MEM[25][13] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25407_ (.D(_06284_),
    .Q(\design_top.MEM[25][14] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25408_ (.D(_06285_),
    .Q(\design_top.MEM[25][15] ),
    .CLK(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25409_ (.D(_06286_),
    .Q(\design_top.MEM[24][24] ),
    .CLK(clknet_leaf_398_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25410_ (.D(_06287_),
    .Q(\design_top.MEM[24][25] ),
    .CLK(clknet_leaf_398_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25411_ (.D(_06288_),
    .Q(\design_top.MEM[24][26] ),
    .CLK(clknet_leaf_392_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25412_ (.D(_06289_),
    .Q(\design_top.MEM[24][27] ),
    .CLK(clknet_leaf_411_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25413_ (.D(_06290_),
    .Q(\design_top.MEM[24][28] ),
    .CLK(clknet_leaf_414_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25414_ (.D(_06291_),
    .Q(\design_top.MEM[24][29] ),
    .CLK(clknet_leaf_414_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25415_ (.D(_06292_),
    .Q(\design_top.MEM[24][30] ),
    .CLK(clknet_leaf_411_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25416_ (.D(_06293_),
    .Q(\design_top.MEM[24][31] ),
    .CLK(clknet_leaf_409_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25417_ (.D(_06294_),
    .Q(\design_top.MEM[24][16] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25418_ (.D(_06295_),
    .Q(\design_top.MEM[24][17] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25419_ (.D(_06296_),
    .Q(\design_top.MEM[24][18] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25420_ (.D(_06297_),
    .Q(\design_top.MEM[24][19] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25421_ (.D(_06298_),
    .Q(\design_top.MEM[24][20] ),
    .CLK(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25422_ (.D(_06299_),
    .Q(\design_top.MEM[24][21] ),
    .CLK(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25423_ (.D(_06300_),
    .Q(\design_top.MEM[24][22] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25424_ (.D(_06301_),
    .Q(\design_top.MEM[24][23] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25425_ (.D(_06302_),
    .Q(\design_top.MEM[38][8] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25426_ (.D(_06303_),
    .Q(\design_top.MEM[38][9] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25427_ (.D(_06304_),
    .Q(\design_top.MEM[38][10] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25428_ (.D(_06305_),
    .Q(\design_top.MEM[38][11] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25429_ (.D(_06306_),
    .Q(\design_top.MEM[38][12] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25430_ (.D(_06307_),
    .Q(\design_top.MEM[38][13] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25431_ (.D(_06308_),
    .Q(\design_top.MEM[38][14] ),
    .CLK(clknet_leaf_84_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25432_ (.D(_06309_),
    .Q(\design_top.MEM[38][15] ),
    .CLK(clknet_leaf_84_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25433_ (.D(_06310_),
    .Q(\design_top.MEM[24][8] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25434_ (.D(_06311_),
    .Q(\design_top.MEM[24][9] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25435_ (.D(_06312_),
    .Q(\design_top.MEM[24][10] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25436_ (.D(_06313_),
    .Q(\design_top.MEM[24][11] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25437_ (.D(_06314_),
    .Q(\design_top.MEM[24][12] ),
    .CLK(clknet_leaf_29_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25438_ (.D(_06315_),
    .Q(\design_top.MEM[24][13] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25439_ (.D(_06316_),
    .Q(\design_top.MEM[24][14] ),
    .CLK(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25440_ (.D(_06317_),
    .Q(\design_top.MEM[24][15] ),
    .CLK(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25441_ (.D(_06318_),
    .Q(\design_top.MEM[23][24] ),
    .CLK(clknet_leaf_399_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25442_ (.D(_06319_),
    .Q(\design_top.MEM[23][25] ),
    .CLK(clknet_leaf_401_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25443_ (.D(_06320_),
    .Q(\design_top.MEM[23][26] ),
    .CLK(clknet_leaf_393_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25444_ (.D(_06321_),
    .Q(\design_top.MEM[23][27] ),
    .CLK(clknet_leaf_411_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25445_ (.D(_06322_),
    .Q(\design_top.MEM[23][28] ),
    .CLK(clknet_leaf_415_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25446_ (.D(_06323_),
    .Q(\design_top.MEM[23][29] ),
    .CLK(clknet_leaf_415_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25447_ (.D(_06324_),
    .Q(\design_top.MEM[23][30] ),
    .CLK(clknet_leaf_411_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25448_ (.D(_06325_),
    .Q(\design_top.MEM[23][31] ),
    .CLK(clknet_leaf_410_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25449_ (.D(_06326_),
    .Q(\design_top.MEM[37][24] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25450_ (.D(_06327_),
    .Q(\design_top.MEM[37][25] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25451_ (.D(_06328_),
    .Q(\design_top.MEM[37][26] ),
    .CLK(clknet_leaf_386_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25452_ (.D(_06329_),
    .Q(\design_top.MEM[37][27] ),
    .CLK(clknet_leaf_361_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25453_ (.D(_06330_),
    .Q(\design_top.MEM[37][28] ),
    .CLK(clknet_leaf_357_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25454_ (.D(_06331_),
    .Q(\design_top.MEM[37][29] ),
    .CLK(clknet_leaf_357_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25455_ (.D(_06332_),
    .Q(\design_top.MEM[37][30] ),
    .CLK(clknet_leaf_358_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25456_ (.D(_06333_),
    .Q(\design_top.MEM[37][31] ),
    .CLK(clknet_leaf_362_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25457_ (.D(_06334_),
    .Q(\design_top.MEM[37][16] ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25458_ (.D(_06335_),
    .Q(\design_top.MEM[37][17] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25459_ (.D(_06336_),
    .Q(\design_top.MEM[37][18] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25460_ (.D(_06337_),
    .Q(\design_top.MEM[37][19] ),
    .CLK(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25461_ (.D(_06338_),
    .Q(\design_top.MEM[37][20] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25462_ (.D(_06339_),
    .Q(\design_top.MEM[37][21] ),
    .CLK(clknet_leaf_143_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25463_ (.D(_06340_),
    .Q(\design_top.MEM[37][22] ),
    .CLK(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25464_ (.D(_06341_),
    .Q(\design_top.MEM[37][23] ),
    .CLK(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25465_ (.D(_06342_),
    .Q(\design_top.MEM[23][16] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25466_ (.D(_06343_),
    .Q(\design_top.MEM[23][17] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25467_ (.D(_06344_),
    .Q(\design_top.MEM[23][18] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25468_ (.D(_06345_),
    .Q(\design_top.MEM[23][19] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25469_ (.D(_06346_),
    .Q(\design_top.MEM[23][20] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25470_ (.D(_06347_),
    .Q(\design_top.MEM[23][21] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25471_ (.D(_06348_),
    .Q(\design_top.MEM[23][22] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25472_ (.D(_06349_),
    .Q(\design_top.MEM[23][23] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25473_ (.D(_06350_),
    .Q(\design_top.MEM[37][8] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25474_ (.D(_06351_),
    .Q(\design_top.MEM[37][9] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25475_ (.D(_06352_),
    .Q(\design_top.MEM[37][10] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25476_ (.D(_06353_),
    .Q(\design_top.MEM[37][11] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25477_ (.D(_06354_),
    .Q(\design_top.MEM[37][12] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25478_ (.D(_06355_),
    .Q(\design_top.MEM[37][13] ),
    .CLK(clknet_leaf_84_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25479_ (.D(_06356_),
    .Q(\design_top.MEM[37][14] ),
    .CLK(clknet_leaf_84_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25480_ (.D(_06357_),
    .Q(\design_top.MEM[37][15] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25481_ (.D(_06358_),
    .Q(\design_top.MEM[23][8] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25482_ (.D(_06359_),
    .Q(\design_top.MEM[23][9] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25483_ (.D(_06360_),
    .Q(\design_top.MEM[23][10] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25484_ (.D(_06361_),
    .Q(\design_top.MEM[23][11] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25485_ (.D(_06362_),
    .Q(\design_top.MEM[23][12] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25486_ (.D(_06363_),
    .Q(\design_top.MEM[23][13] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25487_ (.D(_06364_),
    .Q(\design_top.MEM[23][14] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25488_ (.D(_06365_),
    .Q(\design_top.MEM[23][15] ),
    .CLK(clknet_leaf_31_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25489_ (.D(_06366_),
    .Q(\design_top.MEM[22][24] ),
    .CLK(clknet_leaf_392_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25490_ (.D(_06367_),
    .Q(\design_top.MEM[22][25] ),
    .CLK(clknet_leaf_400_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25491_ (.D(_06368_),
    .Q(\design_top.MEM[22][26] ),
    .CLK(clknet_leaf_389_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25492_ (.D(_06369_),
    .Q(\design_top.MEM[22][27] ),
    .CLK(clknet_leaf_362_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25493_ (.D(_06370_),
    .Q(\design_top.MEM[22][28] ),
    .CLK(clknet_leaf_357_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25494_ (.D(_06371_),
    .Q(\design_top.MEM[22][29] ),
    .CLK(clknet_leaf_415_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25495_ (.D(_06372_),
    .Q(\design_top.MEM[22][30] ),
    .CLK(clknet_leaf_358_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25496_ (.D(_06373_),
    .Q(\design_top.MEM[22][31] ),
    .CLK(clknet_leaf_410_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25497_ (.D(_06374_),
    .Q(\design_top.MEM[1][8] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25498_ (.D(_06375_),
    .Q(\design_top.MEM[1][9] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25499_ (.D(_06376_),
    .Q(\design_top.MEM[1][10] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25500_ (.D(_06377_),
    .Q(\design_top.MEM[1][11] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25501_ (.D(_06378_),
    .Q(\design_top.MEM[1][12] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25502_ (.D(_06379_),
    .Q(\design_top.MEM[1][13] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25503_ (.D(_06380_),
    .Q(\design_top.MEM[1][14] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25504_ (.D(_06381_),
    .Q(\design_top.MEM[1][15] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25505_ (.D(_06382_),
    .Q(\design_top.MEM[1][16] ),
    .CLK(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25506_ (.D(_06383_),
    .Q(\design_top.MEM[1][17] ),
    .CLK(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25507_ (.D(_06384_),
    .Q(\design_top.MEM[1][18] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25508_ (.D(_06385_),
    .Q(\design_top.MEM[1][19] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25509_ (.D(_06386_),
    .Q(\design_top.MEM[1][20] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25510_ (.D(_06387_),
    .Q(\design_top.MEM[1][21] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25511_ (.D(_06388_),
    .Q(\design_top.MEM[1][22] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25512_ (.D(_06389_),
    .Q(\design_top.MEM[1][23] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25513_ (.D(_06390_),
    .Q(\design_top.MEM[1][24] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25514_ (.D(_06391_),
    .Q(\design_top.MEM[1][25] ),
    .CLK(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25515_ (.D(_06392_),
    .Q(\design_top.MEM[1][26] ),
    .CLK(clknet_leaf_388_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25516_ (.D(_06393_),
    .Q(\design_top.MEM[1][27] ),
    .CLK(clknet_leaf_364_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25517_ (.D(_06394_),
    .Q(\design_top.MEM[1][28] ),
    .CLK(clknet_leaf_363_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25518_ (.D(_06395_),
    .Q(\design_top.MEM[1][29] ),
    .CLK(clknet_leaf_363_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25519_ (.D(_06396_),
    .Q(\design_top.MEM[1][30] ),
    .CLK(clknet_leaf_364_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25520_ (.D(_06397_),
    .Q(\design_top.MEM[1][31] ),
    .CLK(clknet_leaf_409_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25521_ (.D(_06398_),
    .Q(\design_top.MEM[45][8] ),
    .CLK(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25522_ (.D(_06399_),
    .Q(\design_top.MEM[45][9] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25523_ (.D(_06400_),
    .Q(\design_top.MEM[45][10] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25524_ (.D(_06401_),
    .Q(\design_top.MEM[45][11] ),
    .CLK(clknet_leaf_76_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25525_ (.D(_06402_),
    .Q(\design_top.MEM[45][12] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25526_ (.D(_06403_),
    .Q(\design_top.MEM[45][13] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25527_ (.D(_06404_),
    .Q(\design_top.MEM[45][14] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25528_ (.D(_06405_),
    .Q(\design_top.MEM[45][15] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25529_ (.D(_06406_),
    .Q(\design_top.MEM[44][24] ),
    .CLK(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25530_ (.D(_06407_),
    .Q(\design_top.MEM[44][25] ),
    .CLK(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25531_ (.D(_06408_),
    .Q(\design_top.MEM[44][26] ),
    .CLK(clknet_leaf_384_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25532_ (.D(_06409_),
    .Q(\design_top.MEM[44][27] ),
    .CLK(clknet_leaf_360_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25533_ (.D(_06410_),
    .Q(\design_top.MEM[44][28] ),
    .CLK(clknet_leaf_358_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25534_ (.D(_06411_),
    .Q(\design_top.MEM[44][29] ),
    .CLK(clknet_leaf_359_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25535_ (.D(_06412_),
    .Q(\design_top.MEM[44][30] ),
    .CLK(clknet_leaf_358_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25536_ (.D(_06413_),
    .Q(\design_top.MEM[44][31] ),
    .CLK(clknet_leaf_361_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25537_ (.D(_06414_),
    .Q(\design_top.MEM[44][16] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25538_ (.D(_06415_),
    .Q(\design_top.MEM[44][17] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25539_ (.D(_06416_),
    .Q(\design_top.MEM[44][18] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25540_ (.D(_06417_),
    .Q(\design_top.MEM[44][19] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25541_ (.D(_06418_),
    .Q(\design_top.MEM[44][20] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25542_ (.D(_06419_),
    .Q(\design_top.MEM[44][21] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25543_ (.D(_06420_),
    .Q(\design_top.MEM[44][22] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25544_ (.D(_06421_),
    .Q(\design_top.MEM[44][23] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25545_ (.D(_06422_),
    .Q(\design_top.MEM[44][8] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25546_ (.D(_06423_),
    .Q(\design_top.MEM[44][9] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25547_ (.D(_06424_),
    .Q(\design_top.MEM[44][10] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25548_ (.D(_06425_),
    .Q(\design_top.MEM[44][11] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25549_ (.D(_06426_),
    .Q(\design_top.MEM[44][12] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25550_ (.D(_06427_),
    .Q(\design_top.MEM[44][13] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25551_ (.D(_06428_),
    .Q(\design_top.MEM[44][14] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25552_ (.D(_06429_),
    .Q(\design_top.MEM[44][15] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25553_ (.D(_06430_),
    .Q(\design_top.MEM[50][16] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25554_ (.D(_06431_),
    .Q(\design_top.MEM[50][17] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25555_ (.D(_06432_),
    .Q(\design_top.MEM[50][18] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25556_ (.D(_06433_),
    .Q(\design_top.MEM[50][19] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25557_ (.D(_06434_),
    .Q(\design_top.MEM[50][20] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25558_ (.D(_06435_),
    .Q(\design_top.MEM[50][21] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25559_ (.D(_06436_),
    .Q(\design_top.MEM[50][22] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25560_ (.D(_06437_),
    .Q(\design_top.MEM[50][23] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25561_ (.D(_06438_),
    .Q(\design_top.MEM[43][24] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25562_ (.D(_06439_),
    .Q(\design_top.MEM[43][25] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25563_ (.D(_06440_),
    .Q(\design_top.MEM[43][26] ),
    .CLK(clknet_leaf_315_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25564_ (.D(_06441_),
    .Q(\design_top.MEM[43][27] ),
    .CLK(clknet_leaf_360_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25565_ (.D(_06442_),
    .Q(\design_top.MEM[43][28] ),
    .CLK(clknet_leaf_354_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25566_ (.D(_06443_),
    .Q(\design_top.MEM[43][29] ),
    .CLK(clknet_leaf_353_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25567_ (.D(_06444_),
    .Q(\design_top.MEM[43][30] ),
    .CLK(clknet_leaf_360_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25568_ (.D(_06445_),
    .Q(\design_top.MEM[43][31] ),
    .CLK(clknet_leaf_367_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25569_ (.D(_06446_),
    .Q(\design_top.MEM[43][16] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25570_ (.D(_06447_),
    .Q(\design_top.MEM[43][17] ),
    .CLK(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25571_ (.D(_06448_),
    .Q(\design_top.MEM[43][18] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25572_ (.D(_06449_),
    .Q(\design_top.MEM[43][19] ),
    .CLK(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25573_ (.D(_06450_),
    .Q(\design_top.MEM[43][20] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25574_ (.D(_06451_),
    .Q(\design_top.MEM[43][21] ),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25575_ (.D(_06452_),
    .Q(\design_top.MEM[43][22] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25576_ (.D(_06453_),
    .Q(\design_top.MEM[43][23] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25577_ (.D(_06454_),
    .Q(\design_top.MEM[50][8] ),
    .CLK(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25578_ (.D(_06455_),
    .Q(\design_top.MEM[50][9] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25579_ (.D(_06456_),
    .Q(\design_top.MEM[50][10] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25580_ (.D(_06457_),
    .Q(\design_top.MEM[50][11] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25581_ (.D(_06458_),
    .Q(\design_top.MEM[50][12] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25582_ (.D(_06459_),
    .Q(\design_top.MEM[50][13] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25583_ (.D(_06460_),
    .Q(\design_top.MEM[50][14] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25584_ (.D(_06461_),
    .Q(\design_top.MEM[50][15] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25585_ (.D(_06462_),
    .Q(\design_top.MEM[43][8] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25586_ (.D(_06463_),
    .Q(\design_top.MEM[43][9] ),
    .CLK(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25587_ (.D(_06464_),
    .Q(\design_top.MEM[43][10] ),
    .CLK(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25588_ (.D(_06465_),
    .Q(\design_top.MEM[43][11] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25589_ (.D(_06466_),
    .Q(\design_top.MEM[43][12] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25590_ (.D(_06467_),
    .Q(\design_top.MEM[43][13] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25591_ (.D(_06468_),
    .Q(\design_top.MEM[43][14] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25592_ (.D(_06469_),
    .Q(\design_top.MEM[43][15] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25593_ (.D(_06470_),
    .Q(\design_top.MEM[4][24] ),
    .CLK(clknet_leaf_387_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25594_ (.D(_06471_),
    .Q(\design_top.MEM[4][25] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25595_ (.D(_06472_),
    .Q(\design_top.MEM[4][26] ),
    .CLK(clknet_leaf_387_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25596_ (.D(_06473_),
    .Q(\design_top.MEM[4][27] ),
    .CLK(clknet_leaf_381_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25597_ (.D(_06474_),
    .Q(\design_top.MEM[4][28] ),
    .CLK(clknet_leaf_393_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25598_ (.D(_06475_),
    .Q(\design_top.MEM[4][29] ),
    .CLK(clknet_leaf_380_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25599_ (.D(_06476_),
    .Q(\design_top.MEM[4][30] ),
    .CLK(clknet_leaf_379_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25600_ (.D(_06477_),
    .Q(\design_top.MEM[4][31] ),
    .CLK(clknet_leaf_393_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25601_ (.D(_06478_),
    .Q(\design_top.MEM[4][16] ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25602_ (.D(_06479_),
    .Q(\design_top.MEM[4][17] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25603_ (.D(_06480_),
    .Q(\design_top.MEM[4][18] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25604_ (.D(_06481_),
    .Q(\design_top.MEM[4][19] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25605_ (.D(_06482_),
    .Q(\design_top.MEM[4][20] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25606_ (.D(_06483_),
    .Q(\design_top.MEM[4][21] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25607_ (.D(_06484_),
    .Q(\design_top.MEM[4][22] ),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25608_ (.D(_06485_),
    .Q(\design_top.MEM[4][23] ),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25609_ (.D(_06486_),
    .Q(\design_top.MEM[42][24] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25610_ (.D(_06487_),
    .Q(\design_top.MEM[42][25] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25611_ (.D(_06488_),
    .Q(\design_top.MEM[42][26] ),
    .CLK(clknet_leaf_315_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25612_ (.D(_06489_),
    .Q(\design_top.MEM[42][27] ),
    .CLK(clknet_leaf_360_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25613_ (.D(_06490_),
    .Q(\design_top.MEM[42][28] ),
    .CLK(clknet_leaf_354_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25614_ (.D(_06491_),
    .Q(\design_top.MEM[42][29] ),
    .CLK(clknet_leaf_353_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25615_ (.D(_06492_),
    .Q(\design_top.MEM[42][30] ),
    .CLK(clknet_leaf_353_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25616_ (.D(_06493_),
    .Q(\design_top.MEM[42][31] ),
    .CLK(clknet_leaf_360_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25617_ (.D(_06494_),
    .Q(\design_top.MEM[42][16] ),
    .CLK(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25618_ (.D(_06495_),
    .Q(\design_top.MEM[42][17] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25619_ (.D(_06496_),
    .Q(\design_top.MEM[42][18] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25620_ (.D(_06497_),
    .Q(\design_top.MEM[42][19] ),
    .CLK(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25621_ (.D(_06498_),
    .Q(\design_top.MEM[42][20] ),
    .CLK(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25622_ (.D(_06499_),
    .Q(\design_top.MEM[42][21] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25623_ (.D(_06500_),
    .Q(\design_top.MEM[42][22] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25624_ (.D(_06501_),
    .Q(\design_top.MEM[42][23] ),
    .CLK(clknet_leaf_143_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25625_ (.D(_06502_),
    .Q(\design_top.MEM[4][8] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25626_ (.D(_06503_),
    .Q(\design_top.MEM[4][9] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25627_ (.D(_06504_),
    .Q(\design_top.MEM[4][10] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25628_ (.D(_06505_),
    .Q(\design_top.MEM[4][11] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25629_ (.D(_06506_),
    .Q(\design_top.MEM[4][12] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25630_ (.D(_06507_),
    .Q(\design_top.MEM[4][13] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25631_ (.D(_06508_),
    .Q(\design_top.MEM[4][14] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25632_ (.D(_06509_),
    .Q(\design_top.MEM[4][15] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25633_ (.D(_06510_),
    .Q(\design_top.MEM[49][24] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25634_ (.D(_06511_),
    .Q(\design_top.MEM[49][25] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25635_ (.D(_06512_),
    .Q(\design_top.MEM[49][26] ),
    .CLK(clknet_leaf_314_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25636_ (.D(_06513_),
    .Q(\design_top.MEM[49][27] ),
    .CLK(clknet_leaf_365_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25637_ (.D(_06514_),
    .Q(\design_top.MEM[49][28] ),
    .CLK(clknet_leaf_363_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25638_ (.D(_06515_),
    .Q(\design_top.MEM[49][29] ),
    .CLK(clknet_leaf_366_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25639_ (.D(_06516_),
    .Q(\design_top.MEM[49][30] ),
    .CLK(clknet_leaf_366_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25640_ (.D(_06517_),
    .Q(\design_top.MEM[49][31] ),
    .CLK(clknet_leaf_365_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25641_ (.D(_06518_),
    .Q(\design_top.MEM[49][16] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25642_ (.D(_06519_),
    .Q(\design_top.MEM[49][17] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25643_ (.D(_06520_),
    .Q(\design_top.MEM[49][18] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25644_ (.D(_06521_),
    .Q(\design_top.MEM[49][19] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25645_ (.D(_06522_),
    .Q(\design_top.MEM[49][20] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25646_ (.D(_06523_),
    .Q(\design_top.MEM[49][21] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25647_ (.D(_06524_),
    .Q(\design_top.MEM[49][22] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25648_ (.D(_06525_),
    .Q(\design_top.MEM[49][23] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25649_ (.D(_06526_),
    .Q(\design_top.MEM[42][8] ),
    .CLK(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25650_ (.D(_06527_),
    .Q(\design_top.MEM[42][9] ),
    .CLK(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25651_ (.D(_06528_),
    .Q(\design_top.MEM[42][10] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25652_ (.D(_06529_),
    .Q(\design_top.MEM[42][11] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25653_ (.D(_06530_),
    .Q(\design_top.MEM[42][12] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25654_ (.D(_06531_),
    .Q(\design_top.MEM[42][13] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25655_ (.D(_06532_),
    .Q(\design_top.MEM[42][14] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25656_ (.D(_06533_),
    .Q(\design_top.MEM[42][15] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25657_ (.D(_06534_),
    .Q(\design_top.MEM[41][24] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25658_ (.D(_06535_),
    .Q(\design_top.MEM[41][25] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25659_ (.D(_06536_),
    .Q(\design_top.MEM[41][26] ),
    .CLK(clknet_leaf_315_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25660_ (.D(_06537_),
    .Q(\design_top.MEM[41][27] ),
    .CLK(clknet_leaf_368_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25661_ (.D(_06538_),
    .Q(\design_top.MEM[41][28] ),
    .CLK(clknet_leaf_354_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25662_ (.D(_06539_),
    .Q(\design_top.MEM[41][29] ),
    .CLK(clknet_leaf_354_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25663_ (.D(_06540_),
    .Q(\design_top.MEM[41][30] ),
    .CLK(clknet_leaf_353_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25664_ (.D(_06541_),
    .Q(\design_top.MEM[41][31] ),
    .CLK(clknet_leaf_368_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25665_ (.D(_06542_),
    .Q(\design_top.MEM[41][16] ),
    .CLK(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25666_ (.D(_06543_),
    .Q(\design_top.MEM[41][17] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25667_ (.D(_06544_),
    .Q(\design_top.MEM[41][18] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25668_ (.D(_06545_),
    .Q(\design_top.MEM[41][19] ),
    .CLK(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25669_ (.D(_06546_),
    .Q(\design_top.MEM[41][20] ),
    .CLK(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25670_ (.D(_06547_),
    .Q(\design_top.MEM[41][21] ),
    .CLK(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25671_ (.D(_06548_),
    .Q(\design_top.MEM[41][22] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25672_ (.D(_06549_),
    .Q(\design_top.MEM[41][23] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25673_ (.D(_06550_),
    .Q(\design_top.MEM[49][8] ),
    .CLK(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25674_ (.D(_06551_),
    .Q(\design_top.MEM[49][9] ),
    .CLK(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25675_ (.D(_06552_),
    .Q(\design_top.MEM[49][10] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25676_ (.D(_06553_),
    .Q(\design_top.MEM[49][11] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25677_ (.D(_06554_),
    .Q(\design_top.MEM[49][12] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25678_ (.D(_06555_),
    .Q(\design_top.MEM[49][13] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25679_ (.D(_06556_),
    .Q(\design_top.MEM[49][14] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25680_ (.D(_06557_),
    .Q(\design_top.MEM[49][15] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25681_ (.D(_06558_),
    .Q(\design_top.MEM[41][8] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25682_ (.D(_06559_),
    .Q(\design_top.MEM[41][9] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25683_ (.D(_06560_),
    .Q(\design_top.MEM[41][10] ),
    .CLK(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25684_ (.D(_06561_),
    .Q(\design_top.MEM[41][11] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25685_ (.D(_06562_),
    .Q(\design_top.MEM[41][12] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25686_ (.D(_06563_),
    .Q(\design_top.MEM[41][13] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25687_ (.D(_06564_),
    .Q(\design_top.MEM[41][14] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25688_ (.D(_06565_),
    .Q(\design_top.MEM[41][15] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25689_ (.D(_06566_),
    .Q(\design_top.MEM[48][24] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25690_ (.D(_06567_),
    .Q(\design_top.MEM[48][25] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25691_ (.D(_06568_),
    .Q(\design_top.MEM[48][26] ),
    .CLK(clknet_leaf_314_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25692_ (.D(_06569_),
    .Q(\design_top.MEM[48][27] ),
    .CLK(clknet_leaf_366_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25693_ (.D(_06570_),
    .Q(\design_top.MEM[48][28] ),
    .CLK(clknet_leaf_363_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25694_ (.D(_06571_),
    .Q(\design_top.MEM[48][29] ),
    .CLK(clknet_leaf_366_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25695_ (.D(_06572_),
    .Q(\design_top.MEM[48][30] ),
    .CLK(clknet_leaf_366_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25696_ (.D(_06573_),
    .Q(\design_top.MEM[48][31] ),
    .CLK(clknet_leaf_365_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25697_ (.D(_06574_),
    .Q(\design_top.MEM[48][16] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25698_ (.D(_06575_),
    .Q(\design_top.MEM[48][17] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25699_ (.D(_06576_),
    .Q(\design_top.MEM[48][18] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25700_ (.D(_06577_),
    .Q(\design_top.MEM[48][19] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25701_ (.D(_06578_),
    .Q(\design_top.MEM[48][20] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25702_ (.D(_06579_),
    .Q(\design_top.MEM[48][21] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25703_ (.D(_06580_),
    .Q(\design_top.MEM[48][22] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25704_ (.D(_06581_),
    .Q(\design_top.MEM[48][23] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25705_ (.D(_06582_),
    .Q(\design_top.MEM[40][24] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25706_ (.D(_06583_),
    .Q(\design_top.MEM[40][25] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25707_ (.D(_06584_),
    .Q(\design_top.MEM[40][26] ),
    .CLK(clknet_leaf_315_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25708_ (.D(_06585_),
    .Q(\design_top.MEM[40][27] ),
    .CLK(clknet_leaf_353_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25709_ (.D(_06586_),
    .Q(\design_top.MEM[40][28] ),
    .CLK(clknet_leaf_354_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25710_ (.D(_06587_),
    .Q(\design_top.MEM[40][29] ),
    .CLK(clknet_leaf_354_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25711_ (.D(_06588_),
    .Q(\design_top.MEM[40][30] ),
    .CLK(clknet_leaf_353_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25712_ (.D(_06589_),
    .Q(\design_top.MEM[40][31] ),
    .CLK(clknet_leaf_367_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25713_ (.D(_06590_),
    .Q(\design_top.MEM[40][16] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25714_ (.D(_06591_),
    .Q(\design_top.MEM[40][17] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25715_ (.D(_06592_),
    .Q(\design_top.MEM[40][18] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25716_ (.D(_06593_),
    .Q(\design_top.MEM[40][19] ),
    .CLK(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25717_ (.D(_06594_),
    .Q(\design_top.MEM[40][20] ),
    .CLK(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25718_ (.D(_06595_),
    .Q(\design_top.MEM[40][21] ),
    .CLK(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25719_ (.D(_06596_),
    .Q(\design_top.MEM[40][22] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25720_ (.D(_06597_),
    .Q(\design_top.MEM[40][23] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25721_ (.D(_06598_),
    .Q(\design_top.MEM[48][8] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25722_ (.D(_06599_),
    .Q(\design_top.MEM[48][9] ),
    .CLK(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25723_ (.D(_06600_),
    .Q(\design_top.MEM[48][10] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25724_ (.D(_06601_),
    .Q(\design_top.MEM[48][11] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25725_ (.D(_06602_),
    .Q(\design_top.MEM[48][12] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25726_ (.D(_06603_),
    .Q(\design_top.MEM[48][13] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25727_ (.D(_06604_),
    .Q(\design_top.MEM[48][14] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25728_ (.D(_06605_),
    .Q(\design_top.MEM[48][15] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25729_ (.D(_06606_),
    .Q(\design_top.MEM[40][8] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25730_ (.D(_06607_),
    .Q(\design_top.MEM[40][9] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25731_ (.D(_06608_),
    .Q(\design_top.MEM[40][10] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25732_ (.D(_06609_),
    .Q(\design_top.MEM[40][11] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25733_ (.D(_06610_),
    .Q(\design_top.MEM[40][12] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25734_ (.D(_06611_),
    .Q(\design_top.MEM[40][13] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25735_ (.D(_06612_),
    .Q(\design_top.MEM[40][14] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25736_ (.D(_06613_),
    .Q(\design_top.MEM[40][15] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25737_ (.D(_06614_),
    .Q(\design_top.MEM[47][24] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25738_ (.D(_06615_),
    .Q(\design_top.MEM[47][25] ),
    .CLK(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25739_ (.D(_06616_),
    .Q(\design_top.MEM[47][26] ),
    .CLK(clknet_leaf_386_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25740_ (.D(_06617_),
    .Q(\design_top.MEM[47][27] ),
    .CLK(clknet_leaf_361_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25741_ (.D(_06618_),
    .Q(\design_top.MEM[47][28] ),
    .CLK(clknet_leaf_357_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25742_ (.D(_06619_),
    .Q(\design_top.MEM[47][29] ),
    .CLK(clknet_leaf_359_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25743_ (.D(_06620_),
    .Q(\design_top.MEM[47][30] ),
    .CLK(clknet_leaf_358_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25744_ (.D(_06621_),
    .Q(\design_top.MEM[47][31] ),
    .CLK(clknet_leaf_361_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25745_ (.D(_06622_),
    .Q(\design_top.MEM[47][16] ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25746_ (.D(_06623_),
    .Q(\design_top.MEM[47][17] ),
    .CLK(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25747_ (.D(_06624_),
    .Q(\design_top.MEM[47][18] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25748_ (.D(_06625_),
    .Q(\design_top.MEM[47][19] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25749_ (.D(_06626_),
    .Q(\design_top.MEM[47][20] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25750_ (.D(_06627_),
    .Q(\design_top.MEM[47][21] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25751_ (.D(_06628_),
    .Q(\design_top.MEM[47][22] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25752_ (.D(_06629_),
    .Q(\design_top.MEM[47][23] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25753_ (.D(_06630_),
    .Q(\design_top.MEM[3][24] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25754_ (.D(_06631_),
    .Q(\design_top.MEM[3][25] ),
    .CLK(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25755_ (.D(_06632_),
    .Q(\design_top.MEM[3][26] ),
    .CLK(clknet_leaf_386_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25756_ (.D(_06633_),
    .Q(\design_top.MEM[3][27] ),
    .CLK(clknet_leaf_362_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25757_ (.D(_06634_),
    .Q(\design_top.MEM[3][28] ),
    .CLK(clknet_leaf_362_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25758_ (.D(_06635_),
    .Q(\design_top.MEM[3][29] ),
    .CLK(clknet_leaf_361_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25759_ (.D(_06636_),
    .Q(\design_top.MEM[3][30] ),
    .CLK(clknet_leaf_362_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25760_ (.D(_06637_),
    .Q(\design_top.MEM[3][31] ),
    .CLK(clknet_leaf_362_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25761_ (.D(_06638_),
    .Q(\design_top.MEM[3][16] ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25762_ (.D(_06639_),
    .Q(\design_top.MEM[3][17] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25763_ (.D(_06640_),
    .Q(\design_top.MEM[3][18] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25764_ (.D(_06641_),
    .Q(\design_top.MEM[3][19] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25765_ (.D(_06642_),
    .Q(\design_top.MEM[3][20] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25766_ (.D(_06643_),
    .Q(\design_top.MEM[3][21] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25767_ (.D(_06644_),
    .Q(\design_top.MEM[3][22] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25768_ (.D(_06645_),
    .Q(\design_top.MEM[3][23] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25769_ (.D(_06646_),
    .Q(\design_top.MEM[3][8] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25770_ (.D(_06647_),
    .Q(\design_top.MEM[3][9] ),
    .CLK(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25771_ (.D(_06648_),
    .Q(\design_top.MEM[3][10] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25772_ (.D(_06649_),
    .Q(\design_top.MEM[3][11] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25773_ (.D(_06650_),
    .Q(\design_top.MEM[3][12] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25774_ (.D(_06651_),
    .Q(\design_top.MEM[3][13] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25775_ (.D(_06652_),
    .Q(\design_top.MEM[3][14] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25776_ (.D(_06653_),
    .Q(\design_top.MEM[3][15] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25777_ (.D(_06654_),
    .Q(\design_top.MEM[47][8] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25778_ (.D(_06655_),
    .Q(\design_top.MEM[47][9] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25779_ (.D(_06656_),
    .Q(\design_top.MEM[47][10] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25780_ (.D(_06657_),
    .Q(\design_top.MEM[47][11] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25781_ (.D(_06658_),
    .Q(\design_top.MEM[47][12] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25782_ (.D(_06659_),
    .Q(\design_top.MEM[47][13] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25783_ (.D(_06660_),
    .Q(\design_top.MEM[47][14] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25784_ (.D(_06661_),
    .Q(\design_top.MEM[47][15] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25785_ (.D(_06662_),
    .Q(\design_top.MEM[39][24] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25786_ (.D(_06663_),
    .Q(\design_top.MEM[39][25] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25787_ (.D(_06664_),
    .Q(\design_top.MEM[39][26] ),
    .CLK(clknet_leaf_386_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25788_ (.D(_06665_),
    .Q(\design_top.MEM[39][27] ),
    .CLK(clknet_leaf_360_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25789_ (.D(_06666_),
    .Q(\design_top.MEM[39][28] ),
    .CLK(clknet_leaf_357_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25790_ (.D(_06667_),
    .Q(\design_top.MEM[39][29] ),
    .CLK(clknet_leaf_359_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25791_ (.D(_06668_),
    .Q(\design_top.MEM[39][30] ),
    .CLK(clknet_leaf_359_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25792_ (.D(_06669_),
    .Q(\design_top.MEM[39][31] ),
    .CLK(clknet_leaf_362_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25793_ (.D(_06670_),
    .Q(\design_top.MEM[46][24] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25794_ (.D(_06671_),
    .Q(\design_top.MEM[46][25] ),
    .CLK(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25795_ (.D(_06672_),
    .Q(\design_top.MEM[46][26] ),
    .CLK(clknet_leaf_386_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25796_ (.D(_06673_),
    .Q(\design_top.MEM[46][27] ),
    .CLK(clknet_leaf_361_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25797_ (.D(_06674_),
    .Q(\design_top.MEM[46][28] ),
    .CLK(clknet_leaf_357_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25798_ (.D(_06675_),
    .Q(\design_top.MEM[46][29] ),
    .CLK(clknet_leaf_357_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25799_ (.D(_06676_),
    .Q(\design_top.MEM[46][30] ),
    .CLK(clknet_leaf_358_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25800_ (.D(_06677_),
    .Q(\design_top.MEM[46][31] ),
    .CLK(clknet_leaf_362_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25801_ (.D(_06678_),
    .Q(\design_top.MEM[46][16] ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25802_ (.D(_06679_),
    .Q(\design_top.MEM[46][17] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25803_ (.D(_06680_),
    .Q(\design_top.MEM[46][18] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25804_ (.D(_06681_),
    .Q(\design_top.MEM[46][19] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25805_ (.D(_06682_),
    .Q(\design_top.MEM[46][20] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25806_ (.D(_06683_),
    .Q(\design_top.MEM[46][21] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25807_ (.D(_06684_),
    .Q(\design_top.MEM[46][22] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25808_ (.D(_06685_),
    .Q(\design_top.MEM[46][23] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25809_ (.D(_06686_),
    .Q(\design_top.MEM[39][16] ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25810_ (.D(_06687_),
    .Q(\design_top.MEM[39][17] ),
    .CLK(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25811_ (.D(_06688_),
    .Q(\design_top.MEM[39][18] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25812_ (.D(_06689_),
    .Q(\design_top.MEM[39][19] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25813_ (.D(_06690_),
    .Q(\design_top.MEM[39][20] ),
    .CLK(clknet_leaf_143_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25814_ (.D(_06691_),
    .Q(\design_top.MEM[39][21] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25815_ (.D(_06692_),
    .Q(\design_top.MEM[39][22] ),
    .CLK(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25816_ (.D(_06693_),
    .Q(\design_top.MEM[39][23] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25817_ (.D(_06694_),
    .Q(\design_top.MEM[46][8] ),
    .CLK(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25818_ (.D(_06695_),
    .Q(\design_top.MEM[46][9] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25819_ (.D(_06696_),
    .Q(\design_top.MEM[46][10] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25820_ (.D(_06697_),
    .Q(\design_top.MEM[46][11] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25821_ (.D(_06698_),
    .Q(\design_top.MEM[46][12] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25822_ (.D(_06699_),
    .Q(\design_top.MEM[46][13] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25823_ (.D(_06700_),
    .Q(\design_top.MEM[46][14] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25824_ (.D(_06701_),
    .Q(\design_top.MEM[46][15] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25825_ (.D(_06702_),
    .Q(\design_top.MEM[39][8] ),
    .CLK(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25826_ (.D(_06703_),
    .Q(\design_top.MEM[39][9] ),
    .CLK(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25827_ (.D(_06704_),
    .Q(\design_top.MEM[39][10] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25828_ (.D(_06705_),
    .Q(\design_top.MEM[39][11] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25829_ (.D(_06706_),
    .Q(\design_top.MEM[39][12] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25830_ (.D(_06707_),
    .Q(\design_top.MEM[39][13] ),
    .CLK(clknet_leaf_84_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25831_ (.D(_06708_),
    .Q(\design_top.MEM[39][14] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25832_ (.D(_06709_),
    .Q(\design_top.MEM[39][15] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25833_ (.D(_06710_),
    .Q(\design_top.MEM[45][24] ),
    .CLK(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25834_ (.D(_06711_),
    .Q(\design_top.MEM[45][25] ),
    .CLK(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25835_ (.D(_06712_),
    .Q(\design_top.MEM[45][26] ),
    .CLK(clknet_leaf_386_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25836_ (.D(_06713_),
    .Q(\design_top.MEM[45][27] ),
    .CLK(clknet_leaf_361_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25837_ (.D(_06714_),
    .Q(\design_top.MEM[45][28] ),
    .CLK(clknet_leaf_358_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25838_ (.D(_06715_),
    .Q(\design_top.MEM[45][29] ),
    .CLK(clknet_leaf_358_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25839_ (.D(_06716_),
    .Q(\design_top.MEM[45][30] ),
    .CLK(clknet_leaf_358_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25840_ (.D(_06717_),
    .Q(\design_top.MEM[45][31] ),
    .CLK(clknet_leaf_361_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25841_ (.D(_06718_),
    .Q(\design_top.MEM[38][24] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25842_ (.D(_06719_),
    .Q(\design_top.MEM[38][25] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25843_ (.D(_06720_),
    .Q(\design_top.MEM[38][26] ),
    .CLK(clknet_leaf_386_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25844_ (.D(_06721_),
    .Q(\design_top.MEM[38][27] ),
    .CLK(clknet_leaf_367_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25845_ (.D(_06722_),
    .Q(\design_top.MEM[38][28] ),
    .CLK(clknet_leaf_363_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25846_ (.D(_06723_),
    .Q(\design_top.MEM[38][29] ),
    .CLK(clknet_leaf_367_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25847_ (.D(_06724_),
    .Q(\design_top.MEM[38][30] ),
    .CLK(clknet_leaf_367_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25848_ (.D(_06725_),
    .Q(\design_top.MEM[38][31] ),
    .CLK(clknet_leaf_363_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25849_ (.D(_06726_),
    .Q(\design_top.MEM[53][8] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25850_ (.D(_06727_),
    .Q(\design_top.MEM[53][9] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25851_ (.D(_06728_),
    .Q(\design_top.MEM[53][10] ),
    .CLK(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25852_ (.D(_06729_),
    .Q(\design_top.MEM[53][11] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25853_ (.D(_06730_),
    .Q(\design_top.MEM[53][12] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25854_ (.D(_06731_),
    .Q(\design_top.MEM[53][13] ),
    .CLK(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25855_ (.D(_06732_),
    .Q(\design_top.MEM[53][14] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25856_ (.D(_06733_),
    .Q(\design_top.MEM[53][15] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25857_ (.D(_06734_),
    .Q(\design_top.MEM[53][24] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25858_ (.D(_06735_),
    .Q(\design_top.MEM[53][25] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25859_ (.D(_06736_),
    .Q(\design_top.MEM[53][26] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25860_ (.D(_06737_),
    .Q(\design_top.MEM[53][27] ),
    .CLK(clknet_leaf_375_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25861_ (.D(_06738_),
    .Q(\design_top.MEM[53][28] ),
    .CLK(clknet_leaf_377_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25862_ (.D(_06739_),
    .Q(\design_top.MEM[53][29] ),
    .CLK(clknet_leaf_377_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25863_ (.D(_06740_),
    .Q(\design_top.MEM[53][30] ),
    .CLK(clknet_leaf_376_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25864_ (.D(_06741_),
    .Q(\design_top.MEM[53][31] ),
    .CLK(clknet_leaf_375_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25865_ (.D(_06742_),
    .Q(\design_top.MEM[53][16] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25866_ (.D(_06743_),
    .Q(\design_top.MEM[53][17] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25867_ (.D(_06744_),
    .Q(\design_top.MEM[53][18] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25868_ (.D(_06745_),
    .Q(\design_top.MEM[53][19] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25869_ (.D(_06746_),
    .Q(\design_top.MEM[53][20] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25870_ (.D(_06747_),
    .Q(\design_top.MEM[53][21] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25871_ (.D(_06748_),
    .Q(\design_top.MEM[53][22] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25872_ (.D(_06749_),
    .Q(\design_top.MEM[53][23] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25873_ (.D(_06750_),
    .Q(\design_top.MEM[52][24] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25874_ (.D(_06751_),
    .Q(\design_top.MEM[52][25] ),
    .CLK(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25875_ (.D(_06752_),
    .Q(\design_top.MEM[52][26] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25876_ (.D(_06753_),
    .Q(\design_top.MEM[52][27] ),
    .CLK(clknet_leaf_375_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25877_ (.D(_06754_),
    .Q(\design_top.MEM[52][28] ),
    .CLK(clknet_leaf_377_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25878_ (.D(_06755_),
    .Q(\design_top.MEM[52][29] ),
    .CLK(clknet_leaf_373_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25879_ (.D(_06756_),
    .Q(\design_top.MEM[52][30] ),
    .CLK(clknet_leaf_374_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25880_ (.D(_06757_),
    .Q(\design_top.MEM[52][31] ),
    .CLK(clknet_leaf_375_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25881_ (.D(_06758_),
    .Q(\design_top.MEM[55][24] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25882_ (.D(_06759_),
    .Q(\design_top.MEM[55][25] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25883_ (.D(_06760_),
    .Q(\design_top.MEM[55][26] ),
    .CLK(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25884_ (.D(_06761_),
    .Q(\design_top.MEM[55][27] ),
    .CLK(clknet_leaf_375_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25885_ (.D(_06762_),
    .Q(\design_top.MEM[55][28] ),
    .CLK(clknet_leaf_377_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25886_ (.D(_06763_),
    .Q(\design_top.MEM[55][29] ),
    .CLK(clknet_leaf_377_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25887_ (.D(_06764_),
    .Q(\design_top.MEM[55][30] ),
    .CLK(clknet_leaf_374_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25888_ (.D(_06765_),
    .Q(\design_top.MEM[55][31] ),
    .CLK(clknet_leaf_375_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25889_ (.D(_06766_),
    .Q(\design_top.MEM[55][16] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25890_ (.D(_06767_),
    .Q(\design_top.MEM[55][17] ),
    .CLK(clknet_leaf_172_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25891_ (.D(_06768_),
    .Q(\design_top.MEM[55][18] ),
    .CLK(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25892_ (.D(_06769_),
    .Q(\design_top.MEM[55][19] ),
    .CLK(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25893_ (.D(_06770_),
    .Q(\design_top.MEM[55][20] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25894_ (.D(_06771_),
    .Q(\design_top.MEM[55][21] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25895_ (.D(_06772_),
    .Q(\design_top.MEM[55][22] ),
    .CLK(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25896_ (.D(_06773_),
    .Q(\design_top.MEM[55][23] ),
    .CLK(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25897_ (.D(_06774_),
    .Q(\design_top.MEM[52][16] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25898_ (.D(_06775_),
    .Q(\design_top.MEM[52][17] ),
    .CLK(clknet_leaf_172_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25899_ (.D(_06776_),
    .Q(\design_top.MEM[52][18] ),
    .CLK(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25900_ (.D(_06777_),
    .Q(\design_top.MEM[52][19] ),
    .CLK(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25901_ (.D(_06778_),
    .Q(\design_top.MEM[52][20] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25902_ (.D(_06779_),
    .Q(\design_top.MEM[52][21] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25903_ (.D(_06780_),
    .Q(\design_top.MEM[52][22] ),
    .CLK(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25904_ (.D(_06781_),
    .Q(\design_top.MEM[52][23] ),
    .CLK(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25905_ (.D(_06782_),
    .Q(\design_top.MEM[54][24] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25906_ (.D(_06783_),
    .Q(\design_top.MEM[54][25] ),
    .CLK(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25907_ (.D(_06784_),
    .Q(\design_top.MEM[54][26] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25908_ (.D(_06785_),
    .Q(\design_top.MEM[54][27] ),
    .CLK(clknet_leaf_375_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25909_ (.D(_06786_),
    .Q(\design_top.MEM[54][28] ),
    .CLK(clknet_leaf_377_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25910_ (.D(_06787_),
    .Q(\design_top.MEM[54][29] ),
    .CLK(clknet_leaf_377_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25911_ (.D(_06788_),
    .Q(\design_top.MEM[54][30] ),
    .CLK(clknet_leaf_376_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25912_ (.D(_06789_),
    .Q(\design_top.MEM[54][31] ),
    .CLK(clknet_leaf_383_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25913_ (.D(_06790_),
    .Q(\design_top.MEM[52][8] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25914_ (.D(_06791_),
    .Q(\design_top.MEM[52][9] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25915_ (.D(_06792_),
    .Q(\design_top.MEM[52][10] ),
    .CLK(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25916_ (.D(_06793_),
    .Q(\design_top.MEM[52][11] ),
    .CLK(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25917_ (.D(_06794_),
    .Q(\design_top.MEM[52][12] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25918_ (.D(_06795_),
    .Q(\design_top.MEM[52][13] ),
    .CLK(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25919_ (.D(_06796_),
    .Q(\design_top.MEM[52][14] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25920_ (.D(_06797_),
    .Q(\design_top.MEM[52][15] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25921_ (.D(_06798_),
    .Q(\design_top.MEM[54][16] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25922_ (.D(_06799_),
    .Q(\design_top.MEM[54][17] ),
    .CLK(clknet_leaf_172_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25923_ (.D(_06800_),
    .Q(\design_top.MEM[54][18] ),
    .CLK(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25924_ (.D(_06801_),
    .Q(\design_top.MEM[54][19] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25925_ (.D(_06802_),
    .Q(\design_top.MEM[54][20] ),
    .CLK(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25926_ (.D(_06803_),
    .Q(\design_top.MEM[54][21] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25927_ (.D(_06804_),
    .Q(\design_top.MEM[54][22] ),
    .CLK(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25928_ (.D(_06805_),
    .Q(\design_top.MEM[54][23] ),
    .CLK(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25929_ (.D(_06806_),
    .Q(\design_top.MEM[51][24] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25930_ (.D(_06807_),
    .Q(\design_top.MEM[51][25] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25931_ (.D(_06808_),
    .Q(\design_top.MEM[51][26] ),
    .CLK(clknet_leaf_314_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25932_ (.D(_06809_),
    .Q(\design_top.MEM[51][27] ),
    .CLK(clknet_leaf_365_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25933_ (.D(_06810_),
    .Q(\design_top.MEM[51][28] ),
    .CLK(clknet_leaf_364_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25934_ (.D(_06811_),
    .Q(\design_top.MEM[51][29] ),
    .CLK(clknet_leaf_367_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25935_ (.D(_06812_),
    .Q(\design_top.MEM[51][30] ),
    .CLK(clknet_leaf_365_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25936_ (.D(_06813_),
    .Q(\design_top.MEM[51][31] ),
    .CLK(clknet_leaf_364_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25937_ (.D(_06814_),
    .Q(\design_top.MEM[51][16] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25938_ (.D(_06815_),
    .Q(\design_top.MEM[51][17] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25939_ (.D(_06816_),
    .Q(\design_top.MEM[51][18] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25940_ (.D(_06817_),
    .Q(\design_top.MEM[51][19] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25941_ (.D(_06818_),
    .Q(\design_top.MEM[51][20] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25942_ (.D(_06819_),
    .Q(\design_top.MEM[51][21] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25943_ (.D(_06820_),
    .Q(\design_top.MEM[51][22] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25944_ (.D(_06821_),
    .Q(\design_top.MEM[51][23] ),
    .CLK(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25945_ (.D(_06822_),
    .Q(\design_top.MEM[51][8] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25946_ (.D(_06823_),
    .Q(\design_top.MEM[51][9] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25947_ (.D(_06824_),
    .Q(\design_top.MEM[51][10] ),
    .CLK(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25948_ (.D(_06825_),
    .Q(\design_top.MEM[51][11] ),
    .CLK(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25949_ (.D(_06826_),
    .Q(\design_top.MEM[51][12] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25950_ (.D(_06827_),
    .Q(\design_top.MEM[51][13] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25951_ (.D(_06828_),
    .Q(\design_top.MEM[51][14] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25952_ (.D(_06829_),
    .Q(\design_top.MEM[51][15] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25953_ (.D(_06830_),
    .Q(\design_top.MEM[54][8] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25954_ (.D(_06831_),
    .Q(\design_top.MEM[54][9] ),
    .CLK(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25955_ (.D(_06832_),
    .Q(\design_top.MEM[54][10] ),
    .CLK(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25956_ (.D(_06833_),
    .Q(\design_top.MEM[54][11] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25957_ (.D(_06834_),
    .Q(\design_top.MEM[54][12] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25958_ (.D(_06835_),
    .Q(\design_top.MEM[54][13] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25959_ (.D(_06836_),
    .Q(\design_top.MEM[54][14] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25960_ (.D(_06837_),
    .Q(\design_top.MEM[54][15] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25961_ (.D(_06838_),
    .Q(\design_top.MEM[50][24] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25962_ (.D(_06839_),
    .Q(\design_top.MEM[50][25] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25963_ (.D(_06840_),
    .Q(\design_top.MEM[50][26] ),
    .CLK(clknet_leaf_314_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25964_ (.D(_06841_),
    .Q(\design_top.MEM[50][27] ),
    .CLK(clknet_leaf_365_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25965_ (.D(_06842_),
    .Q(\design_top.MEM[50][28] ),
    .CLK(clknet_leaf_364_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25966_ (.D(_06843_),
    .Q(\design_top.MEM[50][29] ),
    .CLK(clknet_leaf_365_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25967_ (.D(_06844_),
    .Q(\design_top.MEM[50][30] ),
    .CLK(clknet_leaf_366_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25968_ (.D(_06845_),
    .Q(\design_top.MEM[50][31] ),
    .CLK(clknet_leaf_364_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25969_ (.D(_06846_),
    .Q(\design_top.MEM[36][24] ),
    .CLK(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25970_ (.D(_06847_),
    .Q(\design_top.MEM[36][25] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25971_ (.D(_06848_),
    .Q(\design_top.MEM[36][26] ),
    .CLK(clknet_leaf_386_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25972_ (.D(_06849_),
    .Q(\design_top.MEM[36][27] ),
    .CLK(clknet_leaf_360_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25973_ (.D(_06850_),
    .Q(\design_top.MEM[36][28] ),
    .CLK(clknet_leaf_356_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25974_ (.D(_06851_),
    .Q(\design_top.MEM[36][29] ),
    .CLK(clknet_leaf_355_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25975_ (.D(_06852_),
    .Q(\design_top.MEM[36][30] ),
    .CLK(clknet_leaf_359_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25976_ (.D(_06853_),
    .Q(\design_top.MEM[36][31] ),
    .CLK(clknet_leaf_361_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25977_ (.D(_06854_),
    .Q(\design_top.MEM[36][16] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25978_ (.D(_06855_),
    .Q(\design_top.MEM[36][17] ),
    .CLK(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25979_ (.D(_06856_),
    .Q(\design_top.MEM[36][18] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25980_ (.D(_06857_),
    .Q(\design_top.MEM[36][19] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25981_ (.D(_06858_),
    .Q(\design_top.MEM[36][20] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25982_ (.D(_06859_),
    .Q(\design_top.MEM[36][21] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25983_ (.D(_06860_),
    .Q(\design_top.MEM[36][22] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25984_ (.D(_06861_),
    .Q(\design_top.MEM[36][23] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25985_ (.D(_06862_),
    .Q(\design_top.MEM[22][16] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25986_ (.D(_06863_),
    .Q(\design_top.MEM[22][17] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25987_ (.D(_06864_),
    .Q(\design_top.MEM[22][18] ),
    .CLK(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25988_ (.D(_06865_),
    .Q(\design_top.MEM[22][19] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25989_ (.D(_06866_),
    .Q(\design_top.MEM[22][20] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25990_ (.D(_06867_),
    .Q(\design_top.MEM[22][21] ),
    .CLK(clknet_5_20_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25991_ (.D(_06868_),
    .Q(\design_top.MEM[22][22] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25992_ (.D(_06869_),
    .Q(\design_top.MEM[22][23] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25993_ (.D(_06870_),
    .Q(\design_top.MEM[22][8] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25994_ (.D(_06871_),
    .Q(\design_top.MEM[22][9] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25995_ (.D(_06872_),
    .Q(\design_top.MEM[22][10] ),
    .CLK(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25996_ (.D(_06873_),
    .Q(\design_top.MEM[22][11] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25997_ (.D(_06874_),
    .Q(\design_top.MEM[22][12] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25998_ (.D(_06875_),
    .Q(\design_top.MEM[22][13] ),
    .CLK(clknet_leaf_31_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _25999_ (.D(_06876_),
    .Q(\design_top.MEM[22][14] ),
    .CLK(clknet_leaf_31_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26000_ (.D(_06877_),
    .Q(\design_top.MEM[22][15] ),
    .CLK(clknet_leaf_31_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26001_ (.D(_06878_),
    .Q(\design_top.MEM[21][24] ),
    .CLK(clknet_leaf_391_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26002_ (.D(_06879_),
    .Q(\design_top.MEM[21][25] ),
    .CLK(clknet_leaf_400_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26003_ (.D(_06880_),
    .Q(\design_top.MEM[21][26] ),
    .CLK(clknet_leaf_389_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26004_ (.D(_06881_),
    .Q(\design_top.MEM[21][27] ),
    .CLK(clknet_leaf_362_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26005_ (.D(_06882_),
    .Q(\design_top.MEM[21][28] ),
    .CLK(clknet_leaf_357_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26006_ (.D(_06883_),
    .Q(\design_top.MEM[21][29] ),
    .CLK(clknet_leaf_357_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26007_ (.D(_06884_),
    .Q(\design_top.MEM[21][30] ),
    .CLK(clknet_leaf_362_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26008_ (.D(_06885_),
    .Q(\design_top.MEM[21][31] ),
    .CLK(clknet_leaf_362_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26009_ (.D(_06886_),
    .Q(\design_top.MEM[36][8] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26010_ (.D(_06887_),
    .Q(\design_top.MEM[36][9] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26011_ (.D(_06888_),
    .Q(\design_top.MEM[36][10] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26012_ (.D(_06889_),
    .Q(\design_top.MEM[36][11] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26013_ (.D(_06890_),
    .Q(\design_top.MEM[36][12] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26014_ (.D(_06891_),
    .Q(\design_top.MEM[36][13] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26015_ (.D(_06892_),
    .Q(\design_top.MEM[36][14] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26016_ (.D(_06893_),
    .Q(\design_top.MEM[36][15] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26017_ (.D(_06894_),
    .Q(\design_top.MEM[21][16] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26018_ (.D(_06895_),
    .Q(\design_top.MEM[21][17] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26019_ (.D(_06896_),
    .Q(\design_top.MEM[21][18] ),
    .CLK(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26020_ (.D(_06897_),
    .Q(\design_top.MEM[21][19] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26021_ (.D(_06898_),
    .Q(\design_top.MEM[21][20] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26022_ (.D(_06899_),
    .Q(\design_top.MEM[21][21] ),
    .CLK(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26023_ (.D(_06900_),
    .Q(\design_top.MEM[21][22] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26024_ (.D(_06901_),
    .Q(\design_top.MEM[21][23] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26025_ (.D(_06902_),
    .Q(\design_top.MEM[21][8] ),
    .CLK(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26026_ (.D(_06903_),
    .Q(\design_top.MEM[21][9] ),
    .CLK(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26027_ (.D(_06904_),
    .Q(\design_top.MEM[21][10] ),
    .CLK(clknet_leaf_48_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26028_ (.D(_06905_),
    .Q(\design_top.MEM[21][11] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26029_ (.D(_06906_),
    .Q(\design_top.MEM[21][12] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26030_ (.D(_06907_),
    .Q(\design_top.MEM[21][13] ),
    .CLK(clknet_leaf_31_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26031_ (.D(_06908_),
    .Q(\design_top.MEM[21][14] ),
    .CLK(clknet_leaf_31_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26032_ (.D(_06909_),
    .Q(\design_top.MEM[21][15] ),
    .CLK(clknet_leaf_31_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26033_ (.D(_06910_),
    .Q(\design_top.MEM[20][16] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26034_ (.D(_06911_),
    .Q(\design_top.MEM[20][17] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26035_ (.D(_06912_),
    .Q(\design_top.MEM[20][18] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26036_ (.D(_06913_),
    .Q(\design_top.MEM[20][19] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26037_ (.D(_06914_),
    .Q(\design_top.MEM[20][20] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26038_ (.D(_06915_),
    .Q(\design_top.MEM[20][21] ),
    .CLK(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26039_ (.D(_06916_),
    .Q(\design_top.MEM[20][22] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26040_ (.D(_06917_),
    .Q(\design_top.MEM[20][23] ),
    .CLK(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26041_ (.D(_06918_),
    .Q(\design_top.MEM[35][24] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26042_ (.D(_06919_),
    .Q(\design_top.MEM[35][25] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26043_ (.D(_06920_),
    .Q(\design_top.MEM[35][26] ),
    .CLK(clknet_leaf_385_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26044_ (.D(_06921_),
    .Q(\design_top.MEM[35][27] ),
    .CLK(clknet_leaf_357_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26045_ (.D(_06922_),
    .Q(\design_top.MEM[35][28] ),
    .CLK(clknet_leaf_355_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26046_ (.D(_06923_),
    .Q(\design_top.MEM[35][29] ),
    .CLK(clknet_leaf_355_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26047_ (.D(_06924_),
    .Q(\design_top.MEM[35][30] ),
    .CLK(clknet_leaf_355_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26048_ (.D(_06925_),
    .Q(\design_top.MEM[35][31] ),
    .CLK(clknet_leaf_356_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26049_ (.D(_06926_),
    .Q(\design_top.MEM[20][8] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26050_ (.D(_06927_),
    .Q(\design_top.MEM[20][9] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26051_ (.D(_06928_),
    .Q(\design_top.MEM[20][10] ),
    .CLK(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26052_ (.D(_06929_),
    .Q(\design_top.MEM[20][11] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26053_ (.D(_06930_),
    .Q(\design_top.MEM[20][12] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26054_ (.D(_06931_),
    .Q(\design_top.MEM[20][13] ),
    .CLK(clknet_leaf_31_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26055_ (.D(_06932_),
    .Q(\design_top.MEM[20][14] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26056_ (.D(_06933_),
    .Q(\design_top.MEM[20][15] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26057_ (.D(_06934_),
    .Q(\design_top.MEM[35][16] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26058_ (.D(_06935_),
    .Q(\design_top.MEM[35][17] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26059_ (.D(_06936_),
    .Q(\design_top.MEM[35][18] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26060_ (.D(_06937_),
    .Q(\design_top.MEM[35][19] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26061_ (.D(_06938_),
    .Q(\design_top.MEM[35][20] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26062_ (.D(_06939_),
    .Q(\design_top.MEM[35][21] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26063_ (.D(_06940_),
    .Q(\design_top.MEM[35][22] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26064_ (.D(_06941_),
    .Q(\design_top.MEM[35][23] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26065_ (.D(_06942_),
    .Q(\design_top.MEM[45][16] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26066_ (.D(_06943_),
    .Q(\design_top.MEM[45][17] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26067_ (.D(_06944_),
    .Q(\design_top.MEM[45][18] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26068_ (.D(_06945_),
    .Q(\design_top.MEM[45][19] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26069_ (.D(_06946_),
    .Q(\design_top.MEM[45][20] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26070_ (.D(_06947_),
    .Q(\design_top.MEM[45][21] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26071_ (.D(_06948_),
    .Q(\design_top.MEM[45][22] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26072_ (.D(_06949_),
    .Q(\design_top.MEM[45][23] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26073_ (.D(_06950_),
    .Q(\design_top.MEM[35][8] ),
    .CLK(clknet_leaf_79_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26074_ (.D(_06951_),
    .Q(\design_top.MEM[35][9] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26075_ (.D(_06952_),
    .Q(\design_top.MEM[35][10] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26076_ (.D(_06953_),
    .Q(\design_top.MEM[35][11] ),
    .CLK(clknet_leaf_79_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26077_ (.D(_06954_),
    .Q(\design_top.MEM[35][12] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26078_ (.D(_06955_),
    .Q(\design_top.MEM[35][13] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26079_ (.D(_06956_),
    .Q(\design_top.MEM[35][14] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26080_ (.D(_06957_),
    .Q(\design_top.MEM[35][15] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26081_ (.D(_06958_),
    .Q(\design_top.MEM[34][16] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26082_ (.D(_06959_),
    .Q(\design_top.MEM[34][17] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26083_ (.D(_06960_),
    .Q(\design_top.MEM[34][18] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26084_ (.D(_06961_),
    .Q(\design_top.MEM[34][19] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26085_ (.D(_06962_),
    .Q(\design_top.MEM[34][20] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26086_ (.D(_06963_),
    .Q(\design_top.MEM[34][21] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26087_ (.D(_06964_),
    .Q(\design_top.MEM[34][22] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26088_ (.D(_06965_),
    .Q(\design_top.MEM[34][23] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26089_ (.D(_06966_),
    .Q(\design_top.MEM[34][8] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26090_ (.D(_06967_),
    .Q(\design_top.MEM[34][9] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26091_ (.D(_06968_),
    .Q(\design_top.MEM[34][10] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26092_ (.D(_06969_),
    .Q(\design_top.MEM[34][11] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26093_ (.D(_06970_),
    .Q(\design_top.MEM[34][12] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26094_ (.D(_06971_),
    .Q(\design_top.MEM[34][13] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26095_ (.D(_06972_),
    .Q(\design_top.MEM[34][14] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26096_ (.D(_06973_),
    .Q(\design_top.MEM[34][15] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26097_ (.D(_06974_),
    .Q(\design_top.MEM[19][24] ),
    .CLK(clknet_leaf_400_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26098_ (.D(_06975_),
    .Q(\design_top.MEM[19][25] ),
    .CLK(clknet_leaf_402_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26099_ (.D(_06976_),
    .Q(\design_top.MEM[19][26] ),
    .CLK(clknet_leaf_392_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26100_ (.D(_06977_),
    .Q(\design_top.MEM[19][27] ),
    .CLK(clknet_leaf_416_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26101_ (.D(_06978_),
    .Q(\design_top.MEM[19][28] ),
    .CLK(clknet_leaf_416_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26102_ (.D(_06979_),
    .Q(\design_top.MEM[19][29] ),
    .CLK(clknet_leaf_417_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26103_ (.D(_06980_),
    .Q(\design_top.MEM[19][30] ),
    .CLK(clknet_leaf_417_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26104_ (.D(_06981_),
    .Q(\design_top.MEM[19][31] ),
    .CLK(clknet_leaf_417_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26105_ (.D(_06982_),
    .Q(\design_top.MEM[19][16] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26106_ (.D(_06983_),
    .Q(\design_top.MEM[19][17] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26107_ (.D(_06984_),
    .Q(\design_top.MEM[19][18] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26108_ (.D(_06985_),
    .Q(\design_top.MEM[19][19] ),
    .CLK(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26109_ (.D(_06986_),
    .Q(\design_top.MEM[19][20] ),
    .CLK(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26110_ (.D(_06987_),
    .Q(\design_top.MEM[19][21] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26111_ (.D(_06988_),
    .Q(\design_top.MEM[19][22] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26112_ (.D(_06989_),
    .Q(\design_top.MEM[19][23] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26113_ (.D(_06990_),
    .Q(\design_top.MEM[19][8] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26114_ (.D(_06991_),
    .Q(\design_top.MEM[19][9] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26115_ (.D(_06992_),
    .Q(\design_top.MEM[19][10] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26116_ (.D(_06993_),
    .Q(\design_top.MEM[19][11] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26117_ (.D(_06994_),
    .Q(\design_top.MEM[19][12] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26118_ (.D(_06995_),
    .Q(\design_top.MEM[19][13] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26119_ (.D(_06996_),
    .Q(\design_top.MEM[19][14] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26120_ (.D(_06997_),
    .Q(\design_top.MEM[19][15] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26121_ (.D(_06998_),
    .Q(\design_top.MEM[18][24] ),
    .CLK(clknet_leaf_391_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26122_ (.D(_06999_),
    .Q(\design_top.MEM[18][25] ),
    .CLK(clknet_leaf_402_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26123_ (.D(_07000_),
    .Q(\design_top.MEM[18][26] ),
    .CLK(clknet_leaf_391_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26124_ (.D(_07001_),
    .Q(\design_top.MEM[18][27] ),
    .CLK(clknet_leaf_416_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26125_ (.D(_07002_),
    .Q(\design_top.MEM[18][28] ),
    .CLK(clknet_leaf_418_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26126_ (.D(_07003_),
    .Q(\design_top.MEM[18][29] ),
    .CLK(clknet_leaf_417_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26127_ (.D(_07004_),
    .Q(\design_top.MEM[18][30] ),
    .CLK(clknet_leaf_416_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26128_ (.D(_07005_),
    .Q(\design_top.MEM[18][31] ),
    .CLK(clknet_leaf_418_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26129_ (.D(_07006_),
    .Q(\design_top.MEM[18][16] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26130_ (.D(_07007_),
    .Q(\design_top.MEM[18][17] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26131_ (.D(_07008_),
    .Q(\design_top.MEM[18][18] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26132_ (.D(_07009_),
    .Q(\design_top.MEM[18][19] ),
    .CLK(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26133_ (.D(_07010_),
    .Q(\design_top.MEM[18][20] ),
    .CLK(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26134_ (.D(_07011_),
    .Q(\design_top.MEM[18][21] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26135_ (.D(_07012_),
    .Q(\design_top.MEM[18][22] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26136_ (.D(_07013_),
    .Q(\design_top.MEM[18][23] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26137_ (.D(_07014_),
    .Q(\design_top.MEM[18][8] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26138_ (.D(_07015_),
    .Q(\design_top.MEM[18][9] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26139_ (.D(_07016_),
    .Q(\design_top.MEM[18][10] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26140_ (.D(_07017_),
    .Q(\design_top.MEM[18][11] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26141_ (.D(_07018_),
    .Q(\design_top.MEM[18][12] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26142_ (.D(_07019_),
    .Q(\design_top.MEM[18][13] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26143_ (.D(_07020_),
    .Q(\design_top.MEM[18][14] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26144_ (.D(_07021_),
    .Q(\design_top.MEM[18][15] ),
    .CLK(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26145_ (.D(_07022_),
    .Q(\design_top.MEM[17][24] ),
    .CLK(clknet_leaf_399_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26146_ (.D(_07023_),
    .Q(\design_top.MEM[17][25] ),
    .CLK(clknet_leaf_397_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26147_ (.D(_07024_),
    .Q(\design_top.MEM[17][26] ),
    .CLK(clknet_leaf_392_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26148_ (.D(_07025_),
    .Q(\design_top.MEM[17][27] ),
    .CLK(clknet_leaf_415_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26149_ (.D(_07026_),
    .Q(\design_top.MEM[17][28] ),
    .CLK(clknet_leaf_414_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26150_ (.D(_07027_),
    .Q(\design_top.MEM[17][29] ),
    .CLK(clknet_leaf_417_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26151_ (.D(_07028_),
    .Q(\design_top.MEM[17][30] ),
    .CLK(clknet_leaf_417_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26152_ (.D(_07029_),
    .Q(\design_top.MEM[17][31] ),
    .CLK(clknet_leaf_418_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26153_ (.D(_07030_),
    .Q(\design_top.MEM[17][16] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26154_ (.D(_07031_),
    .Q(\design_top.MEM[17][17] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26155_ (.D(_07032_),
    .Q(\design_top.MEM[17][18] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26156_ (.D(_07033_),
    .Q(\design_top.MEM[17][19] ),
    .CLK(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26157_ (.D(_07034_),
    .Q(\design_top.MEM[17][20] ),
    .CLK(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26158_ (.D(_07035_),
    .Q(\design_top.MEM[17][21] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26159_ (.D(_07036_),
    .Q(\design_top.MEM[17][22] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26160_ (.D(_07037_),
    .Q(\design_top.MEM[17][23] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26161_ (.D(_07038_),
    .Q(\design_top.MEM[34][24] ),
    .CLK(clknet_leaf_390_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26162_ (.D(_07039_),
    .Q(\design_top.MEM[34][25] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26163_ (.D(_07040_),
    .Q(\design_top.MEM[34][26] ),
    .CLK(clknet_leaf_385_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26164_ (.D(_07041_),
    .Q(\design_top.MEM[34][27] ),
    .CLK(clknet_leaf_357_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26165_ (.D(_07042_),
    .Q(\design_top.MEM[34][28] ),
    .CLK(clknet_leaf_356_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26166_ (.D(_07043_),
    .Q(\design_top.MEM[34][29] ),
    .CLK(clknet_leaf_356_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26167_ (.D(_07044_),
    .Q(\design_top.MEM[34][30] ),
    .CLK(clknet_leaf_356_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26168_ (.D(_07045_),
    .Q(\design_top.MEM[34][31] ),
    .CLK(clknet_leaf_356_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26169_ (.D(_07046_),
    .Q(\design_top.MEM[33][24] ),
    .CLK(clknet_leaf_390_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26170_ (.D(_07047_),
    .Q(\design_top.MEM[33][25] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26171_ (.D(_07048_),
    .Q(\design_top.MEM[33][26] ),
    .CLK(clknet_leaf_385_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26172_ (.D(_07049_),
    .Q(\design_top.MEM[33][27] ),
    .CLK(clknet_leaf_356_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26173_ (.D(_07050_),
    .Q(\design_top.MEM[33][28] ),
    .CLK(clknet_leaf_356_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26174_ (.D(_07051_),
    .Q(\design_top.MEM[33][29] ),
    .CLK(clknet_leaf_355_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26175_ (.D(_07052_),
    .Q(\design_top.MEM[33][30] ),
    .CLK(clknet_leaf_355_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26176_ (.D(_07053_),
    .Q(\design_top.MEM[33][31] ),
    .CLK(clknet_leaf_356_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26177_ (.D(_07054_),
    .Q(\design_top.MEM[33][16] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26178_ (.D(_07055_),
    .Q(\design_top.MEM[33][17] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26179_ (.D(_07056_),
    .Q(\design_top.MEM[33][18] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26180_ (.D(_07057_),
    .Q(\design_top.MEM[33][19] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26181_ (.D(_07058_),
    .Q(\design_top.MEM[33][20] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26182_ (.D(_07059_),
    .Q(\design_top.MEM[33][21] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26183_ (.D(_07060_),
    .Q(\design_top.MEM[33][22] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26184_ (.D(_07061_),
    .Q(\design_top.MEM[33][23] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26185_ (.D(_07062_),
    .Q(\design_top.MEM[33][8] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26186_ (.D(_07063_),
    .Q(\design_top.MEM[33][9] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26187_ (.D(_07064_),
    .Q(\design_top.MEM[33][10] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26188_ (.D(_07065_),
    .Q(\design_top.MEM[33][11] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26189_ (.D(_07066_),
    .Q(\design_top.MEM[33][12] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26190_ (.D(_07067_),
    .Q(\design_top.MEM[33][13] ),
    .CLK(clknet_leaf_84_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26191_ (.D(_07068_),
    .Q(\design_top.MEM[33][14] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26192_ (.D(_07069_),
    .Q(\design_top.MEM[33][15] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26193_ (.D(_07070_),
    .Q(\design_top.MEM[32][24] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26194_ (.D(_07071_),
    .Q(\design_top.MEM[32][25] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26195_ (.D(_07072_),
    .Q(\design_top.MEM[32][26] ),
    .CLK(clknet_leaf_388_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26196_ (.D(_07073_),
    .Q(\design_top.MEM[32][27] ),
    .CLK(clknet_leaf_416_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26197_ (.D(_07074_),
    .Q(\design_top.MEM[32][28] ),
    .CLK(clknet_leaf_416_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26198_ (.D(_07075_),
    .Q(\design_top.MEM[32][29] ),
    .CLK(clknet_leaf_356_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26199_ (.D(_07076_),
    .Q(\design_top.MEM[32][30] ),
    .CLK(clknet_leaf_417_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26200_ (.D(_07077_),
    .Q(\design_top.MEM[32][31] ),
    .CLK(clknet_leaf_417_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26201_ (.D(_07078_),
    .Q(\design_top.MEM[17][8] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26202_ (.D(_07079_),
    .Q(\design_top.MEM[17][9] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26203_ (.D(_07080_),
    .Q(\design_top.MEM[17][10] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26204_ (.D(_07081_),
    .Q(\design_top.MEM[17][11] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26205_ (.D(_07082_),
    .Q(\design_top.MEM[17][12] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26206_ (.D(_07083_),
    .Q(\design_top.MEM[17][13] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26207_ (.D(_07084_),
    .Q(\design_top.MEM[17][14] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26208_ (.D(_07085_),
    .Q(\design_top.MEM[17][15] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26209_ (.D(_07086_),
    .Q(\design_top.MEM[16][24] ),
    .CLK(clknet_leaf_391_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26210_ (.D(_07087_),
    .Q(\design_top.MEM[16][25] ),
    .CLK(clknet_leaf_402_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26211_ (.D(_07088_),
    .Q(\design_top.MEM[16][26] ),
    .CLK(clknet_leaf_389_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26212_ (.D(_07089_),
    .Q(\design_top.MEM[16][27] ),
    .CLK(clknet_leaf_416_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26213_ (.D(_07090_),
    .Q(\design_top.MEM[16][28] ),
    .CLK(clknet_leaf_416_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26214_ (.D(_07091_),
    .Q(\design_top.MEM[16][29] ),
    .CLK(clknet_leaf_417_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26215_ (.D(_07092_),
    .Q(\design_top.MEM[16][30] ),
    .CLK(clknet_leaf_416_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26216_ (.D(_07093_),
    .Q(\design_top.MEM[16][31] ),
    .CLK(clknet_leaf_418_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26217_ (.D(_07094_),
    .Q(\design_top.MEM[16][16] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26218_ (.D(_07095_),
    .Q(\design_top.MEM[16][17] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26219_ (.D(_07096_),
    .Q(\design_top.MEM[16][18] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26220_ (.D(_07097_),
    .Q(\design_top.MEM[16][19] ),
    .CLK(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26221_ (.D(_07098_),
    .Q(\design_top.MEM[16][20] ),
    .CLK(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26222_ (.D(_07099_),
    .Q(\design_top.MEM[16][21] ),
    .CLK(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26223_ (.D(_07100_),
    .Q(\design_top.MEM[16][22] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26224_ (.D(_07101_),
    .Q(\design_top.MEM[16][23] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26225_ (.D(_07102_),
    .Q(\design_top.MEM[16][8] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26226_ (.D(_07103_),
    .Q(\design_top.MEM[16][9] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26227_ (.D(_07104_),
    .Q(\design_top.MEM[16][10] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26228_ (.D(_07105_),
    .Q(\design_top.MEM[16][11] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26229_ (.D(_07106_),
    .Q(\design_top.MEM[16][12] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26230_ (.D(_07107_),
    .Q(\design_top.MEM[16][13] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26231_ (.D(_07108_),
    .Q(\design_top.MEM[16][14] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26232_ (.D(_07109_),
    .Q(\design_top.MEM[16][15] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26233_ (.D(_07110_),
    .Q(\design_top.MEM[15][24] ),
    .CLK(clknet_leaf_390_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26234_ (.D(_07111_),
    .Q(\design_top.MEM[15][25] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26235_ (.D(_07112_),
    .Q(\design_top.MEM[15][26] ),
    .CLK(clknet_leaf_390_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26236_ (.D(_07113_),
    .Q(\design_top.MEM[15][27] ),
    .CLK(clknet_leaf_409_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26237_ (.D(_07114_),
    .Q(\design_top.MEM[15][28] ),
    .CLK(clknet_leaf_409_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26238_ (.D(_07115_),
    .Q(\design_top.MEM[15][29] ),
    .CLK(clknet_leaf_396_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26239_ (.D(_07116_),
    .Q(\design_top.MEM[15][30] ),
    .CLK(clknet_leaf_394_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26240_ (.D(_07117_),
    .Q(\design_top.MEM[15][31] ),
    .CLK(clknet_leaf_394_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26241_ (.D(_07118_),
    .Q(\design_top.MEM[15][16] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26242_ (.D(_07119_),
    .Q(\design_top.MEM[15][17] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26243_ (.D(_07120_),
    .Q(\design_top.MEM[15][18] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26244_ (.D(_07121_),
    .Q(\design_top.MEM[15][19] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26245_ (.D(_07122_),
    .Q(\design_top.MEM[15][20] ),
    .CLK(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26246_ (.D(_07123_),
    .Q(\design_top.MEM[15][21] ),
    .CLK(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26247_ (.D(_07124_),
    .Q(\design_top.MEM[15][22] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26248_ (.D(_07125_),
    .Q(\design_top.MEM[15][23] ),
    .CLK(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26249_ (.D(_07126_),
    .Q(\design_top.MEM[15][8] ),
    .CLK(clknet_leaf_79_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26250_ (.D(_07127_),
    .Q(\design_top.MEM[15][9] ),
    .CLK(clknet_leaf_79_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26251_ (.D(_07128_),
    .Q(\design_top.MEM[15][10] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26252_ (.D(_07129_),
    .Q(\design_top.MEM[15][11] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26253_ (.D(_07130_),
    .Q(\design_top.MEM[15][12] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26254_ (.D(_07131_),
    .Q(\design_top.MEM[15][13] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26255_ (.D(_07132_),
    .Q(\design_top.MEM[15][14] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26256_ (.D(_07133_),
    .Q(\design_top.MEM[15][15] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26257_ (.D(_07134_),
    .Q(\design_top.MEM[14][24] ),
    .CLK(clknet_leaf_390_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26258_ (.D(_07135_),
    .Q(\design_top.MEM[14][25] ),
    .CLK(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26259_ (.D(_07136_),
    .Q(\design_top.MEM[14][26] ),
    .CLK(clknet_leaf_390_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26260_ (.D(_07137_),
    .Q(\design_top.MEM[14][27] ),
    .CLK(clknet_leaf_396_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26261_ (.D(_07138_),
    .Q(\design_top.MEM[14][28] ),
    .CLK(clknet_leaf_395_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26262_ (.D(_07139_),
    .Q(\design_top.MEM[14][29] ),
    .CLK(clknet_leaf_396_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26263_ (.D(_07140_),
    .Q(\design_top.MEM[14][30] ),
    .CLK(clknet_leaf_396_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26264_ (.D(_07141_),
    .Q(\design_top.MEM[14][31] ),
    .CLK(clknet_leaf_394_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26265_ (.D(_07142_),
    .Q(\design_top.MEM[14][16] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26266_ (.D(_07143_),
    .Q(\design_top.MEM[14][17] ),
    .CLK(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26267_ (.D(_07144_),
    .Q(\design_top.MEM[14][18] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26268_ (.D(_07145_),
    .Q(\design_top.MEM[14][19] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26269_ (.D(_07146_),
    .Q(\design_top.MEM[14][20] ),
    .CLK(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26270_ (.D(_07147_),
    .Q(\design_top.MEM[14][21] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26271_ (.D(_07148_),
    .Q(\design_top.MEM[14][22] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26272_ (.D(_07149_),
    .Q(\design_top.MEM[14][23] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26273_ (.D(_07150_),
    .Q(\design_top.MEM[14][8] ),
    .CLK(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26274_ (.D(_07151_),
    .Q(\design_top.MEM[14][9] ),
    .CLK(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26275_ (.D(_07152_),
    .Q(\design_top.MEM[14][10] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26276_ (.D(_07153_),
    .Q(\design_top.MEM[14][11] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26277_ (.D(_07154_),
    .Q(\design_top.MEM[14][12] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26278_ (.D(_07155_),
    .Q(\design_top.MEM[14][13] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26279_ (.D(_07156_),
    .Q(\design_top.MEM[14][14] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26280_ (.D(_07157_),
    .Q(\design_top.MEM[14][15] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26281_ (.D(_07158_),
    .Q(\design_top.MEM[13][24] ),
    .CLK(clknet_leaf_390_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26282_ (.D(_07159_),
    .Q(\design_top.MEM[13][25] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26283_ (.D(_07160_),
    .Q(\design_top.MEM[13][26] ),
    .CLK(clknet_leaf_390_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26284_ (.D(_07161_),
    .Q(\design_top.MEM[13][27] ),
    .CLK(clknet_leaf_396_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26285_ (.D(_07162_),
    .Q(\design_top.MEM[13][28] ),
    .CLK(clknet_leaf_395_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26286_ (.D(_07163_),
    .Q(\design_top.MEM[13][29] ),
    .CLK(clknet_leaf_396_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26287_ (.D(_07164_),
    .Q(\design_top.MEM[13][30] ),
    .CLK(clknet_leaf_396_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26288_ (.D(_07165_),
    .Q(\design_top.MEM[13][31] ),
    .CLK(clknet_leaf_392_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26289_ (.D(_07166_),
    .Q(\design_top.MEM[13][16] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26290_ (.D(_07167_),
    .Q(\design_top.MEM[13][17] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26291_ (.D(_07168_),
    .Q(\design_top.MEM[13][18] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26292_ (.D(_07169_),
    .Q(\design_top.MEM[13][19] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26293_ (.D(_07170_),
    .Q(\design_top.MEM[13][20] ),
    .CLK(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26294_ (.D(_07171_),
    .Q(\design_top.MEM[13][21] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26295_ (.D(_07172_),
    .Q(\design_top.MEM[13][22] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26296_ (.D(_07173_),
    .Q(\design_top.MEM[13][23] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26297_ (.D(_07174_),
    .Q(\design_top.MEM[13][8] ),
    .CLK(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26298_ (.D(_07175_),
    .Q(\design_top.MEM[13][9] ),
    .CLK(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26299_ (.D(_07176_),
    .Q(\design_top.MEM[13][10] ),
    .CLK(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26300_ (.D(_07177_),
    .Q(\design_top.MEM[13][11] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26301_ (.D(_07178_),
    .Q(\design_top.MEM[13][12] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26302_ (.D(_07179_),
    .Q(\design_top.MEM[13][13] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26303_ (.D(_07180_),
    .Q(\design_top.MEM[13][14] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26304_ (.D(_07181_),
    .Q(\design_top.MEM[13][15] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26305_ (.D(_07182_),
    .Q(\design_top.MEM[12][24] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26306_ (.D(_07183_),
    .Q(\design_top.MEM[12][25] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26307_ (.D(_07184_),
    .Q(\design_top.MEM[12][26] ),
    .CLK(clknet_leaf_390_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26308_ (.D(_07185_),
    .Q(\design_top.MEM[12][27] ),
    .CLK(clknet_leaf_408_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26309_ (.D(_07186_),
    .Q(\design_top.MEM[12][28] ),
    .CLK(clknet_leaf_397_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26310_ (.D(_07187_),
    .Q(\design_top.MEM[12][29] ),
    .CLK(clknet_leaf_396_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26311_ (.D(_07188_),
    .Q(\design_top.MEM[12][30] ),
    .CLK(clknet_leaf_396_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26312_ (.D(_07189_),
    .Q(\design_top.MEM[12][31] ),
    .CLK(clknet_leaf_399_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26313_ (.D(_07190_),
    .Q(\design_top.MEM[12][16] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26314_ (.D(_07191_),
    .Q(\design_top.MEM[12][17] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26315_ (.D(_07192_),
    .Q(\design_top.MEM[12][18] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26316_ (.D(_07193_),
    .Q(\design_top.MEM[12][19] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26317_ (.D(_07194_),
    .Q(\design_top.MEM[12][20] ),
    .CLK(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26318_ (.D(_07195_),
    .Q(\design_top.MEM[12][21] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26319_ (.D(_07196_),
    .Q(\design_top.MEM[12][22] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26320_ (.D(_07197_),
    .Q(\design_top.MEM[12][23] ),
    .CLK(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26321_ (.D(_07198_),
    .Q(\design_top.MEM[12][8] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26322_ (.D(_07199_),
    .Q(\design_top.MEM[12][9] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26323_ (.D(_07200_),
    .Q(\design_top.MEM[12][10] ),
    .CLK(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26324_ (.D(_07201_),
    .Q(\design_top.MEM[12][11] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26325_ (.D(_07202_),
    .Q(\design_top.MEM[12][12] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26326_ (.D(_07203_),
    .Q(\design_top.MEM[12][13] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26327_ (.D(_07204_),
    .Q(\design_top.MEM[12][14] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26328_ (.D(_07205_),
    .Q(\design_top.MEM[12][15] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26329_ (.D(_07206_),
    .Q(\design_top.MEM[11][24] ),
    .CLK(clknet_leaf_390_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26330_ (.D(_07207_),
    .Q(\design_top.MEM[11][25] ),
    .CLK(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26331_ (.D(_07208_),
    .Q(\design_top.MEM[11][26] ),
    .CLK(clknet_leaf_388_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26332_ (.D(_07209_),
    .Q(\design_top.MEM[11][27] ),
    .CLK(clknet_leaf_379_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26333_ (.D(_07210_),
    .Q(\design_top.MEM[11][28] ),
    .CLK(clknet_leaf_395_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26334_ (.D(_07211_),
    .Q(\design_top.MEM[11][29] ),
    .CLK(clknet_leaf_379_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26335_ (.D(_07212_),
    .Q(\design_top.MEM[11][30] ),
    .CLK(clknet_leaf_379_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26336_ (.D(_07213_),
    .Q(\design_top.MEM[11][31] ),
    .CLK(clknet_leaf_394_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26337_ (.D(_07214_),
    .Q(\design_top.MEM[11][16] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26338_ (.D(_07215_),
    .Q(\design_top.MEM[11][17] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26339_ (.D(_07216_),
    .Q(\design_top.MEM[11][18] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26340_ (.D(_07217_),
    .Q(\design_top.MEM[11][19] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26341_ (.D(_07218_),
    .Q(\design_top.MEM[11][20] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26342_ (.D(_07219_),
    .Q(\design_top.MEM[11][21] ),
    .CLK(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26343_ (.D(_07220_),
    .Q(\design_top.MEM[11][22] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26344_ (.D(_07221_),
    .Q(\design_top.MEM[11][23] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26345_ (.D(_07222_),
    .Q(\design_top.MEM[11][8] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26346_ (.D(_07223_),
    .Q(\design_top.MEM[11][9] ),
    .CLK(clknet_leaf_76_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26347_ (.D(_07224_),
    .Q(\design_top.MEM[11][10] ),
    .CLK(clknet_leaf_76_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26348_ (.D(_07225_),
    .Q(\design_top.MEM[11][11] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26349_ (.D(_07226_),
    .Q(\design_top.MEM[11][12] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26350_ (.D(_07227_),
    .Q(\design_top.MEM[11][13] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26351_ (.D(_07228_),
    .Q(\design_top.MEM[11][14] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26352_ (.D(_07229_),
    .Q(\design_top.MEM[11][15] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26353_ (.D(_07230_),
    .Q(\design_top.MEM[10][24] ),
    .CLK(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26354_ (.D(_07231_),
    .Q(\design_top.MEM[10][25] ),
    .CLK(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26355_ (.D(_07232_),
    .Q(\design_top.MEM[10][26] ),
    .CLK(clknet_leaf_388_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26356_ (.D(_07233_),
    .Q(\design_top.MEM[10][27] ),
    .CLK(clknet_leaf_395_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26357_ (.D(_07234_),
    .Q(\design_top.MEM[10][28] ),
    .CLK(clknet_leaf_395_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26358_ (.D(_07235_),
    .Q(\design_top.MEM[10][29] ),
    .CLK(clknet_leaf_395_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26359_ (.D(_07236_),
    .Q(\design_top.MEM[10][30] ),
    .CLK(clknet_leaf_394_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26360_ (.D(_07237_),
    .Q(\design_top.MEM[10][31] ),
    .CLK(clknet_leaf_394_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26361_ (.D(_07238_),
    .Q(\design_top.MEM[10][16] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26362_ (.D(_07239_),
    .Q(\design_top.MEM[10][17] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26363_ (.D(_07240_),
    .Q(\design_top.MEM[10][18] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26364_ (.D(_07241_),
    .Q(\design_top.MEM[10][19] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26365_ (.D(_07242_),
    .Q(\design_top.MEM[10][20] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26366_ (.D(_07243_),
    .Q(\design_top.MEM[10][21] ),
    .CLK(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26367_ (.D(_07244_),
    .Q(\design_top.MEM[10][22] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26368_ (.D(_07245_),
    .Q(\design_top.MEM[10][23] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26369_ (.D(_07246_),
    .Q(\design_top.MEM[10][8] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26370_ (.D(_07247_),
    .Q(\design_top.MEM[10][9] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26371_ (.D(_07248_),
    .Q(\design_top.MEM[10][10] ),
    .CLK(clknet_leaf_76_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26372_ (.D(_07249_),
    .Q(\design_top.MEM[10][11] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26373_ (.D(_07250_),
    .Q(\design_top.MEM[10][12] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26374_ (.D(_07251_),
    .Q(\design_top.MEM[10][13] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26375_ (.D(_07252_),
    .Q(\design_top.MEM[10][14] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26376_ (.D(_07253_),
    .Q(\design_top.MEM[10][15] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26377_ (.D(_07254_),
    .Q(\design_top.MEM[0][24] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26378_ (.D(_07255_),
    .Q(\design_top.MEM[0][25] ),
    .CLK(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26379_ (.D(_07256_),
    .Q(\design_top.MEM[0][26] ),
    .CLK(clknet_leaf_388_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26380_ (.D(_07257_),
    .Q(\design_top.MEM[0][27] ),
    .CLK(clknet_leaf_364_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26381_ (.D(_07258_),
    .Q(\design_top.MEM[0][28] ),
    .CLK(clknet_leaf_409_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26382_ (.D(_07259_),
    .Q(\design_top.MEM[0][29] ),
    .CLK(clknet_leaf_363_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26383_ (.D(_07260_),
    .Q(\design_top.MEM[0][30] ),
    .CLK(clknet_leaf_364_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26384_ (.D(_07261_),
    .Q(\design_top.MEM[0][31] ),
    .CLK(clknet_leaf_409_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26385_ (.D(_07262_),
    .Q(\design_top.MEM[0][16] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26386_ (.D(_07263_),
    .Q(\design_top.MEM[0][17] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26387_ (.D(_07264_),
    .Q(\design_top.MEM[0][18] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26388_ (.D(_07265_),
    .Q(\design_top.MEM[0][19] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26389_ (.D(_07266_),
    .Q(\design_top.MEM[0][20] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26390_ (.D(_07267_),
    .Q(\design_top.MEM[0][21] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26391_ (.D(_07268_),
    .Q(\design_top.MEM[0][22] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26392_ (.D(_07269_),
    .Q(\design_top.MEM[0][23] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26393_ (.D(_07270_),
    .Q(\design_top.MEM[32][16] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26394_ (.D(_07271_),
    .Q(\design_top.MEM[32][17] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26395_ (.D(_07272_),
    .Q(\design_top.MEM[32][18] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26396_ (.D(_07273_),
    .Q(\design_top.MEM[32][19] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26397_ (.D(_07274_),
    .Q(\design_top.MEM[32][20] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26398_ (.D(_07275_),
    .Q(\design_top.MEM[32][21] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26399_ (.D(_07276_),
    .Q(\design_top.MEM[32][22] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26400_ (.D(_07277_),
    .Q(\design_top.MEM[32][23] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26401_ (.D(_07278_),
    .Q(\design_top.MEM[32][8] ),
    .CLK(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26402_ (.D(_07279_),
    .Q(\design_top.MEM[32][9] ),
    .CLK(clknet_leaf_79_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26403_ (.D(_07280_),
    .Q(\design_top.MEM[32][10] ),
    .CLK(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26404_ (.D(_07281_),
    .Q(\design_top.MEM[32][11] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26405_ (.D(_07282_),
    .Q(\design_top.MEM[32][12] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26406_ (.D(_07283_),
    .Q(\design_top.MEM[32][13] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26407_ (.D(_07284_),
    .Q(\design_top.MEM[32][14] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26408_ (.D(_07285_),
    .Q(\design_top.MEM[32][15] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26409_ (.D(_07286_),
    .Q(\design_top.MEM[31][24] ),
    .CLK(clknet_leaf_397_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26410_ (.D(_07287_),
    .Q(\design_top.MEM[31][25] ),
    .CLK(clknet_leaf_400_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26411_ (.D(_07288_),
    .Q(\design_top.MEM[31][26] ),
    .CLK(clknet_leaf_390_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26412_ (.D(_07289_),
    .Q(\design_top.MEM[31][27] ),
    .CLK(clknet_leaf_407_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26413_ (.D(_07290_),
    .Q(\design_top.MEM[31][28] ),
    .CLK(clknet_leaf_407_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26414_ (.D(_07291_),
    .Q(\design_top.MEM[31][29] ),
    .CLK(clknet_leaf_407_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26415_ (.D(_07292_),
    .Q(\design_top.MEM[31][30] ),
    .CLK(clknet_leaf_407_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26416_ (.D(_07293_),
    .Q(\design_top.MEM[31][31] ),
    .CLK(clknet_leaf_408_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26417_ (.D(_07294_),
    .Q(\design_top.MEM[31][16] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26418_ (.D(_07295_),
    .Q(\design_top.MEM[31][17] ),
    .CLK(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26419_ (.D(_07296_),
    .Q(\design_top.MEM[31][18] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26420_ (.D(_07297_),
    .Q(\design_top.MEM[31][19] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26421_ (.D(_07298_),
    .Q(\design_top.MEM[31][20] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26422_ (.D(_07299_),
    .Q(\design_top.MEM[31][21] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26423_ (.D(_07300_),
    .Q(\design_top.MEM[31][22] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26424_ (.D(_07301_),
    .Q(\design_top.MEM[31][23] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26425_ (.D(_07302_),
    .Q(\design_top.MEM[31][8] ),
    .CLK(clknet_leaf_79_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26426_ (.D(_07303_),
    .Q(\design_top.MEM[31][9] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26427_ (.D(_07304_),
    .Q(\design_top.MEM[31][10] ),
    .CLK(clknet_leaf_79_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26428_ (.D(_07305_),
    .Q(\design_top.MEM[31][11] ),
    .CLK(clknet_leaf_79_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26429_ (.D(_07306_),
    .Q(\design_top.MEM[31][12] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26430_ (.D(_07307_),
    .Q(\design_top.MEM[31][13] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26431_ (.D(_07308_),
    .Q(\design_top.MEM[31][14] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26432_ (.D(_07309_),
    .Q(\design_top.MEM[31][15] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26433_ (.D(_07310_),
    .Q(\design_top.MEM[30][24] ),
    .CLK(clknet_leaf_397_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26434_ (.D(_07311_),
    .Q(\design_top.MEM[30][25] ),
    .CLK(clknet_leaf_400_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26435_ (.D(_07312_),
    .Q(\design_top.MEM[30][26] ),
    .CLK(clknet_leaf_391_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26436_ (.D(_07313_),
    .Q(\design_top.MEM[30][27] ),
    .CLK(clknet_leaf_406_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26437_ (.D(_07314_),
    .Q(\design_top.MEM[30][28] ),
    .CLK(clknet_leaf_413_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26438_ (.D(_07315_),
    .Q(\design_top.MEM[30][29] ),
    .CLK(clknet_leaf_412_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26439_ (.D(_07316_),
    .Q(\design_top.MEM[30][30] ),
    .CLK(clknet_leaf_412_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26440_ (.D(_07317_),
    .Q(\design_top.MEM[30][31] ),
    .CLK(clknet_leaf_408_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26441_ (.D(_07318_),
    .Q(\design_top.MEM[30][16] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26442_ (.D(_07319_),
    .Q(\design_top.MEM[30][17] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26443_ (.D(_07320_),
    .Q(\design_top.MEM[30][18] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26444_ (.D(_07321_),
    .Q(\design_top.MEM[30][19] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26445_ (.D(_07322_),
    .Q(\design_top.MEM[30][20] ),
    .CLK(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26446_ (.D(_07323_),
    .Q(\design_top.MEM[30][21] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26447_ (.D(_07324_),
    .Q(\design_top.MEM[30][22] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26448_ (.D(_07325_),
    .Q(\design_top.MEM[30][23] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26449_ (.D(_07326_),
    .Q(\design_top.MEM[30][8] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26450_ (.D(_07327_),
    .Q(\design_top.MEM[30][9] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26451_ (.D(_07328_),
    .Q(\design_top.MEM[30][10] ),
    .CLK(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26452_ (.D(_07329_),
    .Q(\design_top.MEM[30][11] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26453_ (.D(_07330_),
    .Q(\design_top.MEM[30][12] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26454_ (.D(_07331_),
    .Q(\design_top.MEM[30][13] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26455_ (.D(_07332_),
    .Q(\design_top.MEM[30][14] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26456_ (.D(_07333_),
    .Q(\design_top.MEM[30][15] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26457_ (.D(_07334_),
    .Q(\design_top.MEM[2][24] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26458_ (.D(_07335_),
    .Q(\design_top.MEM[2][25] ),
    .CLK(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26459_ (.D(_07336_),
    .Q(\design_top.MEM[2][26] ),
    .CLK(clknet_leaf_388_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26460_ (.D(_07337_),
    .Q(\design_top.MEM[2][27] ),
    .CLK(clknet_leaf_409_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26461_ (.D(_07338_),
    .Q(\design_top.MEM[2][28] ),
    .CLK(clknet_leaf_409_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26462_ (.D(_07339_),
    .Q(\design_top.MEM[2][29] ),
    .CLK(clknet_leaf_409_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26463_ (.D(_07340_),
    .Q(\design_top.MEM[2][30] ),
    .CLK(clknet_leaf_409_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26464_ (.D(_07341_),
    .Q(\design_top.MEM[2][31] ),
    .CLK(clknet_leaf_409_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26465_ (.D(_07342_),
    .Q(\design_top.MEM[2][16] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26466_ (.D(_07343_),
    .Q(\design_top.MEM[2][17] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26467_ (.D(_07344_),
    .Q(\design_top.MEM[2][18] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26468_ (.D(_07345_),
    .Q(\design_top.MEM[2][19] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26469_ (.D(_07346_),
    .Q(\design_top.MEM[2][20] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26470_ (.D(_07347_),
    .Q(\design_top.MEM[2][21] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26471_ (.D(_07348_),
    .Q(\design_top.MEM[2][22] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26472_ (.D(_07349_),
    .Q(\design_top.MEM[2][23] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26473_ (.D(_07350_),
    .Q(\design_top.MEM[2][8] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26474_ (.D(_07351_),
    .Q(\design_top.MEM[2][9] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26475_ (.D(_07352_),
    .Q(\design_top.MEM[2][10] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26476_ (.D(_07353_),
    .Q(\design_top.MEM[2][11] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26477_ (.D(_07354_),
    .Q(\design_top.MEM[2][12] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26478_ (.D(_07355_),
    .Q(\design_top.MEM[2][13] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26479_ (.D(_07356_),
    .Q(\design_top.MEM[2][14] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26480_ (.D(_07357_),
    .Q(\design_top.MEM[2][15] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26481_ (.D(_07358_),
    .Q(\design_top.MEM[29][24] ),
    .CLK(clknet_leaf_397_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26482_ (.D(_07359_),
    .Q(\design_top.MEM[29][25] ),
    .CLK(clknet_leaf_400_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26483_ (.D(_07360_),
    .Q(\design_top.MEM[29][26] ),
    .CLK(clknet_leaf_391_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26484_ (.D(_07361_),
    .Q(\design_top.MEM[29][27] ),
    .CLK(clknet_leaf_407_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26485_ (.D(_07362_),
    .Q(\design_top.MEM[29][28] ),
    .CLK(clknet_leaf_413_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26486_ (.D(_07363_),
    .Q(\design_top.MEM[29][29] ),
    .CLK(clknet_leaf_413_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26487_ (.D(_07364_),
    .Q(\design_top.MEM[29][30] ),
    .CLK(clknet_leaf_412_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26488_ (.D(_07365_),
    .Q(\design_top.MEM[29][31] ),
    .CLK(clknet_leaf_408_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26489_ (.D(_07366_),
    .Q(\design_top.MEM[29][16] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26490_ (.D(_07367_),
    .Q(\design_top.MEM[29][17] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26491_ (.D(_07368_),
    .Q(\design_top.MEM[29][18] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26492_ (.D(_07369_),
    .Q(\design_top.MEM[29][19] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26493_ (.D(_07370_),
    .Q(\design_top.MEM[29][20] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26494_ (.D(_07371_),
    .Q(\design_top.MEM[29][21] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26495_ (.D(_07372_),
    .Q(\design_top.MEM[29][22] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26496_ (.D(_07373_),
    .Q(\design_top.MEM[29][23] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26497_ (.D(_07374_),
    .Q(\design_top.MEM[29][8] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26498_ (.D(_07375_),
    .Q(\design_top.MEM[29][9] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26499_ (.D(_07376_),
    .Q(\design_top.MEM[29][10] ),
    .CLK(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26500_ (.D(_07377_),
    .Q(\design_top.MEM[29][11] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26501_ (.D(_07378_),
    .Q(\design_top.MEM[29][12] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26502_ (.D(_07379_),
    .Q(\design_top.MEM[29][13] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26503_ (.D(_07380_),
    .Q(\design_top.MEM[29][14] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26504_ (.D(_07381_),
    .Q(\design_top.MEM[29][15] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26505_ (.D(_07382_),
    .Q(\design_top.MEM[28][24] ),
    .CLK(clknet_leaf_397_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26506_ (.D(_07383_),
    .Q(\design_top.MEM[28][25] ),
    .CLK(clknet_leaf_400_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26507_ (.D(_07384_),
    .Q(\design_top.MEM[28][26] ),
    .CLK(clknet_leaf_391_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26508_ (.D(_07385_),
    .Q(\design_top.MEM[28][27] ),
    .CLK(clknet_leaf_412_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26509_ (.D(_07386_),
    .Q(\design_top.MEM[28][28] ),
    .CLK(clknet_leaf_413_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26510_ (.D(_07387_),
    .Q(\design_top.MEM[28][29] ),
    .CLK(clknet_leaf_412_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26511_ (.D(_07388_),
    .Q(\design_top.MEM[28][30] ),
    .CLK(clknet_leaf_412_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26512_ (.D(_07389_),
    .Q(\design_top.MEM[28][31] ),
    .CLK(clknet_leaf_407_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26513_ (.D(_07390_),
    .Q(\design_top.MEM[28][16] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26514_ (.D(_07391_),
    .Q(\design_top.MEM[28][17] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26515_ (.D(_07392_),
    .Q(\design_top.MEM[28][18] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26516_ (.D(_07393_),
    .Q(\design_top.MEM[28][19] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26517_ (.D(_07394_),
    .Q(\design_top.MEM[28][20] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26518_ (.D(_07395_),
    .Q(\design_top.MEM[28][21] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26519_ (.D(_07396_),
    .Q(\design_top.MEM[28][22] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26520_ (.D(_07397_),
    .Q(\design_top.MEM[28][23] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26521_ (.D(_07398_),
    .Q(\design_top.MEM[28][8] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26522_ (.D(_07399_),
    .Q(\design_top.MEM[28][9] ),
    .CLK(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26523_ (.D(_07400_),
    .Q(\design_top.MEM[28][10] ),
    .CLK(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26524_ (.D(_07401_),
    .Q(\design_top.MEM[28][11] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26525_ (.D(_07402_),
    .Q(\design_top.MEM[28][12] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26526_ (.D(_07403_),
    .Q(\design_top.MEM[28][13] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26527_ (.D(_07404_),
    .Q(\design_top.MEM[28][14] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26528_ (.D(_07405_),
    .Q(\design_top.MEM[28][15] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26529_ (.D(_07406_),
    .Q(\design_top.MEM[27][24] ),
    .CLK(clknet_leaf_396_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26530_ (.D(_07407_),
    .Q(\design_top.MEM[27][25] ),
    .CLK(clknet_leaf_399_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26531_ (.D(_07408_),
    .Q(\design_top.MEM[27][26] ),
    .CLK(clknet_leaf_392_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26532_ (.D(_07409_),
    .Q(\design_top.MEM[27][27] ),
    .CLK(clknet_leaf_411_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26533_ (.D(_07410_),
    .Q(\design_top.MEM[27][28] ),
    .CLK(clknet_leaf_413_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26534_ (.D(_07411_),
    .Q(\design_top.MEM[27][29] ),
    .CLK(clknet_leaf_414_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26535_ (.D(_07412_),
    .Q(\design_top.MEM[27][30] ),
    .CLK(clknet_leaf_411_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26536_ (.D(_07413_),
    .Q(\design_top.MEM[27][31] ),
    .CLK(clknet_leaf_409_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26537_ (.D(_07414_),
    .Q(\design_top.MEM[27][16] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26538_ (.D(_07415_),
    .Q(\design_top.MEM[27][17] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26539_ (.D(_07416_),
    .Q(\design_top.MEM[27][18] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26540_ (.D(_07417_),
    .Q(\design_top.MEM[27][19] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26541_ (.D(_07418_),
    .Q(\design_top.MEM[27][20] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26542_ (.D(_07419_),
    .Q(\design_top.MEM[27][21] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26543_ (.D(_07420_),
    .Q(\design_top.MEM[27][22] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26544_ (.D(_07421_),
    .Q(\design_top.MEM[27][23] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26545_ (.D(_07422_),
    .Q(\design_top.IREQ[7] ),
    .CLK(clknet_leaf_371_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26546_ (.D(_07423_),
    .Q(\design_top.IACK[7] ),
    .CLK(clknet_leaf_369_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26547_ (.D(_07424_),
    .Q(\design_top.MEM[0][8] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26548_ (.D(_07425_),
    .Q(\design_top.MEM[0][9] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26549_ (.D(_07426_),
    .Q(\design_top.MEM[0][10] ),
    .CLK(clknet_leaf_76_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26550_ (.D(_07427_),
    .Q(\design_top.MEM[0][11] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26551_ (.D(_07428_),
    .Q(\design_top.MEM[0][12] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26552_ (.D(_07429_),
    .Q(\design_top.MEM[0][13] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26553_ (.D(_07430_),
    .Q(\design_top.MEM[0][14] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _26554_ (.D(_07431_),
    .Q(\design_top.MEM[0][15] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_29_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_31_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_37_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_39_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_48_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_user_clock2 (.A(clknet_opt_6_user_clock2),
    .X(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_user_clock2 (.A(clknet_opt_11_user_clock2),
    .X(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_76_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_79_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_84_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_user_clock2 (.A(clknet_opt_1_user_clock2),
    .X(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_user_clock2 (.A(clknet_opt_10_user_clock2),
    .X(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_user_clock2 (.A(clknet_opt_16_user_clock2),
    .X(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_120_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_143_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_155_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_user_clock2 (.A(clknet_opt_15_user_clock2),
    .X(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_172_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_user_clock2 (.A(clknet_opt_12_user_clock2),
    .X(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_user_clock2 (.A(clknet_opt_13_user_clock2),
    .X(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_187_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_193_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_194_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_195_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_196_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_197_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_198_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_199_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_200_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_201_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_202_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_203_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_204_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_205_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_206_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_207_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_208_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_209_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_210_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_211_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_212_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_213_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_214_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_215_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_216_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_217_user_clock2 (.A(clknet_opt_21_user_clock2),
    .X(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_218_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_219_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_220_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_221_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_222_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_223_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_224_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_225_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_226_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_227_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_228_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_229_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_230_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_231_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_232_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_233_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_234_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_235_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_235_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_236_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_237_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_238_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_239_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_240_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_241_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_242_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_243_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_244_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_244_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_245_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_245_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_246_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_246_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_247_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_247_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_248_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_248_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_249_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_249_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_250_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_250_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_251_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_251_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_252_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_253_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_253_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_254_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_254_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_255_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_255_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_256_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_256_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_257_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_258_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_258_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_259_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_259_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_260_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_260_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_261_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_261_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_262_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_262_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_263_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_263_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_264_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_264_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_265_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_266_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_266_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_267_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_267_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_268_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_268_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_269_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_269_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_270_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_270_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_271_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_271_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_272_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_272_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_273_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_274_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_275_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_276_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_277_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_277_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_278_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_278_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_279_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_280_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_281_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_281_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_282_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_282_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_283_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_283_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_284_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_284_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_285_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_286_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_286_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_287_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_287_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_288_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_288_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_289_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_289_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_290_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_290_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_291_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_291_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_292_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_292_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_293_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_294_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_294_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_295_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_295_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_296_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_296_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_297_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_298_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_298_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_299_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_300_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_300_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_301_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_301_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_302_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_302_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_303_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_304_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_305_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_305_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_307_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_307_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_308_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_308_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_309_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_309_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_310_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_310_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_311_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_311_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_312_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_312_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_313_user_clock2 (.A(clknet_opt_14_user_clock2),
    .X(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_314_user_clock2 (.A(clknet_opt_17_user_clock2),
    .X(clknet_leaf_314_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_315_user_clock2 (.A(clknet_opt_18_user_clock2),
    .X(clknet_leaf_315_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_316_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_316_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_317_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_318_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_318_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_319_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_319_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_320_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_320_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_321_user_clock2 (.A(clknet_opt_19_user_clock2),
    .X(clknet_leaf_321_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_322_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_322_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_325_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_325_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_327_user_clock2 (.A(clknet_opt_8_user_clock2),
    .X(clknet_leaf_327_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_328_user_clock2 (.A(clknet_opt_9_user_clock2),
    .X(clknet_leaf_328_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_329_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_329_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_330_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_330_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_331_user_clock2 (.A(clknet_opt_20_user_clock2),
    .X(clknet_leaf_331_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_332_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_332_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_333_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_333_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_334_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_334_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_335_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_335_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_337_user_clock2 (.A(clknet_opt_4_user_clock2),
    .X(clknet_leaf_337_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_338_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_338_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_339_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_339_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_340_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_340_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_341_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_341_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_342_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_342_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_343_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_343_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_344_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_344_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_345_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_345_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_346_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_346_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_347_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_347_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_348_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_348_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_349_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_349_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_350_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_350_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_351_user_clock2 (.A(clknet_opt_5_user_clock2),
    .X(clknet_leaf_351_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_352_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_352_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_353_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_353_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_354_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_354_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_355_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_355_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_356_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_356_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_357_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_357_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_358_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_358_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_359_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_359_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_360_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_360_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_361_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_361_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_362_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_362_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_363_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_363_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_364_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_364_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_365_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_365_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_366_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_366_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_367_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_367_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_368_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_368_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_369_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_369_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_370_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_370_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_371_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_371_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_372_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_372_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_373_user_clock2 (.A(clknet_5_14_0_user_clock2),
    .X(clknet_leaf_373_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_374_user_clock2 (.A(clknet_5_14_0_user_clock2),
    .X(clknet_leaf_374_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_375_user_clock2 (.A(clknet_5_14_0_user_clock2),
    .X(clknet_leaf_375_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_376_user_clock2 (.A(clknet_5_14_0_user_clock2),
    .X(clknet_leaf_376_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_377_user_clock2 (.A(clknet_5_14_0_user_clock2),
    .X(clknet_leaf_377_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_378_user_clock2 (.A(clknet_5_14_0_user_clock2),
    .X(clknet_leaf_378_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_379_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_379_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_380_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_380_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_381_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_381_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_382_user_clock2 (.A(clknet_5_14_0_user_clock2),
    .X(clknet_leaf_382_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_383_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_383_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_384_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_384_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_385_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_385_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_386_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_386_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_387_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_387_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_388_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_388_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_389_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_389_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_390_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_390_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_391_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_391_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_392_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_392_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_393_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_393_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_394_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_394_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_395_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_395_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_396_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_396_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_397_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_397_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_398_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_398_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_399_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_399_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_400_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_400_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_401_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_401_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_402_user_clock2 (.A(clknet_opt_0_user_clock2),
    .X(clknet_leaf_402_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_403_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_403_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_404_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_404_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_405_user_clock2 (.A(clknet_opt_2_user_clock2),
    .X(clknet_leaf_405_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_406_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_406_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_407_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_407_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_408_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_408_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_409_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_409_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_410_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_410_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_411_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_411_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_412_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_412_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_413_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_413_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_414_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_414_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_415_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_415_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_416_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_416_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_417_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_417_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_418_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_418_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_419_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_419_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_420_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_420_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_421_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_421_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_422_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_422_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_423_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_423_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_424_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_424_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_425_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_425_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_426_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_426_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_427_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_427_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_428_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_428_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_429_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_429_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_430_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_430_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_431_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_431_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_432_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_432_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_433_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_433_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_434_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_434_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_435_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_435_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_436_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_436_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_437_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_437_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_438_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_438_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_439_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_439_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_440_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_440_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_441_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_441_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_442_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_442_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_443_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_443_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_444_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_444_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_445_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_445_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_446_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_446_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_user_clock2 (.A(user_clock2),
    .X(clknet_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_0_user_clock2 (.A(clknet_0_user_clock2),
    .X(clknet_1_0_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_1_user_clock2 (.A(clknet_1_0_0_user_clock2),
    .X(clknet_1_0_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_0_user_clock2 (.A(clknet_0_user_clock2),
    .X(clknet_1_1_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_1_user_clock2 (.A(clknet_1_1_0_user_clock2),
    .X(clknet_1_1_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_0_0_user_clock2 (.A(clknet_1_0_1_user_clock2),
    .X(clknet_2_0_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_0_1_user_clock2 (.A(clknet_2_0_0_user_clock2),
    .X(clknet_2_0_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_1_0_user_clock2 (.A(clknet_1_0_1_user_clock2),
    .X(clknet_2_1_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_1_1_user_clock2 (.A(clknet_2_1_0_user_clock2),
    .X(clknet_2_1_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_2_0_user_clock2 (.A(clknet_1_1_1_user_clock2),
    .X(clknet_2_2_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_2_1_user_clock2 (.A(clknet_2_2_0_user_clock2),
    .X(clknet_2_2_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_3_0_user_clock2 (.A(clknet_1_1_1_user_clock2),
    .X(clknet_2_3_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_3_1_user_clock2 (.A(clknet_2_3_0_user_clock2),
    .X(clknet_2_3_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_0_0_user_clock2 (.A(clknet_2_0_1_user_clock2),
    .X(clknet_3_0_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_1_0_user_clock2 (.A(clknet_2_0_1_user_clock2),
    .X(clknet_3_1_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_2_0_user_clock2 (.A(clknet_2_1_1_user_clock2),
    .X(clknet_3_2_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_3_0_user_clock2 (.A(clknet_2_1_1_user_clock2),
    .X(clknet_3_3_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_4_0_user_clock2 (.A(clknet_2_2_1_user_clock2),
    .X(clknet_3_4_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_5_0_user_clock2 (.A(clknet_2_2_1_user_clock2),
    .X(clknet_3_5_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_6_0_user_clock2 (.A(clknet_2_3_1_user_clock2),
    .X(clknet_3_6_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_7_0_user_clock2 (.A(clknet_2_3_1_user_clock2),
    .X(clknet_3_7_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_0_0_user_clock2 (.A(clknet_3_0_0_user_clock2),
    .X(clknet_4_0_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_1_0_user_clock2 (.A(clknet_3_0_0_user_clock2),
    .X(clknet_4_1_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_2_0_user_clock2 (.A(clknet_3_1_0_user_clock2),
    .X(clknet_4_2_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_3_0_user_clock2 (.A(clknet_3_1_0_user_clock2),
    .X(clknet_4_3_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_4_0_user_clock2 (.A(clknet_3_2_0_user_clock2),
    .X(clknet_4_4_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_5_0_user_clock2 (.A(clknet_3_2_0_user_clock2),
    .X(clknet_4_5_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_6_0_user_clock2 (.A(clknet_3_3_0_user_clock2),
    .X(clknet_4_6_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_7_0_user_clock2 (.A(clknet_3_3_0_user_clock2),
    .X(clknet_4_7_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_8_0_user_clock2 (.A(clknet_3_4_0_user_clock2),
    .X(clknet_4_8_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_9_0_user_clock2 (.A(clknet_3_4_0_user_clock2),
    .X(clknet_4_9_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_10_0_user_clock2 (.A(clknet_3_5_0_user_clock2),
    .X(clknet_4_10_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_11_0_user_clock2 (.A(clknet_3_5_0_user_clock2),
    .X(clknet_4_11_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_12_0_user_clock2 (.A(clknet_3_6_0_user_clock2),
    .X(clknet_4_12_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_13_0_user_clock2 (.A(clknet_3_6_0_user_clock2),
    .X(clknet_4_13_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_14_0_user_clock2 (.A(clknet_3_7_0_user_clock2),
    .X(clknet_4_14_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_15_0_user_clock2 (.A(clknet_3_7_0_user_clock2),
    .X(clknet_4_15_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_0_0_user_clock2 (.A(clknet_4_0_0_user_clock2),
    .X(clknet_5_0_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_1_0_user_clock2 (.A(clknet_4_0_0_user_clock2),
    .X(clknet_5_1_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_2_0_user_clock2 (.A(clknet_4_1_0_user_clock2),
    .X(clknet_5_2_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_3_0_user_clock2 (.A(clknet_4_1_0_user_clock2),
    .X(clknet_5_3_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_4_0_user_clock2 (.A(clknet_4_2_0_user_clock2),
    .X(clknet_5_4_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_5_0_user_clock2 (.A(clknet_4_2_0_user_clock2),
    .X(clknet_5_5_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_6_0_user_clock2 (.A(clknet_4_3_0_user_clock2),
    .X(clknet_5_6_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_7_0_user_clock2 (.A(clknet_4_3_0_user_clock2),
    .X(clknet_5_7_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_8_0_user_clock2 (.A(clknet_4_4_0_user_clock2),
    .X(clknet_5_8_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_9_0_user_clock2 (.A(clknet_4_4_0_user_clock2),
    .X(clknet_5_9_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_10_0_user_clock2 (.A(clknet_4_5_0_user_clock2),
    .X(clknet_5_10_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_11_0_user_clock2 (.A(clknet_4_5_0_user_clock2),
    .X(clknet_5_11_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_12_0_user_clock2 (.A(clknet_4_6_0_user_clock2),
    .X(clknet_5_12_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_13_0_user_clock2 (.A(clknet_4_6_0_user_clock2),
    .X(clknet_5_13_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_14_0_user_clock2 (.A(clknet_4_7_0_user_clock2),
    .X(clknet_5_14_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_15_0_user_clock2 (.A(clknet_4_7_0_user_clock2),
    .X(clknet_5_15_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_16_0_user_clock2 (.A(clknet_4_8_0_user_clock2),
    .X(clknet_5_16_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_17_0_user_clock2 (.A(clknet_4_8_0_user_clock2),
    .X(clknet_5_17_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_18_0_user_clock2 (.A(clknet_4_9_0_user_clock2),
    .X(clknet_5_18_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_19_0_user_clock2 (.A(clknet_4_9_0_user_clock2),
    .X(clknet_5_19_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_20_0_user_clock2 (.A(clknet_4_10_0_user_clock2),
    .X(clknet_5_20_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_21_0_user_clock2 (.A(clknet_4_10_0_user_clock2),
    .X(clknet_5_21_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_22_0_user_clock2 (.A(clknet_4_11_0_user_clock2),
    .X(clknet_5_22_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_23_0_user_clock2 (.A(clknet_4_11_0_user_clock2),
    .X(clknet_5_23_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_24_0_user_clock2 (.A(clknet_4_12_0_user_clock2),
    .X(clknet_5_24_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_25_0_user_clock2 (.A(clknet_4_12_0_user_clock2),
    .X(clknet_5_25_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_26_0_user_clock2 (.A(clknet_4_13_0_user_clock2),
    .X(clknet_5_26_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_27_0_user_clock2 (.A(clknet_4_13_0_user_clock2),
    .X(clknet_5_27_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_28_0_user_clock2 (.A(clknet_4_14_0_user_clock2),
    .X(clknet_5_28_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_29_0_user_clock2 (.A(clknet_4_14_0_user_clock2),
    .X(clknet_5_29_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_30_0_user_clock2 (.A(clknet_4_15_0_user_clock2),
    .X(clknet_5_30_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_31_0_user_clock2 (.A(clknet_4_15_0_user_clock2),
    .X(clknet_5_31_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_0_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_opt_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_opt_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_opt_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_3_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_opt_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_4_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_opt_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_5_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_opt_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_6_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_opt_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_7_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_opt_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_8_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_opt_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_9_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_opt_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_10_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_opt_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_11_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_opt_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_12_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_opt_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_13_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_opt_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_14_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_opt_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_15_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_opt_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_16_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_opt_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_17_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_opt_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_18_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_opt_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_19_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_opt_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_20_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_opt_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_21_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_opt_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
endmodule
