module user_project_wrapper (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    vccd1,
    vssd1,
    vccd2,
    vssd2,
    vdda1,
    vssa1,
    vdda2,
    vssa2,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input vccd1;
 input vssd1;
 input vccd2;
 input vssd2;
 input vdda1;
 input vssa1;
 input vdda2;
 input vssa2;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 sky130_fd_sc_hd__inv_2 _08563_ (.A(\design_top.DATAO[30] ),
    .Y(_06655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08564_ (.A(_06655_),
    .X(_06656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08565_ (.A(_06656_),
    .X(_06657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08566_ (.A(\design_top.DACK[0] ),
    .Y(_02944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08567_ (.A(\design_top.core0.FLUSH[1] ),
    .Y(_06658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08568_ (.A(\design_top.core0.FLUSH[0] ),
    .Y(_06659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _08569_ (.A(_06658_),
    .B(_06659_),
    .C(\design_top.core0.XLCC ),
    .X(_06660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08570_ (.A(_06660_),
    .X(io_out[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08571_ (.A1(\design_top.DACK[1] ),
    .A2(_02944_),
    .B1(io_out[12]),
    .Y(_06661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08572_ (.A(_06661_),
    .Y(_06662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08573_ (.A(\design_top.core0.FLUSH[1] ),
    .B(\design_top.core0.FLUSH[0] ),
    .X(_06663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08574_ (.A(_06663_),
    .Y(_00786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _08575_ (.A(\design_top.core0.XSCC ),
    .B(_00786_),
    .Y(_06664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08576_ (.A(\design_top.core0.SIMM[30] ),
    .Y(_01338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08577_ (.A(_00856_),
    .X(_06665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08578_ (.A(_06665_),
    .Y(_06666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08579_ (.A1(\design_top.core0.SIMM[30] ),
    .A2(_06665_),
    .B1(_01338_),
    .B2(_06666_),
    .X(_06667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08580_ (.A(\design_top.core0.SIMM[29] ),
    .X(_06668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08581_ (.A(_00870_),
    .X(_06669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08582_ (.A(\design_top.core0.SIMM[29] ),
    .B(_00870_),
    .Y(_06670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _08583_ (.A1(_06668_),
    .A2(_06669_),
    .B1(_06670_),
    .Y(_06671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08584_ (.A(_06671_),
    .Y(_06672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08585_ (.A(\design_top.core0.SIMM[28] ),
    .Y(_01340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08586_ (.A(_00884_),
    .Y(_06673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08587_ (.A(\design_top.core0.SIMM[28] ),
    .X(_06674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08588_ (.A1(_01340_),
    .A2(_06673_),
    .B1(_06674_),
    .B2(_00884_),
    .X(_06675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08589_ (.A(_06675_),
    .Y(_06676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08590_ (.A(\design_top.core0.SIMM[26] ),
    .Y(_06677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08591_ (.A(_00911_),
    .Y(_06678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08592_ (.A1(\design_top.core0.SIMM[26] ),
    .A2(_00911_),
    .B1(_06677_),
    .B2(_06678_),
    .X(_06679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08593_ (.A(\design_top.core0.SIMM[27] ),
    .B(_00897_),
    .Y(_06680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _08594_ (.A1(\design_top.core0.SIMM[27] ),
    .A2(_00897_),
    .B1(_06680_),
    .X(_06681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08595_ (.A(_06679_),
    .B(_06681_),
    .X(_06682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08596_ (.A(\design_top.core0.SIMM[25] ),
    .X(_06683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08597_ (.A(_00924_),
    .X(_06684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08598_ (.A(\design_top.core0.SIMM[24] ),
    .X(_06685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08599_ (.A(_00938_),
    .X(_06686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08600_ (.A1(_06685_),
    .A2(_06686_),
    .B1(_06683_),
    .B2(_06684_),
    .X(_06687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08601_ (.A1(_06683_),
    .A2(_06684_),
    .B1(_06687_),
    .Y(_06688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08602_ (.A(\design_top.core0.SIMM[20] ),
    .Y(_01348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08603_ (.A(_00992_),
    .Y(_06689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08604_ (.A(\design_top.core0.SIMM[20] ),
    .X(_06690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08605_ (.A(_00992_),
    .X(_06691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08606_ (.A1(_01348_),
    .A2(_06689_),
    .B1(_06690_),
    .B2(_06691_),
    .X(_06692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08607_ (.A(_06692_),
    .Y(_06693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08608_ (.A(\design_top.core0.SIMM[21] ),
    .Y(_01347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08609_ (.A(_00978_),
    .Y(_06694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08610_ (.A1(_01347_),
    .A2(_06694_),
    .B1(\design_top.core0.SIMM[21] ),
    .B2(_00978_),
    .X(_06695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08611_ (.A(_06695_),
    .Y(_06696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08612_ (.A(\design_top.core0.SIMM[22] ),
    .Y(_06697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08613_ (.A(_00965_),
    .Y(_06698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08614_ (.A(\design_top.core0.SIMM[22] ),
    .X(_06699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08615_ (.A1(_06697_),
    .A2(_06698_),
    .B1(_06699_),
    .B2(_00965_),
    .X(_06700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08616_ (.A(_06700_),
    .Y(_06701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08617_ (.A(_00951_),
    .X(_06702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08618_ (.A(\design_top.core0.SIMM[23] ),
    .B(_00951_),
    .Y(_06703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _08619_ (.A1(\design_top.core0.SIMM[23] ),
    .A2(_06702_),
    .B1(_06703_),
    .Y(_06704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08620_ (.A(_06704_),
    .Y(_06705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08621_ (.A(_06693_),
    .B(_06696_),
    .C(_06701_),
    .D(_06705_),
    .X(_06706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08622_ (.A(\design_top.core0.SIMM[19] ),
    .B(_01005_),
    .Y(_06707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _08623_ (.A1(\design_top.core0.SIMM[19] ),
    .A2(_01005_),
    .B1(_06707_),
    .Y(_06708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08624_ (.A(_06708_),
    .Y(_06709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08625_ (.A(\design_top.core0.SIMM[18] ),
    .Y(_06710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08626_ (.A(_01019_),
    .Y(_06711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08627_ (.A1(_06710_),
    .A2(_06711_),
    .B1(\design_top.core0.SIMM[18] ),
    .B2(_01019_),
    .X(_06712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08628_ (.A(_06712_),
    .Y(_06713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08629_ (.A(\design_top.core0.SIMM[17] ),
    .X(_06714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08630_ (.A(_01048_),
    .Y(_06715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08631_ (.A(_06715_),
    .X(_06716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08632_ (.A(\design_top.core0.SIMM[16] ),
    .X(_06717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08633_ (.A(_01061_),
    .X(_06718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08634_ (.A1(_06714_),
    .A2(_06716_),
    .B1(_06717_),
    .B2(_06718_),
    .X(_06719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08635_ (.A1(_06714_),
    .A2(_06716_),
    .B1(_06719_),
    .Y(_06720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08636_ (.A(\design_top.core0.SIMM[19] ),
    .Y(_01349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08637_ (.A(_01005_),
    .Y(_06721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _08638_ (.A1(_06710_),
    .A2(_06711_),
    .A3(_06707_),
    .B1(_01349_),
    .B2(_06721_),
    .X(_06722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _08639_ (.A1(_06709_),
    .A2(_06713_),
    .A3(_06720_),
    .B1(_06722_),
    .X(_06723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08640_ (.A(\design_top.core0.SIMM[12] ),
    .Y(_01356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08641_ (.A(_01115_),
    .Y(_06724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08642_ (.A(\design_top.core0.SIMM[12] ),
    .X(_06725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08643_ (.A(_01115_),
    .X(_06726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08644_ (.A1(_01356_),
    .A2(_06724_),
    .B1(_06725_),
    .B2(_06726_),
    .X(_06727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08645_ (.A(_06727_),
    .Y(_06728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08646_ (.A(\design_top.core0.SIMM[13] ),
    .Y(_01355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08647_ (.A(_01101_),
    .Y(_06729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08648_ (.A(\design_top.core0.SIMM[13] ),
    .X(_06730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08649_ (.A1(_01355_),
    .A2(_06729_),
    .B1(_06730_),
    .B2(_01101_),
    .X(_06731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08650_ (.A(_06731_),
    .Y(_06732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08651_ (.A(\design_top.core0.SIMM[14] ),
    .Y(_06733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08652_ (.A(_01088_),
    .Y(_06734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08653_ (.A1(_06733_),
    .A2(_06734_),
    .B1(\design_top.core0.SIMM[14] ),
    .B2(_01088_),
    .X(_06735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08654_ (.A(_06735_),
    .Y(_06736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08655_ (.A(\design_top.core0.SIMM[15] ),
    .B(_01074_),
    .Y(_06737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _08656_ (.A1(\design_top.core0.SIMM[15] ),
    .A2(_01074_),
    .B1(_06737_),
    .Y(_06738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08657_ (.A(_06738_),
    .Y(_06739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08658_ (.A(_06728_),
    .B(_06732_),
    .C(_06736_),
    .D(_06739_),
    .X(_06740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08659_ (.A(\design_top.core0.SIMM[10] ),
    .Y(_06741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08660_ (.A(_01141_),
    .Y(_06742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08661_ (.A1(_06741_),
    .A2(_06742_),
    .B1(\design_top.core0.SIMM[10] ),
    .B2(_01141_),
    .X(_06743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08662_ (.A(_06743_),
    .Y(_06744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08663_ (.A(\design_top.core0.SIMM[11] ),
    .B(_01128_),
    .Y(_06745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _08664_ (.A1(\design_top.core0.SIMM[11] ),
    .A2(_01128_),
    .B1(_06745_),
    .Y(_06746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08665_ (.A(_06746_),
    .Y(_06747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08666_ (.A(\design_top.core0.SIMM[9] ),
    .X(_06748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08667_ (.A(_01164_),
    .X(_06749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08668_ (.A(\design_top.core0.SIMM[8] ),
    .X(_06750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08669_ (.A(_01170_),
    .X(_06751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08670_ (.A1(_06750_),
    .A2(_06751_),
    .B1(\design_top.core0.SIMM[9] ),
    .B2(_06749_),
    .X(_06752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08671_ (.A1(_06748_),
    .A2(_06749_),
    .B1(_06752_),
    .Y(_06753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08672_ (.A(_06742_),
    .X(_01142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08673_ (.A(\design_top.core0.SIMM[11] ),
    .Y(_01357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08674_ (.A(_01128_),
    .X(_06754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08675_ (.A(_06754_),
    .Y(_01540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _08676_ (.A1(_06741_),
    .A2(_01142_),
    .A3(_06745_),
    .B1(_01357_),
    .B2(_01540_),
    .X(_06755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _08677_ (.A1(_06744_),
    .A2(_06747_),
    .A3(_06753_),
    .B1(_06755_),
    .X(_06756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08678_ (.A(\design_top.core0.SIMM[7] ),
    .Y(_01361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08679_ (.A(_01183_),
    .Y(_06757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08680_ (.A(_06757_),
    .X(_01184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08681_ (.A(\design_top.core0.SIMM[6] ),
    .Y(_01336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08682_ (.A(_01197_),
    .Y(_06758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _08683_ (.A1(_01361_),
    .A2(_06757_),
    .B1(_01336_),
    .C1(_06758_),
    .X(_06759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08684_ (.A(\design_top.core0.SIMM[6] ),
    .X(_06760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08685_ (.A(_01197_),
    .X(_06761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08686_ (.A1(_06760_),
    .A2(_06761_),
    .B1(_01336_),
    .B2(_06758_),
    .X(_06762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08687_ (.A(\design_top.core0.SIMM[7] ),
    .X(_06763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08688_ (.A(_01183_),
    .X(_06764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08689_ (.A1(_06763_),
    .A2(_06764_),
    .B1(_01361_),
    .B2(_06757_),
    .X(_06765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08690_ (.A(_06762_),
    .B(_06765_),
    .X(_06766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08691_ (.A(\design_top.core0.SIMM[5] ),
    .X(_06767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08692_ (.A(_01210_),
    .X(_06768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08693_ (.A(_01223_),
    .X(_06769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08694_ (.A1(\design_top.core0.SIMM[5] ),
    .A2(_06768_),
    .B1(\design_top.core0.SIMM[4] ),
    .B2(_06769_),
    .X(_06770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08695_ (.A1(_06767_),
    .A2(_06768_),
    .B1(_06770_),
    .Y(_06771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08696_ (.A(_06766_),
    .B(_06771_),
    .X(_06772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08697_ (.A(\design_top.core0.SIMM[5] ),
    .Y(_01334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08698_ (.A(_01210_),
    .Y(_06773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08699_ (.A1(_01334_),
    .A2(_06773_),
    .B1(\design_top.core0.SIMM[5] ),
    .B2(_01210_),
    .X(_06774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08700_ (.A(_06774_),
    .Y(_06775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08701_ (.A(\design_top.core0.SIMM[4] ),
    .Y(_01332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08702_ (.A(_01223_),
    .Y(_06776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08703_ (.A1(_01332_),
    .A2(_06776_),
    .B1(\design_top.core0.SIMM[4] ),
    .B2(_01223_),
    .X(_06777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08704_ (.A(_06777_),
    .Y(_06778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08705_ (.A(_00818_),
    .X(_06779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08706_ (.A(\design_top.core0.SIMM[1] ),
    .X(_06780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08707_ (.A(_00800_),
    .X(_06781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08708_ (.A(\design_top.core0.SIMM[0] ),
    .Y(_00802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08709_ (.A(_00809_),
    .Y(_06782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08710_ (.A(_00802_),
    .B(_06782_),
    .Y(_06783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _08711_ (.A1_N(_06780_),
    .A2_N(_00800_),
    .B1(\design_top.core0.SIMM[1] ),
    .B2(_00800_),
    .X(_06784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08712_ (.A1(_06780_),
    .A2(_06781_),
    .B1(_06783_),
    .B2(_06784_),
    .X(_06785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08713_ (.A(\design_top.core0.SIMM[2] ),
    .Y(_00819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08714_ (.A(_00432_),
    .X(_06786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08715_ (.A(_00432_),
    .Y(_06787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08716_ (.A1(_00789_),
    .A2(_06786_),
    .B1(_00792_),
    .B2(_06787_),
    .X(_06788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08717_ (.A(_06788_),
    .Y(_00793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08718_ (.A1(_00819_),
    .A2(_00793_),
    .B1(\design_top.core0.SIMM[2] ),
    .B2(_06788_),
    .X(_06789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _08719_ (.A(_06785_),
    .B(_06789_),
    .Y(_06790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08720_ (.A(_06790_),
    .Y(_06791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08721_ (.A(\design_top.core0.SIMM[2] ),
    .X(_06792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08722_ (.A1(_06792_),
    .A2(_06788_),
    .B1(\design_top.core0.SIMM[3] ),
    .B2(_00818_),
    .X(_06793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08723_ (.A1(\design_top.core0.SIMM[3] ),
    .A2(_06779_),
    .B1(_06791_),
    .B2(_06793_),
    .X(_06794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08724_ (.A(_06794_),
    .Y(_06795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08725_ (.A(_06775_),
    .B(_06778_),
    .C(_06766_),
    .D(_06795_),
    .X(_06796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2111a_2 _08726_ (.A1(_01361_),
    .A2(_01184_),
    .B1(_06759_),
    .C1(_06772_),
    .D1(_06796_),
    .X(_06797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08727_ (.A(\design_top.core0.SIMM[8] ),
    .Y(_01360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08728_ (.A(_01170_),
    .Y(_06798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08729_ (.A1(_01360_),
    .A2(_06798_),
    .B1(_06750_),
    .B2(_01170_),
    .X(_06799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08730_ (.A(_06799_),
    .Y(_06800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _08731_ (.A1_N(\design_top.core0.SIMM[9] ),
    .A2_N(_01164_),
    .B1(\design_top.core0.SIMM[9] ),
    .B2(_01164_),
    .X(_06801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08732_ (.A(_06801_),
    .Y(_06802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08733_ (.A(_06800_),
    .B(_06802_),
    .C(_06744_),
    .D(_06747_),
    .X(_06803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08734_ (.A(_06803_),
    .B(_06740_),
    .X(_06804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08735_ (.A(_01101_),
    .X(_06805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08736_ (.A1(_06725_),
    .A2(_06726_),
    .B1(_06730_),
    .B2(_06805_),
    .X(_06806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08737_ (.A1(_06730_),
    .A2(_06805_),
    .B1(_06806_),
    .Y(_06807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08738_ (.A(\design_top.core0.SIMM[15] ),
    .X(_06808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08739_ (.A(_06808_),
    .Y(_01353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08740_ (.A(_01074_),
    .X(_06809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08741_ (.A(_06809_),
    .Y(_06810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _08742_ (.A1(_06733_),
    .A2(_06734_),
    .A3(_06737_),
    .B1(_01353_),
    .B2(_06810_),
    .X(_06811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _08743_ (.A1(_06736_),
    .A2(_06739_),
    .A3(_06807_),
    .B1(_06811_),
    .X(_06812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08744_ (.A1(_06740_),
    .A2(_06756_),
    .B1(_06797_),
    .B2(_06804_),
    .C1(_06812_),
    .X(_06813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08745_ (.A(\design_top.core0.SIMM[17] ),
    .Y(_01351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08746_ (.A1(\design_top.core0.SIMM[17] ),
    .A2(_06715_),
    .B1(_01351_),
    .B2(_01048_),
    .X(_06814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08747_ (.A(\design_top.core0.SIMM[16] ),
    .Y(_01352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08748_ (.A(_01061_),
    .Y(_06815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08749_ (.A1(_01352_),
    .A2(_06815_),
    .B1(\design_top.core0.SIMM[16] ),
    .B2(_01061_),
    .X(_06816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08750_ (.A(_06816_),
    .Y(_06817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08751_ (.A(_06709_),
    .B(_06713_),
    .C(_06814_),
    .D(_06817_),
    .X(_06818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08752_ (.A(_06706_),
    .B(_06818_),
    .X(_06819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08753_ (.A(\design_top.core0.SIMM[21] ),
    .X(_06820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08754_ (.A(_00978_),
    .X(_06821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08755_ (.A1(_06690_),
    .A2(_06691_),
    .B1(_06820_),
    .B2(_06821_),
    .X(_06822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08756_ (.A1(_06820_),
    .A2(_06821_),
    .B1(_06822_),
    .Y(_06823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08757_ (.A(_06697_),
    .X(_01346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08758_ (.A(\design_top.core0.SIMM[23] ),
    .Y(_01345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08759_ (.A(_06702_),
    .Y(_00952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _08760_ (.A1(_01346_),
    .A2(_06698_),
    .A3(_06703_),
    .B1(_01345_),
    .B2(_00952_),
    .X(_06824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _08761_ (.A1(_06701_),
    .A2(_06705_),
    .A3(_06823_),
    .B1(_06824_),
    .X(_06825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08762_ (.A1(_06706_),
    .A2(_06723_),
    .B1(_06813_),
    .B2(_06819_),
    .C1(_06825_),
    .X(_06826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08763_ (.A(\design_top.core0.SIMM[24] ),
    .Y(_01344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08764_ (.A(_00938_),
    .Y(_06827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08765_ (.A1(_01344_),
    .A2(_06827_),
    .B1(_06685_),
    .B2(_06686_),
    .X(_06828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08766_ (.A(_06828_),
    .Y(_06829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08767_ (.A(\design_top.core0.SIMM[25] ),
    .Y(_01343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08768_ (.A(_00924_),
    .Y(_06830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08769_ (.A1(_01343_),
    .A2(_06830_),
    .B1(_06683_),
    .B2(_00924_),
    .X(_06831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08770_ (.A(_06831_),
    .Y(_06832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _08771_ (.A(_06829_),
    .B(_06832_),
    .C(_06682_),
    .X(_06833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08772_ (.A(\design_top.core0.SIMM[27] ),
    .Y(_01341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08773_ (.A(_00897_),
    .Y(_06834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _08774_ (.A1(_06677_),
    .A2(_06678_),
    .A3(_06680_),
    .B1(_01341_),
    .B2(_06834_),
    .X(_06835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08775_ (.A1(_06682_),
    .A2(_06688_),
    .B1(_06826_),
    .B2(_06833_),
    .C1(_06835_),
    .X(_06836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08776_ (.A(\design_top.core0.SIMM[29] ),
    .Y(_01339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08777_ (.A(_00870_),
    .Y(_06837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _08778_ (.A1(_01340_),
    .A2(_06673_),
    .A3(_06670_),
    .B1(_01339_),
    .B2(_06837_),
    .X(_06838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _08779_ (.A1(_06672_),
    .A2(_06676_),
    .A3(_06836_),
    .B1(_06838_),
    .X(_06839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _08780_ (.A1(_01338_),
    .A2(_06666_),
    .B1(_06667_),
    .B2(_06839_),
    .Y(_06840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08781_ (.A(_00843_),
    .Y(_06841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08782_ (.A(\design_top.core0.SIMM[31] ),
    .Y(_00763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08783_ (.A1(\design_top.core0.SIMM[31] ),
    .A2(_06841_),
    .B1(_00763_),
    .B2(_00843_),
    .X(_06842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08784_ (.A1_N(_06840_),
    .A2_N(_06842_),
    .B1(_06840_),
    .B2(_06842_),
    .X(\design_top.DADDR[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _08785_ (.A(_06662_),
    .B(_06664_),
    .C(\design_top.DADDR[31] ),
    .X(_06843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08786_ (.A(_01374_),
    .B(_06843_),
    .X(_06844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08787_ (.A(_06844_),
    .X(_06845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08788_ (.A(_06845_),
    .X(_06846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08789_ (.A(\design_top.core0.SIMM[3] ),
    .X(_06847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08790_ (.A(_06847_),
    .Y(_00811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08791_ (.A(_06779_),
    .Y(_06848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08792_ (.A1(_00811_),
    .A2(_06848_),
    .B1(_06847_),
    .B2(_06779_),
    .X(_06849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _08793_ (.A1(_00819_),
    .A2(_00793_),
    .B1(_06790_),
    .X(_06850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08794_ (.A1_N(_06849_),
    .A2_N(_06850_),
    .B1(_06849_),
    .B2(_06850_),
    .X(_00820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08795_ (.A(_00820_),
    .Y(\design_top.DADDR[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _08796_ (.A1(_06785_),
    .A2(_06789_),
    .B1(_06790_),
    .Y(_00810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08797_ (.A(\design_top.DADDR[3] ),
    .B(_00810_),
    .X(_06851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _08798_ (.A1(_06794_),
    .A2(_06777_),
    .B1(_06795_),
    .B2(_06778_),
    .X(_06852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08799_ (.A(_06852_),
    .X(_01371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08800_ (.A(\design_top.core0.SIMM[4] ),
    .X(_06853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _08801_ (.A1(_06853_),
    .A2(_06769_),
    .B1(_06794_),
    .B2(_06777_),
    .X(_06854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _08802_ (.A1_N(_06774_),
    .A2_N(_06854_),
    .B1(_06774_),
    .B2(_06854_),
    .X(_02480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08803_ (.A(_02480_),
    .Y(_01335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _08804_ (.A1(_06775_),
    .A2(_06778_),
    .A3(_06795_),
    .B1(_06771_),
    .X(_06855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08805_ (.A1_N(_06762_),
    .A2_N(_06855_),
    .B1(_06762_),
    .B2(_06855_),
    .X(_01337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08806_ (.A(_01337_),
    .Y(_02484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08807_ (.A(_01335_),
    .B(_02484_),
    .X(_06856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08808_ (.A(_01371_),
    .B(_06856_),
    .X(_06857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08809_ (.A(_06851_),
    .B(_06857_),
    .X(_06858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08810_ (.A(_06846_),
    .B(_06858_),
    .X(_06859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08811_ (.A(_06859_),
    .X(_06860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08812_ (.A(\design_top.XRES ),
    .Y(_06861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08813_ (.A(_06861_),
    .X(_06862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08814_ (.A(wbs_we_i),
    .Y(_06863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _08815_ (.A(_06862_),
    .B(_06863_),
    .C_N(wbs_sel_i[1]),
    .X(_06864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08816_ (.A(_06864_),
    .X(_06865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08817_ (.A(_06865_),
    .X(_06866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08818_ (.A(wbs_adr_i[1]),
    .Y(_06867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _08819_ (.A(wbs_adr_i[2]),
    .B(_06867_),
    .C(wbs_adr_i[0]),
    .X(_06868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08820_ (.A(_06868_),
    .X(_06869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08821_ (.A(_06869_),
    .X(_06870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _08822_ (.A1(_06866_),
    .A2(_06870_),
    .B1(_06859_),
    .X(_06871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08823_ (.A(_06871_),
    .X(_06872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08824_ (.A1_N(_06657_),
    .A2_N(_06860_),
    .B1(\design_top.MEM[9][30] ),
    .B2(_06872_),
    .X(_05493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08825_ (.A(\design_top.DATAO[29] ),
    .Y(_06873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08826_ (.A(_06873_),
    .X(_06874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08827_ (.A(_06874_),
    .X(_06875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08828_ (.A1_N(_06875_),
    .A2_N(_06860_),
    .B1(\design_top.MEM[9][29] ),
    .B2(_06872_),
    .X(_05492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08829_ (.A(\design_top.DATAO[28] ),
    .Y(_06876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08830_ (.A(_06876_),
    .X(_06877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08831_ (.A(_06877_),
    .X(_06878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08832_ (.A1_N(_06878_),
    .A2_N(_06860_),
    .B1(\design_top.MEM[9][28] ),
    .B2(_06872_),
    .X(_05491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08833_ (.A(\design_top.DATAO[27] ),
    .Y(_06879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08834_ (.A(_06879_),
    .X(_06880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08835_ (.A(_06880_),
    .X(_06881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08836_ (.A1_N(_06881_),
    .A2_N(_06860_),
    .B1(\design_top.MEM[9][27] ),
    .B2(_06872_),
    .X(_05490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08837_ (.A(\design_top.DATAO[26] ),
    .Y(_06882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08838_ (.A(_06882_),
    .X(_06883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08839_ (.A(_06883_),
    .X(_06884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08840_ (.A1_N(_06884_),
    .A2_N(_06860_),
    .B1(\design_top.MEM[9][26] ),
    .B2(_06872_),
    .X(_05489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08841_ (.A(\design_top.DATAO[25] ),
    .Y(_06885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08842_ (.A(_06885_),
    .X(_06886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08843_ (.A(_06886_),
    .X(_06887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08844_ (.A1_N(_06887_),
    .A2_N(_06859_),
    .B1(\design_top.MEM[9][25] ),
    .B2(_06871_),
    .X(_05488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08845_ (.A(\design_top.DATAO[24] ),
    .Y(_06888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08846_ (.A(_06888_),
    .X(_06889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08847_ (.A(_06889_),
    .X(_06890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08848_ (.A1_N(_06890_),
    .A2_N(_06859_),
    .B1(\design_top.MEM[9][24] ),
    .B2(_06871_),
    .X(_05487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08849_ (.A(\design_top.DATAO[31] ),
    .Y(_06891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08850_ (.A(_06891_),
    .X(_06892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08851_ (.A(_06892_),
    .X(_06893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08852_ (.A(_00810_),
    .Y(\design_top.DADDR[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08853_ (.A(\design_top.DADDR[3] ),
    .B(\design_top.DADDR[2] ),
    .X(_06894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08854_ (.A(_02480_),
    .B(_02484_),
    .X(_06895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08855_ (.A(_01371_),
    .B(_06895_),
    .X(_06896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08856_ (.A(_06894_),
    .B(_06896_),
    .X(_06897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08857_ (.A(_06846_),
    .B(_06897_),
    .X(_06898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08858_ (.A(_06898_),
    .X(_06899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _08859_ (.A(_06861_),
    .B(_06863_),
    .C_N(wbs_sel_i[0]),
    .X(_06900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08860_ (.A(_06900_),
    .X(_06901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08861_ (.A(_06901_),
    .X(_06902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _08862_ (.A(wbs_adr_i[2]),
    .B(wbs_adr_i[1]),
    .C(wbs_adr_i[0]),
    .X(_06903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08863_ (.A(_06903_),
    .X(_06904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08864_ (.A(_06904_),
    .X(_06905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _08865_ (.A1(_06902_),
    .A2(_06905_),
    .B1(_06898_),
    .X(_06906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08866_ (.A(_06906_),
    .X(_06907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08867_ (.A1_N(_06893_),
    .A2_N(_06899_),
    .B1(\design_top.MEM[0][31] ),
    .B2(_06907_),
    .X(_05486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08868_ (.A1_N(_06657_),
    .A2_N(_06899_),
    .B1(\design_top.MEM[0][30] ),
    .B2(_06907_),
    .X(_05485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08869_ (.A1_N(_06875_),
    .A2_N(_06899_),
    .B1(\design_top.MEM[0][29] ),
    .B2(_06907_),
    .X(_05484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08870_ (.A1_N(_06878_),
    .A2_N(_06899_),
    .B1(\design_top.MEM[0][28] ),
    .B2(_06907_),
    .X(_05483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08871_ (.A1_N(_06881_),
    .A2_N(_06899_),
    .B1(\design_top.MEM[0][27] ),
    .B2(_06907_),
    .X(_05482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08872_ (.A1_N(_06884_),
    .A2_N(_06898_),
    .B1(\design_top.MEM[0][26] ),
    .B2(_06906_),
    .X(_05481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08873_ (.A1_N(_06887_),
    .A2_N(_06898_),
    .B1(\design_top.MEM[0][25] ),
    .B2(_06906_),
    .X(_05480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08874_ (.A1_N(_06890_),
    .A2_N(_06898_),
    .B1(\design_top.MEM[0][24] ),
    .B2(_06906_),
    .X(_05479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08875_ (.A(\design_top.DATAO[15] ),
    .Y(_06908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08876_ (.A(_06908_),
    .X(_06909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08877_ (.A(_06909_),
    .X(_06910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08878_ (.A(_01380_),
    .B(_06843_),
    .X(_06911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08879_ (.A(_06911_),
    .X(_06912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08880_ (.A(_06912_),
    .X(_06913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08881_ (.A(_06897_),
    .B(_06913_),
    .X(_06914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08882_ (.A(_06914_),
    .X(_06915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _08883_ (.A1(_06902_),
    .A2(_06905_),
    .B1(_06914_),
    .X(_06916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08884_ (.A(_06916_),
    .X(_06917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08885_ (.A1_N(_06910_),
    .A2_N(_06915_),
    .B1(\design_top.MEM[0][15] ),
    .B2(_06917_),
    .X(_05478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08886_ (.A(\design_top.DATAO[14] ),
    .Y(_06918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08887_ (.A(_06918_),
    .X(_06919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08888_ (.A(_06919_),
    .X(_06920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08889_ (.A1_N(_06920_),
    .A2_N(_06915_),
    .B1(\design_top.MEM[0][14] ),
    .B2(_06917_),
    .X(_05477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08890_ (.A(\design_top.DATAO[13] ),
    .Y(_06921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08891_ (.A(_06921_),
    .X(_06922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08892_ (.A(_06922_),
    .X(_06923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08893_ (.A1_N(_06923_),
    .A2_N(_06915_),
    .B1(\design_top.MEM[0][13] ),
    .B2(_06917_),
    .X(_05476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08894_ (.A(\design_top.DATAO[12] ),
    .Y(_06924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08895_ (.A(_06924_),
    .X(_06925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08896_ (.A(_06925_),
    .X(_06926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08897_ (.A1_N(_06926_),
    .A2_N(_06915_),
    .B1(\design_top.MEM[0][12] ),
    .B2(_06917_),
    .X(_05475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08898_ (.A(\design_top.DATAO[11] ),
    .Y(_06927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08899_ (.A(_06927_),
    .X(_06928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08900_ (.A(_06928_),
    .X(_06929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08901_ (.A1_N(_06929_),
    .A2_N(_06915_),
    .B1(\design_top.MEM[0][11] ),
    .B2(_06917_),
    .X(_05474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08902_ (.A(\design_top.DATAO[10] ),
    .Y(_06930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08903_ (.A(_06930_),
    .X(_06931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08904_ (.A(_06931_),
    .X(_06932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08905_ (.A1_N(_06932_),
    .A2_N(_06914_),
    .B1(\design_top.MEM[0][10] ),
    .B2(_06916_),
    .X(_05473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08906_ (.A(\design_top.DATAO[9] ),
    .Y(_06933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08907_ (.A(_06933_),
    .X(_06934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08908_ (.A(_06934_),
    .X(_06935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08909_ (.A1_N(_06935_),
    .A2_N(_06914_),
    .B1(\design_top.MEM[0][9] ),
    .B2(_06916_),
    .X(_05472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08910_ (.A(\design_top.DATAO[8] ),
    .Y(_06936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08911_ (.A(_06936_),
    .X(_06937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08912_ (.A(_06937_),
    .X(_06938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08913_ (.A1_N(_06938_),
    .A2_N(_06914_),
    .B1(\design_top.MEM[0][8] ),
    .B2(_06916_),
    .X(_05471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08914_ (.A(\design_top.DATAO[23] ),
    .Y(_06939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08915_ (.A(_06939_),
    .X(_06940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08916_ (.A(_06940_),
    .X(_06941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08917_ (.A(_01369_),
    .B(_06843_),
    .X(_06942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08918_ (.A(_06942_),
    .X(_06943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08919_ (.A(_06943_),
    .X(_06944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08920_ (.A(_06897_),
    .B(_06944_),
    .X(_06945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08921_ (.A(_06945_),
    .X(_06946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _08922_ (.A1(_06902_),
    .A2(_06905_),
    .B1(_06945_),
    .X(_06947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08923_ (.A(_06947_),
    .X(_06948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08924_ (.A1_N(_06941_),
    .A2_N(_06946_),
    .B1(\design_top.MEM[0][23] ),
    .B2(_06948_),
    .X(_05470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08925_ (.A(\design_top.DATAO[22] ),
    .Y(_06949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08926_ (.A(_06949_),
    .X(_06950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08927_ (.A(_06950_),
    .X(_06951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08928_ (.A1_N(_06951_),
    .A2_N(_06946_),
    .B1(\design_top.MEM[0][22] ),
    .B2(_06948_),
    .X(_05469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08929_ (.A(\design_top.DATAO[21] ),
    .Y(_06952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08930_ (.A(_06952_),
    .X(_06953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08931_ (.A(_06953_),
    .X(_06954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08932_ (.A1_N(_06954_),
    .A2_N(_06946_),
    .B1(\design_top.MEM[0][21] ),
    .B2(_06948_),
    .X(_05468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08933_ (.A(\design_top.DATAO[20] ),
    .Y(_06955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08934_ (.A(_06955_),
    .X(_06956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08935_ (.A(_06956_),
    .X(_06957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08936_ (.A1_N(_06957_),
    .A2_N(_06946_),
    .B1(\design_top.MEM[0][20] ),
    .B2(_06948_),
    .X(_05467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08937_ (.A(\design_top.DATAO[19] ),
    .Y(_06958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08938_ (.A(_06958_),
    .X(_06959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08939_ (.A(_06959_),
    .X(_06960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08940_ (.A1_N(_06960_),
    .A2_N(_06946_),
    .B1(\design_top.MEM[0][19] ),
    .B2(_06948_),
    .X(_05466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08941_ (.A(\design_top.DATAO[18] ),
    .Y(_06961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08942_ (.A(_06961_),
    .X(_06962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08943_ (.A(_06962_),
    .X(_06963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08944_ (.A1_N(_06963_),
    .A2_N(_06945_),
    .B1(\design_top.MEM[0][18] ),
    .B2(_06947_),
    .X(_05465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08945_ (.A(\design_top.DATAO[17] ),
    .Y(_06964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08946_ (.A(_06964_),
    .X(_06965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08947_ (.A(_06965_),
    .X(_06966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08948_ (.A1_N(_06966_),
    .A2_N(_06945_),
    .B1(\design_top.MEM[0][17] ),
    .B2(_06947_),
    .X(_05464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08949_ (.A(\design_top.DATAO[16] ),
    .Y(_06967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08950_ (.A(_06967_),
    .X(_06968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08951_ (.A(_06968_),
    .X(_06969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08952_ (.A1_N(_06969_),
    .A2_N(_06945_),
    .B1(\design_top.MEM[0][16] ),
    .B2(_06947_),
    .X(_05463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08953_ (.A(_00820_),
    .B(\design_top.DADDR[2] ),
    .X(_06970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08954_ (.A(_06970_),
    .X(_06971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08955_ (.A(_06857_),
    .B(_06971_),
    .X(_06972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08956_ (.A(_06913_),
    .B(_06972_),
    .X(_06973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08957_ (.A(_06973_),
    .X(_06974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08958_ (.A(_06869_),
    .X(_06975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _08959_ (.A(_06861_),
    .B(_06863_),
    .C_N(wbs_sel_i[2]),
    .X(_06976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08960_ (.A(_06976_),
    .X(_06977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08961_ (.A(_06977_),
    .X(_06978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _08962_ (.A1(_06975_),
    .A2(_06978_),
    .B1(_06973_),
    .X(_06979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08963_ (.A(_06979_),
    .X(_06980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08964_ (.A1_N(_06910_),
    .A2_N(_06974_),
    .B1(\design_top.MEM[10][15] ),
    .B2(_06980_),
    .X(_05462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08965_ (.A1_N(_06920_),
    .A2_N(_06974_),
    .B1(\design_top.MEM[10][14] ),
    .B2(_06980_),
    .X(_05461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08966_ (.A1_N(_06923_),
    .A2_N(_06974_),
    .B1(\design_top.MEM[10][13] ),
    .B2(_06980_),
    .X(_05460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08967_ (.A1_N(_06926_),
    .A2_N(_06974_),
    .B1(\design_top.MEM[10][12] ),
    .B2(_06980_),
    .X(_05459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08968_ (.A1_N(_06929_),
    .A2_N(_06974_),
    .B1(\design_top.MEM[10][11] ),
    .B2(_06980_),
    .X(_05458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08969_ (.A1_N(_06932_),
    .A2_N(_06973_),
    .B1(\design_top.MEM[10][10] ),
    .B2(_06979_),
    .X(_05457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08970_ (.A1_N(_06935_),
    .A2_N(_06973_),
    .B1(\design_top.MEM[10][9] ),
    .B2(_06979_),
    .X(_05456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _08971_ (.A1_N(_06938_),
    .A2_N(_06973_),
    .B1(\design_top.MEM[10][8] ),
    .B2(_06979_),
    .X(_05455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08972_ (.A(_06784_),
    .Y(_06981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _08973_ (.A1(_00802_),
    .A2(_06782_),
    .B1(_06783_),
    .Y(_06982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08974_ (.A(_06982_),
    .Y(_06983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08975_ (.A(_06981_),
    .B(_06983_),
    .X(_06984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08976_ (.A(_06894_),
    .X(_06985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08977_ (.A(\design_top.DADDR[31] ),
    .Y(_06986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08978_ (.A(_06664_),
    .B(_06986_),
    .X(_06987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08979_ (.A(_06891_),
    .B(_06984_),
    .C(_06985_),
    .D(_06987_),
    .X(_06988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08980_ (.A(_06988_),
    .Y(_06989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _08981_ (.A(\design_top.IRES[7] ),
    .Y(_06990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08982_ (.A(_06990_),
    .X(_06991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _08983_ (.A(_06991_),
    .X(_06992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _08984_ (.A1(\design_top.IREQ[7] ),
    .A2(_06988_),
    .B1(\design_top.IACK[7] ),
    .B2(_06989_),
    .C1(_06992_),
    .X(_05454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08985_ (.A(\design_top.IOMUX[3][11] ),
    .B(\design_top.IOMUX[3][10] ),
    .C(\design_top.IOMUX[3][9] ),
    .D(\design_top.IOMUX[3][8] ),
    .X(_06993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08986_ (.A(\design_top.IOMUX[3][15] ),
    .B(\design_top.IOMUX[3][14] ),
    .C(\design_top.IOMUX[3][13] ),
    .D(\design_top.IOMUX[3][12] ),
    .X(_06994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08987_ (.A(\design_top.IOMUX[3][3] ),
    .B(\design_top.IOMUX[3][2] ),
    .C(\design_top.IOMUX[3][1] ),
    .D(\design_top.IOMUX[3][0] ),
    .X(_06995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08988_ (.A(\design_top.IOMUX[3][7] ),
    .B(\design_top.IOMUX[3][6] ),
    .C(\design_top.IOMUX[3][5] ),
    .D(\design_top.IOMUX[3][4] ),
    .X(_06996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08989_ (.A(_06993_),
    .B(_06994_),
    .C(_06995_),
    .D(_06996_),
    .X(_06997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08990_ (.A(\design_top.IOMUX[3][27] ),
    .B(\design_top.IOMUX[3][26] ),
    .C(\design_top.IOMUX[3][25] ),
    .D(\design_top.IOMUX[3][24] ),
    .X(_06998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08991_ (.A(\design_top.IOMUX[3][31] ),
    .B(\design_top.IOMUX[3][30] ),
    .C(\design_top.IOMUX[3][29] ),
    .D(\design_top.IOMUX[3][28] ),
    .X(_06999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08992_ (.A(\design_top.IOMUX[3][19] ),
    .B(\design_top.IOMUX[3][18] ),
    .C(\design_top.IOMUX[3][17] ),
    .D(\design_top.IOMUX[3][16] ),
    .X(_07000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08993_ (.A(\design_top.IOMUX[3][23] ),
    .B(\design_top.IOMUX[3][22] ),
    .C(\design_top.IOMUX[3][21] ),
    .D(\design_top.IOMUX[3][20] ),
    .X(_07001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _08994_ (.A(_06998_),
    .B(_06999_),
    .C(_07000_),
    .D(_07001_),
    .X(_07002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _08995_ (.A(_06997_),
    .B(_07002_),
    .Y(_07003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08996_ (.A(\design_top.TIMER[31] ),
    .B(\design_top.TIMER[30] ),
    .X(_07004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08997_ (.A(\design_top.TIMER[1] ),
    .B(\design_top.TIMER[0] ),
    .X(_07005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08998_ (.A(\design_top.TIMER[2] ),
    .B(_07005_),
    .X(_07006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _08999_ (.A(\design_top.TIMER[3] ),
    .B(_07006_),
    .X(_07007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09000_ (.A(\design_top.TIMER[4] ),
    .B(_07007_),
    .X(_07008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09001_ (.A(\design_top.TIMER[5] ),
    .B(_07008_),
    .X(_07009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09002_ (.A(\design_top.TIMER[6] ),
    .B(_07009_),
    .X(_07010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09003_ (.A(\design_top.TIMER[7] ),
    .B(_07010_),
    .X(_07011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09004_ (.A(\design_top.TIMER[8] ),
    .B(_07011_),
    .X(_07012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09005_ (.A(\design_top.TIMER[9] ),
    .B(_07012_),
    .X(_07013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09006_ (.A(\design_top.TIMER[10] ),
    .B(_07013_),
    .X(_07014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09007_ (.A(\design_top.TIMER[11] ),
    .B(_07014_),
    .X(_07015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09008_ (.A(\design_top.TIMER[12] ),
    .B(_07015_),
    .X(_07016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09009_ (.A(\design_top.TIMER[13] ),
    .B(_07016_),
    .X(_07017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09010_ (.A(\design_top.TIMER[14] ),
    .B(_07017_),
    .X(_07018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09011_ (.A(\design_top.TIMER[15] ),
    .B(_07018_),
    .X(_07019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _09012_ (.A(\design_top.TIMER[17] ),
    .B(\design_top.TIMER[16] ),
    .C(_07019_),
    .X(_07020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _09013_ (.A(\design_top.TIMER[19] ),
    .B(\design_top.TIMER[18] ),
    .C(_07020_),
    .X(_07021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _09014_ (.A(\design_top.TIMER[21] ),
    .B(\design_top.TIMER[20] ),
    .C(_07021_),
    .X(_07022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _09015_ (.A(\design_top.TIMER[23] ),
    .B(\design_top.TIMER[22] ),
    .C(_07022_),
    .X(_07023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _09016_ (.A(\design_top.TIMER[25] ),
    .B(\design_top.TIMER[24] ),
    .C(_07023_),
    .X(_07024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09017_ (.A(\design_top.TIMER[26] ),
    .B(_07024_),
    .X(_07025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09018_ (.A(\design_top.TIMER[27] ),
    .B(_07025_),
    .X(_07026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _09019_ (.A(\design_top.TIMER[29] ),
    .B(\design_top.TIMER[28] ),
    .C(_07004_),
    .D(_07026_),
    .X(_07027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09020_ (.A(_07003_),
    .B(_07027_),
    .X(_07028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09021_ (.A(_07028_),
    .Y(_07029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09022_ (.A(\design_top.IACK[7] ),
    .Y(_07030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09023_ (.A(_06990_),
    .X(_07031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09024_ (.A(_07031_),
    .X(_07032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _09025_ (.A1(\design_top.IREQ[7] ),
    .A2(_07029_),
    .B1(_07030_),
    .B2(_07028_),
    .C1(_07032_),
    .X(_05453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09026_ (.A(_06944_),
    .B(_06972_),
    .X(_07033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09027_ (.A(_07033_),
    .X(_07034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09028_ (.A1(_06975_),
    .A2(_06978_),
    .B1(_07033_),
    .X(_07035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09029_ (.A(_07035_),
    .X(_07036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09030_ (.A1_N(_06941_),
    .A2_N(_07034_),
    .B1(\design_top.MEM[10][23] ),
    .B2(_07036_),
    .X(_05452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09031_ (.A1_N(_06951_),
    .A2_N(_07034_),
    .B1(\design_top.MEM[10][22] ),
    .B2(_07036_),
    .X(_05451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09032_ (.A1_N(_06954_),
    .A2_N(_07034_),
    .B1(\design_top.MEM[10][21] ),
    .B2(_07036_),
    .X(_05450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09033_ (.A1_N(_06957_),
    .A2_N(_07034_),
    .B1(\design_top.MEM[10][20] ),
    .B2(_07036_),
    .X(_05449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09034_ (.A1_N(_06960_),
    .A2_N(_07034_),
    .B1(\design_top.MEM[10][19] ),
    .B2(_07036_),
    .X(_05448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09035_ (.A1_N(_06963_),
    .A2_N(_07033_),
    .B1(\design_top.MEM[10][18] ),
    .B2(_07035_),
    .X(_05447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09036_ (.A1_N(_06966_),
    .A2_N(_07033_),
    .B1(\design_top.MEM[10][17] ),
    .B2(_07035_),
    .X(_05446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09037_ (.A1_N(_06969_),
    .A2_N(_07033_),
    .B1(\design_top.MEM[10][16] ),
    .B2(_07035_),
    .X(_05445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09038_ (.A(_06846_),
    .B(_06972_),
    .X(_07037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09039_ (.A(_07037_),
    .X(_07038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09040_ (.A(_06976_),
    .X(_07039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09041_ (.A1(_06975_),
    .A2(_07039_),
    .B1(_07037_),
    .X(_07040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09042_ (.A(_07040_),
    .X(_07041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09043_ (.A1_N(_06893_),
    .A2_N(_07038_),
    .B1(\design_top.MEM[10][31] ),
    .B2(_07041_),
    .X(_05444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09044_ (.A1_N(_06657_),
    .A2_N(_07038_),
    .B1(\design_top.MEM[10][30] ),
    .B2(_07041_),
    .X(_05443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09045_ (.A1_N(_06875_),
    .A2_N(_07038_),
    .B1(\design_top.MEM[10][29] ),
    .B2(_07041_),
    .X(_05442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09046_ (.A1_N(_06878_),
    .A2_N(_07038_),
    .B1(\design_top.MEM[10][28] ),
    .B2(_07041_),
    .X(_05441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09047_ (.A1_N(_06881_),
    .A2_N(_07038_),
    .B1(\design_top.MEM[10][27] ),
    .B2(_07041_),
    .X(_05440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09048_ (.A1_N(_06884_),
    .A2_N(_07037_),
    .B1(\design_top.MEM[10][26] ),
    .B2(_07040_),
    .X(_05439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09049_ (.A1_N(_06887_),
    .A2_N(_07037_),
    .B1(\design_top.MEM[10][25] ),
    .B2(_07040_),
    .X(_05438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09050_ (.A1_N(_06890_),
    .A2_N(_07037_),
    .B1(\design_top.MEM[10][24] ),
    .B2(_07040_),
    .X(_05437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09051_ (.A(_00820_),
    .B(_00810_),
    .X(_07042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09052_ (.A(_07042_),
    .X(_07043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09053_ (.A(_06857_),
    .B(_07043_),
    .X(_07044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09054_ (.A(_06913_),
    .B(_07044_),
    .X(_07045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09055_ (.A(_07045_),
    .X(_07046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _09056_ (.A(_06861_),
    .B(_06863_),
    .C_N(wbs_sel_i[3]),
    .X(_07047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09057_ (.A(_07047_),
    .X(_07048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09058_ (.A(_07048_),
    .X(_07049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09059_ (.A1(_06975_),
    .A2(_07049_),
    .B1(_07045_),
    .X(_07050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09060_ (.A(_07050_),
    .X(_07051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09061_ (.A1_N(_06910_),
    .A2_N(_07046_),
    .B1(\design_top.MEM[11][15] ),
    .B2(_07051_),
    .X(_05436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09062_ (.A1_N(_06920_),
    .A2_N(_07046_),
    .B1(\design_top.MEM[11][14] ),
    .B2(_07051_),
    .X(_05435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09063_ (.A1_N(_06923_),
    .A2_N(_07046_),
    .B1(\design_top.MEM[11][13] ),
    .B2(_07051_),
    .X(_05434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09064_ (.A1_N(_06926_),
    .A2_N(_07046_),
    .B1(\design_top.MEM[11][12] ),
    .B2(_07051_),
    .X(_05433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09065_ (.A1_N(_06929_),
    .A2_N(_07046_),
    .B1(\design_top.MEM[11][11] ),
    .B2(_07051_),
    .X(_05432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09066_ (.A1_N(_06932_),
    .A2_N(_07045_),
    .B1(\design_top.MEM[11][10] ),
    .B2(_07050_),
    .X(_05431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09067_ (.A1_N(_06935_),
    .A2_N(_07045_),
    .B1(\design_top.MEM[11][9] ),
    .B2(_07050_),
    .X(_05430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09068_ (.A1_N(_06938_),
    .A2_N(_07045_),
    .B1(\design_top.MEM[11][8] ),
    .B2(_07050_),
    .X(_05429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09069_ (.A(_06896_),
    .B(_06971_),
    .X(_07052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09070_ (.A(_06846_),
    .B(_07052_),
    .X(_07053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09071_ (.A(_07053_),
    .X(_07054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09072_ (.A(_06904_),
    .X(_07055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09073_ (.A1(_07055_),
    .A2(_07039_),
    .B1(_07053_),
    .X(_07056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09074_ (.A(_07056_),
    .X(_07057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09075_ (.A1_N(_06893_),
    .A2_N(_07054_),
    .B1(\design_top.MEM[2][31] ),
    .B2(_07057_),
    .X(_05428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09076_ (.A1_N(_06657_),
    .A2_N(_07054_),
    .B1(\design_top.MEM[2][30] ),
    .B2(_07057_),
    .X(_05427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09077_ (.A1_N(_06875_),
    .A2_N(_07054_),
    .B1(\design_top.MEM[2][29] ),
    .B2(_07057_),
    .X(_05426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09078_ (.A1_N(_06878_),
    .A2_N(_07054_),
    .B1(\design_top.MEM[2][28] ),
    .B2(_07057_),
    .X(_05425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09079_ (.A1_N(_06881_),
    .A2_N(_07054_),
    .B1(\design_top.MEM[2][27] ),
    .B2(_07057_),
    .X(_05424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09080_ (.A1_N(_06884_),
    .A2_N(_07053_),
    .B1(\design_top.MEM[2][26] ),
    .B2(_07056_),
    .X(_05423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09081_ (.A1_N(_06887_),
    .A2_N(_07053_),
    .B1(\design_top.MEM[2][25] ),
    .B2(_07056_),
    .X(_05422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09082_ (.A1_N(_06890_),
    .A2_N(_07053_),
    .B1(\design_top.MEM[2][24] ),
    .B2(_07056_),
    .X(_05421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09083_ (.A(_06852_),
    .Y(_01333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09084_ (.A(_01335_),
    .B(_01337_),
    .X(_07058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09085_ (.A(_01333_),
    .B(_07058_),
    .X(_07059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09086_ (.A(_06971_),
    .B(_07059_),
    .X(_07060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09087_ (.A(_06913_),
    .B(_07060_),
    .X(_07061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09088_ (.A(_07061_),
    .X(_07062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09089_ (.A(_07039_),
    .X(_07063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09090_ (.A(wbs_adr_i[2]),
    .Y(_07064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _09091_ (.A(wbs_adr_i[0]),
    .Y(_07065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _09092_ (.A(_07064_),
    .B(_06867_),
    .C(_07065_),
    .X(_07066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09093_ (.A(_07066_),
    .X(_07067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09094_ (.A(_07067_),
    .X(_07068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09095_ (.A1(_07063_),
    .A2(_07068_),
    .B1(_07061_),
    .X(_07069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09096_ (.A(_07069_),
    .X(_07070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09097_ (.A1_N(_06910_),
    .A2_N(_07062_),
    .B1(\design_top.MEM[30][15] ),
    .B2(_07070_),
    .X(_05420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09098_ (.A1_N(_06920_),
    .A2_N(_07062_),
    .B1(\design_top.MEM[30][14] ),
    .B2(_07070_),
    .X(_05419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09099_ (.A1_N(_06923_),
    .A2_N(_07062_),
    .B1(\design_top.MEM[30][13] ),
    .B2(_07070_),
    .X(_05418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09100_ (.A1_N(_06926_),
    .A2_N(_07062_),
    .B1(\design_top.MEM[30][12] ),
    .B2(_07070_),
    .X(_05417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09101_ (.A1_N(_06929_),
    .A2_N(_07062_),
    .B1(\design_top.MEM[30][11] ),
    .B2(_07070_),
    .X(_05416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09102_ (.A1_N(_06932_),
    .A2_N(_07061_),
    .B1(\design_top.MEM[30][10] ),
    .B2(_07069_),
    .X(_05415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09103_ (.A1_N(_06935_),
    .A2_N(_07061_),
    .B1(\design_top.MEM[30][9] ),
    .B2(_07069_),
    .X(_05414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09104_ (.A1_N(_06938_),
    .A2_N(_07061_),
    .B1(\design_top.MEM[30][8] ),
    .B2(_07069_),
    .X(_05413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09105_ (.A(_06944_),
    .B(_07060_),
    .X(_07071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09106_ (.A(_07071_),
    .X(_07072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09107_ (.A1(_07063_),
    .A2(_07068_),
    .B1(_07071_),
    .X(_07073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09108_ (.A(_07073_),
    .X(_07074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09109_ (.A1_N(_06941_),
    .A2_N(_07072_),
    .B1(\design_top.MEM[30][23] ),
    .B2(_07074_),
    .X(_05412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09110_ (.A1_N(_06951_),
    .A2_N(_07072_),
    .B1(\design_top.MEM[30][22] ),
    .B2(_07074_),
    .X(_05411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09111_ (.A1_N(_06954_),
    .A2_N(_07072_),
    .B1(\design_top.MEM[30][21] ),
    .B2(_07074_),
    .X(_05410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09112_ (.A1_N(_06957_),
    .A2_N(_07072_),
    .B1(\design_top.MEM[30][20] ),
    .B2(_07074_),
    .X(_05409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09113_ (.A1_N(_06960_),
    .A2_N(_07072_),
    .B1(\design_top.MEM[30][19] ),
    .B2(_07074_),
    .X(_05408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09114_ (.A1_N(_06963_),
    .A2_N(_07071_),
    .B1(\design_top.MEM[30][18] ),
    .B2(_07073_),
    .X(_05407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09115_ (.A1_N(_06966_),
    .A2_N(_07071_),
    .B1(\design_top.MEM[30][17] ),
    .B2(_07073_),
    .X(_05406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09116_ (.A1_N(_06969_),
    .A2_N(_07071_),
    .B1(\design_top.MEM[30][16] ),
    .B2(_07073_),
    .X(_05405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09117_ (.A(_06846_),
    .B(_07060_),
    .X(_07075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09118_ (.A(_07075_),
    .X(_07076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09119_ (.A1(_07063_),
    .A2(_07068_),
    .B1(_07075_),
    .X(_07077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09120_ (.A(_07077_),
    .X(_07078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09121_ (.A1_N(_06893_),
    .A2_N(_07076_),
    .B1(\design_top.MEM[30][31] ),
    .B2(_07078_),
    .X(_05404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09122_ (.A1_N(_06657_),
    .A2_N(_07076_),
    .B1(\design_top.MEM[30][30] ),
    .B2(_07078_),
    .X(_05403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09123_ (.A1_N(_06875_),
    .A2_N(_07076_),
    .B1(\design_top.MEM[30][29] ),
    .B2(_07078_),
    .X(_05402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09124_ (.A1_N(_06878_),
    .A2_N(_07076_),
    .B1(\design_top.MEM[30][28] ),
    .B2(_07078_),
    .X(_05401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09125_ (.A1_N(_06881_),
    .A2_N(_07076_),
    .B1(\design_top.MEM[30][27] ),
    .B2(_07078_),
    .X(_05400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09126_ (.A1_N(_06884_),
    .A2_N(_07075_),
    .B1(\design_top.MEM[30][26] ),
    .B2(_07077_),
    .X(_05399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09127_ (.A1_N(_06887_),
    .A2_N(_07075_),
    .B1(\design_top.MEM[30][25] ),
    .B2(_07077_),
    .X(_05398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09128_ (.A1_N(_06890_),
    .A2_N(_07075_),
    .B1(\design_top.MEM[30][24] ),
    .B2(_07077_),
    .X(_05397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09129_ (.A(_06912_),
    .X(_07079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09130_ (.A(_07043_),
    .B(_07059_),
    .X(_07080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09131_ (.A(_07079_),
    .B(_07080_),
    .X(_07081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09132_ (.A(_07081_),
    .X(_07082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09133_ (.A(_07047_),
    .X(_07083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09134_ (.A(_07083_),
    .X(_07084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09135_ (.A1(_07084_),
    .A2(_07068_),
    .B1(_07081_),
    .X(_07085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09136_ (.A(_07085_),
    .X(_07086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09137_ (.A1_N(_06910_),
    .A2_N(_07082_),
    .B1(\design_top.MEM[31][15] ),
    .B2(_07086_),
    .X(_05396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09138_ (.A1_N(_06920_),
    .A2_N(_07082_),
    .B1(\design_top.MEM[31][14] ),
    .B2(_07086_),
    .X(_05395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09139_ (.A1_N(_06923_),
    .A2_N(_07082_),
    .B1(\design_top.MEM[31][13] ),
    .B2(_07086_),
    .X(_05394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09140_ (.A1_N(_06926_),
    .A2_N(_07082_),
    .B1(\design_top.MEM[31][12] ),
    .B2(_07086_),
    .X(_05393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09141_ (.A1_N(_06929_),
    .A2_N(_07082_),
    .B1(\design_top.MEM[31][11] ),
    .B2(_07086_),
    .X(_05392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09142_ (.A1_N(_06932_),
    .A2_N(_07081_),
    .B1(\design_top.MEM[31][10] ),
    .B2(_07085_),
    .X(_05391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09143_ (.A1_N(_06935_),
    .A2_N(_07081_),
    .B1(\design_top.MEM[31][9] ),
    .B2(_07085_),
    .X(_05390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09144_ (.A1_N(_06938_),
    .A2_N(_07081_),
    .B1(\design_top.MEM[31][8] ),
    .B2(_07085_),
    .X(_05389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09145_ (.A(_06944_),
    .B(_07080_),
    .X(_07087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09146_ (.A(_07087_),
    .X(_07088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09147_ (.A1(_07084_),
    .A2(_07068_),
    .B1(_07087_),
    .X(_07089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09148_ (.A(_07089_),
    .X(_07090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09149_ (.A1_N(_06941_),
    .A2_N(_07088_),
    .B1(\design_top.MEM[31][23] ),
    .B2(_07090_),
    .X(_05388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09150_ (.A1_N(_06951_),
    .A2_N(_07088_),
    .B1(\design_top.MEM[31][22] ),
    .B2(_07090_),
    .X(_05387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09151_ (.A1_N(_06954_),
    .A2_N(_07088_),
    .B1(\design_top.MEM[31][21] ),
    .B2(_07090_),
    .X(_05386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09152_ (.A1_N(_06957_),
    .A2_N(_07088_),
    .B1(\design_top.MEM[31][20] ),
    .B2(_07090_),
    .X(_05385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09153_ (.A1_N(_06960_),
    .A2_N(_07088_),
    .B1(\design_top.MEM[31][19] ),
    .B2(_07090_),
    .X(_05384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09154_ (.A1_N(_06963_),
    .A2_N(_07087_),
    .B1(\design_top.MEM[31][18] ),
    .B2(_07089_),
    .X(_05383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09155_ (.A1_N(_06966_),
    .A2_N(_07087_),
    .B1(\design_top.MEM[31][17] ),
    .B2(_07089_),
    .X(_05382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09156_ (.A1_N(_06969_),
    .A2_N(_07087_),
    .B1(\design_top.MEM[31][16] ),
    .B2(_07089_),
    .X(_05381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09157_ (.A(_06845_),
    .X(_07091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09158_ (.A(_07091_),
    .B(_07080_),
    .X(_07092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09159_ (.A(_07092_),
    .X(_07093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09160_ (.A(_07067_),
    .X(_07094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09161_ (.A1(_07084_),
    .A2(_07094_),
    .B1(_07092_),
    .X(_07095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09162_ (.A(_07095_),
    .X(_07096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09163_ (.A1_N(_06893_),
    .A2_N(_07093_),
    .B1(\design_top.MEM[31][31] ),
    .B2(_07096_),
    .X(_05380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09164_ (.A(_06656_),
    .X(_07097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09165_ (.A1_N(_07097_),
    .A2_N(_07093_),
    .B1(\design_top.MEM[31][30] ),
    .B2(_07096_),
    .X(_05379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09166_ (.A(_06874_),
    .X(_07098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09167_ (.A1_N(_07098_),
    .A2_N(_07093_),
    .B1(\design_top.MEM[31][29] ),
    .B2(_07096_),
    .X(_05378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09168_ (.A(_06877_),
    .X(_07099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09169_ (.A1_N(_07099_),
    .A2_N(_07093_),
    .B1(\design_top.MEM[31][28] ),
    .B2(_07096_),
    .X(_05377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09170_ (.A(_06880_),
    .X(_07100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09171_ (.A1_N(_07100_),
    .A2_N(_07093_),
    .B1(\design_top.MEM[31][27] ),
    .B2(_07096_),
    .X(_05376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09172_ (.A(_06883_),
    .X(_07101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09173_ (.A1_N(_07101_),
    .A2_N(_07092_),
    .B1(\design_top.MEM[31][26] ),
    .B2(_07095_),
    .X(_05375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09174_ (.A(_06886_),
    .X(_07102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09175_ (.A1_N(_07102_),
    .A2_N(_07092_),
    .B1(\design_top.MEM[31][25] ),
    .B2(_07095_),
    .X(_05374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09176_ (.A(_06889_),
    .X(_07103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09177_ (.A1_N(_07103_),
    .A2_N(_07092_),
    .B1(\design_top.MEM[31][24] ),
    .B2(_07095_),
    .X(_05373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09178_ (.A(_06909_),
    .X(_07104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09179_ (.A(_06896_),
    .B(_07043_),
    .X(_07105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09180_ (.A(_07079_),
    .B(_07105_),
    .X(_07106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09181_ (.A(_07106_),
    .X(_07107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09182_ (.A1(_07055_),
    .A2(_07049_),
    .B1(_07106_),
    .X(_07108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09183_ (.A(_07108_),
    .X(_07109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09184_ (.A1_N(_07104_),
    .A2_N(_07107_),
    .B1(\design_top.MEM[3][15] ),
    .B2(_07109_),
    .X(_05372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09185_ (.A(_06919_),
    .X(_07110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09186_ (.A1_N(_07110_),
    .A2_N(_07107_),
    .B1(\design_top.MEM[3][14] ),
    .B2(_07109_),
    .X(_05371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09187_ (.A(_06922_),
    .X(_07111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09188_ (.A1_N(_07111_),
    .A2_N(_07107_),
    .B1(\design_top.MEM[3][13] ),
    .B2(_07109_),
    .X(_05370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09189_ (.A(_06925_),
    .X(_07112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09190_ (.A1_N(_07112_),
    .A2_N(_07107_),
    .B1(\design_top.MEM[3][12] ),
    .B2(_07109_),
    .X(_05369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09191_ (.A(_06928_),
    .X(_07113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09192_ (.A1_N(_07113_),
    .A2_N(_07107_),
    .B1(\design_top.MEM[3][11] ),
    .B2(_07109_),
    .X(_05368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09193_ (.A(_06931_),
    .X(_07114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09194_ (.A1_N(_07114_),
    .A2_N(_07106_),
    .B1(\design_top.MEM[3][10] ),
    .B2(_07108_),
    .X(_05367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09195_ (.A(_06934_),
    .X(_07115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09196_ (.A1_N(_07115_),
    .A2_N(_07106_),
    .B1(\design_top.MEM[3][9] ),
    .B2(_07108_),
    .X(_05366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09197_ (.A(_06937_),
    .X(_07116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09198_ (.A1_N(_07116_),
    .A2_N(_07106_),
    .B1(\design_top.MEM[3][8] ),
    .B2(_07108_),
    .X(_05365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09199_ (.A(_06943_),
    .X(_07117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09200_ (.A(_07117_),
    .B(_07105_),
    .X(_07118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09201_ (.A(_07118_),
    .X(_07119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09202_ (.A1(_07055_),
    .A2(_07083_),
    .B1(_07118_),
    .X(_07120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09203_ (.A(_07120_),
    .X(_07121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09204_ (.A1_N(_06941_),
    .A2_N(_07119_),
    .B1(\design_top.MEM[3][23] ),
    .B2(_07121_),
    .X(_05364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09205_ (.A1_N(_06951_),
    .A2_N(_07119_),
    .B1(\design_top.MEM[3][22] ),
    .B2(_07121_),
    .X(_05363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09206_ (.A1_N(_06954_),
    .A2_N(_07119_),
    .B1(\design_top.MEM[3][21] ),
    .B2(_07121_),
    .X(_05362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09207_ (.A1_N(_06957_),
    .A2_N(_07119_),
    .B1(\design_top.MEM[3][20] ),
    .B2(_07121_),
    .X(_05361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09208_ (.A1_N(_06960_),
    .A2_N(_07119_),
    .B1(\design_top.MEM[3][19] ),
    .B2(_07121_),
    .X(_05360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09209_ (.A1_N(_06963_),
    .A2_N(_07118_),
    .B1(\design_top.MEM[3][18] ),
    .B2(_07120_),
    .X(_05359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09210_ (.A1_N(_06966_),
    .A2_N(_07118_),
    .B1(\design_top.MEM[3][17] ),
    .B2(_07120_),
    .X(_05358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09211_ (.A1_N(_06969_),
    .A2_N(_07118_),
    .B1(\design_top.MEM[3][16] ),
    .B2(_07120_),
    .X(_05357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09212_ (.A(_06892_),
    .X(_07122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09213_ (.A(_07091_),
    .B(_07105_),
    .X(_07123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09214_ (.A(_07123_),
    .X(_07124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09215_ (.A1(_07055_),
    .A2(_07083_),
    .B1(_07123_),
    .X(_07125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09216_ (.A(_07125_),
    .X(_07126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09217_ (.A1_N(_07122_),
    .A2_N(_07124_),
    .B1(\design_top.MEM[3][31] ),
    .B2(_07126_),
    .X(_05356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09218_ (.A1_N(_07097_),
    .A2_N(_07124_),
    .B1(\design_top.MEM[3][30] ),
    .B2(_07126_),
    .X(_05355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09219_ (.A1_N(_07098_),
    .A2_N(_07124_),
    .B1(\design_top.MEM[3][29] ),
    .B2(_07126_),
    .X(_05354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09220_ (.A1_N(_07099_),
    .A2_N(_07124_),
    .B1(\design_top.MEM[3][28] ),
    .B2(_07126_),
    .X(_05353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09221_ (.A1_N(_07100_),
    .A2_N(_07124_),
    .B1(\design_top.MEM[3][27] ),
    .B2(_07126_),
    .X(_05352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09222_ (.A1_N(_07101_),
    .A2_N(_07123_),
    .B1(\design_top.MEM[3][26] ),
    .B2(_07125_),
    .X(_05351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09223_ (.A1_N(_07102_),
    .A2_N(_07123_),
    .B1(\design_top.MEM[3][25] ),
    .B2(_07125_),
    .X(_05350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09224_ (.A1_N(_07103_),
    .A2_N(_07123_),
    .B1(\design_top.MEM[3][24] ),
    .B2(_07125_),
    .X(_05349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09225_ (.A(_01333_),
    .B(_06895_),
    .X(_07127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09226_ (.A(_06985_),
    .B(_07127_),
    .X(_07128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09227_ (.A(_07079_),
    .B(_07128_),
    .X(_07129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09228_ (.A(_07129_),
    .X(_07130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _09229_ (.A(wbs_adr_i[2]),
    .B(wbs_adr_i[1]),
    .C(_07065_),
    .X(_07131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09230_ (.A(_07131_),
    .X(_07132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09231_ (.A(_07132_),
    .X(_07133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09232_ (.A1(_06902_),
    .A2(_07133_),
    .B1(_07129_),
    .X(_07134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09233_ (.A(_07134_),
    .X(_07135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09234_ (.A1_N(_07104_),
    .A2_N(_07130_),
    .B1(\design_top.MEM[4][15] ),
    .B2(_07135_),
    .X(_05348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09235_ (.A1_N(_07110_),
    .A2_N(_07130_),
    .B1(\design_top.MEM[4][14] ),
    .B2(_07135_),
    .X(_05347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09236_ (.A1_N(_07111_),
    .A2_N(_07130_),
    .B1(\design_top.MEM[4][13] ),
    .B2(_07135_),
    .X(_05346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09237_ (.A1_N(_07112_),
    .A2_N(_07130_),
    .B1(\design_top.MEM[4][12] ),
    .B2(_07135_),
    .X(_05345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09238_ (.A1_N(_07113_),
    .A2_N(_07130_),
    .B1(\design_top.MEM[4][11] ),
    .B2(_07135_),
    .X(_05344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09239_ (.A1_N(_07114_),
    .A2_N(_07129_),
    .B1(\design_top.MEM[4][10] ),
    .B2(_07134_),
    .X(_05343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09240_ (.A1_N(_07115_),
    .A2_N(_07129_),
    .B1(\design_top.MEM[4][9] ),
    .B2(_07134_),
    .X(_05342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09241_ (.A1_N(_07116_),
    .A2_N(_07129_),
    .B1(\design_top.MEM[4][8] ),
    .B2(_07134_),
    .X(_05341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09242_ (.A(_06940_),
    .X(_07136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09243_ (.A(_07117_),
    .B(_07128_),
    .X(_07137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09244_ (.A(_07137_),
    .X(_07138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09245_ (.A1(_06902_),
    .A2(_07133_),
    .B1(_07137_),
    .X(_07139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09246_ (.A(_07139_),
    .X(_07140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09247_ (.A1_N(_07136_),
    .A2_N(_07138_),
    .B1(\design_top.MEM[4][23] ),
    .B2(_07140_),
    .X(_05340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09248_ (.A(_06950_),
    .X(_07141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09249_ (.A1_N(_07141_),
    .A2_N(_07138_),
    .B1(\design_top.MEM[4][22] ),
    .B2(_07140_),
    .X(_05339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09250_ (.A(_06953_),
    .X(_07142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09251_ (.A1_N(_07142_),
    .A2_N(_07138_),
    .B1(\design_top.MEM[4][21] ),
    .B2(_07140_),
    .X(_05338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09252_ (.A(_06956_),
    .X(_07143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09253_ (.A1_N(_07143_),
    .A2_N(_07138_),
    .B1(\design_top.MEM[4][20] ),
    .B2(_07140_),
    .X(_05337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09254_ (.A(_06959_),
    .X(_07144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09255_ (.A1_N(_07144_),
    .A2_N(_07138_),
    .B1(\design_top.MEM[4][19] ),
    .B2(_07140_),
    .X(_05336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09256_ (.A(_06962_),
    .X(_07145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09257_ (.A1_N(_07145_),
    .A2_N(_07137_),
    .B1(\design_top.MEM[4][18] ),
    .B2(_07139_),
    .X(_05335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09258_ (.A(_06965_),
    .X(_07146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09259_ (.A1_N(_07146_),
    .A2_N(_07137_),
    .B1(\design_top.MEM[4][17] ),
    .B2(_07139_),
    .X(_05334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09260_ (.A(_06968_),
    .X(_07147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09261_ (.A1_N(_07147_),
    .A2_N(_07137_),
    .B1(\design_top.MEM[4][16] ),
    .B2(_07139_),
    .X(_05333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09262_ (.A(_07091_),
    .B(_07128_),
    .X(_07148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09263_ (.A(_07148_),
    .X(_07149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09264_ (.A(_06900_),
    .X(_07150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09265_ (.A(_07150_),
    .X(_07151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09266_ (.A1(_07151_),
    .A2(_07133_),
    .B1(_07148_),
    .X(_07152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09267_ (.A(_07152_),
    .X(_07153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09268_ (.A1_N(_07122_),
    .A2_N(_07149_),
    .B1(\design_top.MEM[4][31] ),
    .B2(_07153_),
    .X(_05332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09269_ (.A1_N(_07097_),
    .A2_N(_07149_),
    .B1(\design_top.MEM[4][30] ),
    .B2(_07153_),
    .X(_05331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09270_ (.A1_N(_07098_),
    .A2_N(_07149_),
    .B1(\design_top.MEM[4][29] ),
    .B2(_07153_),
    .X(_05330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09271_ (.A1_N(_07099_),
    .A2_N(_07149_),
    .B1(\design_top.MEM[4][28] ),
    .B2(_07153_),
    .X(_05329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09272_ (.A1_N(_07100_),
    .A2_N(_07149_),
    .B1(\design_top.MEM[4][27] ),
    .B2(_07153_),
    .X(_05328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09273_ (.A1_N(_07101_),
    .A2_N(_07148_),
    .B1(\design_top.MEM[4][26] ),
    .B2(_07152_),
    .X(_05327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09274_ (.A1_N(_07102_),
    .A2_N(_07148_),
    .B1(\design_top.MEM[4][25] ),
    .B2(_07152_),
    .X(_05326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09275_ (.A1_N(_07103_),
    .A2_N(_07148_),
    .B1(\design_top.MEM[4][24] ),
    .B2(_07152_),
    .X(_05325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09276_ (.A(_06851_),
    .X(_07154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09277_ (.A(_07154_),
    .B(_07127_),
    .X(_07155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09278_ (.A(_07079_),
    .B(_07155_),
    .X(_07156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09279_ (.A(_07156_),
    .X(_07157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09280_ (.A1(_06866_),
    .A2(_07133_),
    .B1(_07156_),
    .X(_07158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09281_ (.A(_07158_),
    .X(_07159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09282_ (.A1_N(_07104_),
    .A2_N(_07157_),
    .B1(\design_top.MEM[5][15] ),
    .B2(_07159_),
    .X(_05324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09283_ (.A1_N(_07110_),
    .A2_N(_07157_),
    .B1(\design_top.MEM[5][14] ),
    .B2(_07159_),
    .X(_05323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09284_ (.A1_N(_07111_),
    .A2_N(_07157_),
    .B1(\design_top.MEM[5][13] ),
    .B2(_07159_),
    .X(_05322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09285_ (.A1_N(_07112_),
    .A2_N(_07157_),
    .B1(\design_top.MEM[5][12] ),
    .B2(_07159_),
    .X(_05321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09286_ (.A1_N(_07113_),
    .A2_N(_07157_),
    .B1(\design_top.MEM[5][11] ),
    .B2(_07159_),
    .X(_05320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09287_ (.A1_N(_07114_),
    .A2_N(_07156_),
    .B1(\design_top.MEM[5][10] ),
    .B2(_07158_),
    .X(_05319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09288_ (.A1_N(_07115_),
    .A2_N(_07156_),
    .B1(\design_top.MEM[5][9] ),
    .B2(_07158_),
    .X(_05318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09289_ (.A1_N(_07116_),
    .A2_N(_07156_),
    .B1(\design_top.MEM[5][8] ),
    .B2(_07158_),
    .X(_05317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09290_ (.A(_07117_),
    .B(_07155_),
    .X(_07160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09291_ (.A(_07160_),
    .X(_07161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09292_ (.A1(_06866_),
    .A2(_07133_),
    .B1(_07160_),
    .X(_07162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09293_ (.A(_07162_),
    .X(_07163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09294_ (.A1_N(_07136_),
    .A2_N(_07161_),
    .B1(\design_top.MEM[5][23] ),
    .B2(_07163_),
    .X(_05316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09295_ (.A1_N(_07141_),
    .A2_N(_07161_),
    .B1(\design_top.MEM[5][22] ),
    .B2(_07163_),
    .X(_05315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09296_ (.A1_N(_07142_),
    .A2_N(_07161_),
    .B1(\design_top.MEM[5][21] ),
    .B2(_07163_),
    .X(_05314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09297_ (.A1_N(_07143_),
    .A2_N(_07161_),
    .B1(\design_top.MEM[5][20] ),
    .B2(_07163_),
    .X(_05313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09298_ (.A1_N(_07144_),
    .A2_N(_07161_),
    .B1(\design_top.MEM[5][19] ),
    .B2(_07163_),
    .X(_05312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09299_ (.A1_N(_07145_),
    .A2_N(_07160_),
    .B1(\design_top.MEM[5][18] ),
    .B2(_07162_),
    .X(_05311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09300_ (.A1_N(_07146_),
    .A2_N(_07160_),
    .B1(\design_top.MEM[5][17] ),
    .B2(_07162_),
    .X(_05310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09301_ (.A1_N(_07147_),
    .A2_N(_07160_),
    .B1(\design_top.MEM[5][16] ),
    .B2(_07162_),
    .X(_05309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09302_ (.A(_07091_),
    .B(_07155_),
    .X(_07164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09303_ (.A(_07164_),
    .X(_07165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09304_ (.A(_07132_),
    .X(_07166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09305_ (.A1(_06866_),
    .A2(_07166_),
    .B1(_07164_),
    .X(_07167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09306_ (.A(_07167_),
    .X(_07168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09307_ (.A1_N(_07122_),
    .A2_N(_07165_),
    .B1(\design_top.MEM[5][31] ),
    .B2(_07168_),
    .X(_05308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09308_ (.A1_N(_07097_),
    .A2_N(_07165_),
    .B1(\design_top.MEM[5][30] ),
    .B2(_07168_),
    .X(_05307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09309_ (.A1_N(_07098_),
    .A2_N(_07165_),
    .B1(\design_top.MEM[5][29] ),
    .B2(_07168_),
    .X(_05306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09310_ (.A1_N(_07099_),
    .A2_N(_07165_),
    .B1(\design_top.MEM[5][28] ),
    .B2(_07168_),
    .X(_05305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09311_ (.A1_N(_07100_),
    .A2_N(_07165_),
    .B1(\design_top.MEM[5][27] ),
    .B2(_07168_),
    .X(_05304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09312_ (.A1_N(_07101_),
    .A2_N(_07164_),
    .B1(\design_top.MEM[5][26] ),
    .B2(_07167_),
    .X(_05303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09313_ (.A1_N(_07102_),
    .A2_N(_07164_),
    .B1(\design_top.MEM[5][25] ),
    .B2(_07167_),
    .X(_05302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09314_ (.A1_N(_07103_),
    .A2_N(_07164_),
    .B1(\design_top.MEM[5][24] ),
    .B2(_07167_),
    .X(_05301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09315_ (.A(_06971_),
    .B(_07127_),
    .X(_07169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09316_ (.A(_07079_),
    .B(_07169_),
    .X(_07170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09317_ (.A(_07170_),
    .X(_07171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09318_ (.A1(_07063_),
    .A2(_07166_),
    .B1(_07170_),
    .X(_07172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09319_ (.A(_07172_),
    .X(_07173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09320_ (.A1_N(_07104_),
    .A2_N(_07171_),
    .B1(\design_top.MEM[6][15] ),
    .B2(_07173_),
    .X(_05300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09321_ (.A1_N(_07110_),
    .A2_N(_07171_),
    .B1(\design_top.MEM[6][14] ),
    .B2(_07173_),
    .X(_05299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09322_ (.A1_N(_07111_),
    .A2_N(_07171_),
    .B1(\design_top.MEM[6][13] ),
    .B2(_07173_),
    .X(_05298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09323_ (.A1_N(_07112_),
    .A2_N(_07171_),
    .B1(\design_top.MEM[6][12] ),
    .B2(_07173_),
    .X(_05297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09324_ (.A1_N(_07113_),
    .A2_N(_07171_),
    .B1(\design_top.MEM[6][11] ),
    .B2(_07173_),
    .X(_05296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09325_ (.A1_N(_07114_),
    .A2_N(_07170_),
    .B1(\design_top.MEM[6][10] ),
    .B2(_07172_),
    .X(_05295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09326_ (.A1_N(_07115_),
    .A2_N(_07170_),
    .B1(\design_top.MEM[6][9] ),
    .B2(_07172_),
    .X(_05294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09327_ (.A1_N(_07116_),
    .A2_N(_07170_),
    .B1(\design_top.MEM[6][8] ),
    .B2(_07172_),
    .X(_05293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09328_ (.A(_07117_),
    .B(_07169_),
    .X(_07174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09329_ (.A(_07174_),
    .X(_07175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09330_ (.A1(_07063_),
    .A2(_07166_),
    .B1(_07174_),
    .X(_07176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09331_ (.A(_07176_),
    .X(_07177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09332_ (.A1_N(_07136_),
    .A2_N(_07175_),
    .B1(\design_top.MEM[6][23] ),
    .B2(_07177_),
    .X(_05292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09333_ (.A1_N(_07141_),
    .A2_N(_07175_),
    .B1(\design_top.MEM[6][22] ),
    .B2(_07177_),
    .X(_05291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09334_ (.A1_N(_07142_),
    .A2_N(_07175_),
    .B1(\design_top.MEM[6][21] ),
    .B2(_07177_),
    .X(_05290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09335_ (.A1_N(_07143_),
    .A2_N(_07175_),
    .B1(\design_top.MEM[6][20] ),
    .B2(_07177_),
    .X(_05289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09336_ (.A1_N(_07144_),
    .A2_N(_07175_),
    .B1(\design_top.MEM[6][19] ),
    .B2(_07177_),
    .X(_05288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09337_ (.A1_N(_07145_),
    .A2_N(_07174_),
    .B1(\design_top.MEM[6][18] ),
    .B2(_07176_),
    .X(_05287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09338_ (.A1_N(_07146_),
    .A2_N(_07174_),
    .B1(\design_top.MEM[6][17] ),
    .B2(_07176_),
    .X(_05286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09339_ (.A1_N(_07147_),
    .A2_N(_07174_),
    .B1(\design_top.MEM[6][16] ),
    .B2(_07176_),
    .X(_05285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09340_ (.A(_01333_),
    .B(_06856_),
    .X(_07178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09341_ (.A(_07154_),
    .B(_07178_),
    .X(_07179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09342_ (.A(_07117_),
    .B(_07179_),
    .X(_07180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09343_ (.A(_07180_),
    .X(_07181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _09344_ (.A(wbs_adr_i[2]),
    .B(_06867_),
    .C(_07065_),
    .X(_07182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09345_ (.A(_07182_),
    .X(_07183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09346_ (.A(_07183_),
    .X(_07184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09347_ (.A1(_06866_),
    .A2(_07184_),
    .B1(_07180_),
    .X(_07185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09348_ (.A(_07185_),
    .X(_07186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09349_ (.A1_N(_07136_),
    .A2_N(_07181_),
    .B1(\design_top.MEM[13][23] ),
    .B2(_07186_),
    .X(_05284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09350_ (.A1_N(_07141_),
    .A2_N(_07181_),
    .B1(\design_top.MEM[13][22] ),
    .B2(_07186_),
    .X(_05283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09351_ (.A1_N(_07142_),
    .A2_N(_07181_),
    .B1(\design_top.MEM[13][21] ),
    .B2(_07186_),
    .X(_05282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09352_ (.A1_N(_07143_),
    .A2_N(_07181_),
    .B1(\design_top.MEM[13][20] ),
    .B2(_07186_),
    .X(_05281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09353_ (.A1_N(_07144_),
    .A2_N(_07181_),
    .B1(\design_top.MEM[13][19] ),
    .B2(_07186_),
    .X(_05280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09354_ (.A1_N(_07145_),
    .A2_N(_07180_),
    .B1(\design_top.MEM[13][18] ),
    .B2(_07185_),
    .X(_05279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09355_ (.A1_N(_07146_),
    .A2_N(_07180_),
    .B1(\design_top.MEM[13][17] ),
    .B2(_07185_),
    .X(_05278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09356_ (.A1_N(_07147_),
    .A2_N(_07180_),
    .B1(\design_top.MEM[13][16] ),
    .B2(_07185_),
    .X(_05277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09357_ (.A(_07091_),
    .B(_07179_),
    .X(_07187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09358_ (.A(_07187_),
    .X(_07188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09359_ (.A(_06864_),
    .X(_07189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09360_ (.A(_07189_),
    .X(_07190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09361_ (.A1(_07190_),
    .A2(_07184_),
    .B1(_07187_),
    .X(_07191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09362_ (.A(_07191_),
    .X(_07192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09363_ (.A1_N(_07122_),
    .A2_N(_07188_),
    .B1(\design_top.MEM[13][31] ),
    .B2(_07192_),
    .X(_05276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09364_ (.A1_N(_07097_),
    .A2_N(_07188_),
    .B1(\design_top.MEM[13][30] ),
    .B2(_07192_),
    .X(_05275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09365_ (.A1_N(_07098_),
    .A2_N(_07188_),
    .B1(\design_top.MEM[13][29] ),
    .B2(_07192_),
    .X(_05274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09366_ (.A1_N(_07099_),
    .A2_N(_07188_),
    .B1(\design_top.MEM[13][28] ),
    .B2(_07192_),
    .X(_05273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09367_ (.A1_N(_07100_),
    .A2_N(_07188_),
    .B1(\design_top.MEM[13][27] ),
    .B2(_07192_),
    .X(_05272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09368_ (.A1_N(_07101_),
    .A2_N(_07187_),
    .B1(\design_top.MEM[13][26] ),
    .B2(_07191_),
    .X(_05271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09369_ (.A1_N(_07102_),
    .A2_N(_07187_),
    .B1(\design_top.MEM[13][25] ),
    .B2(_07191_),
    .X(_05270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09370_ (.A1_N(_07103_),
    .A2_N(_07187_),
    .B1(\design_top.MEM[13][24] ),
    .B2(_07191_),
    .X(_05269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09371_ (.A(_06912_),
    .X(_07193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09372_ (.A(_06971_),
    .B(_07178_),
    .X(_07194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09373_ (.A(_07193_),
    .B(_07194_),
    .X(_07195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09374_ (.A(_07195_),
    .X(_07196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09375_ (.A(_06977_),
    .X(_07197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09376_ (.A1(_07197_),
    .A2(_07184_),
    .B1(_07195_),
    .X(_07198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09377_ (.A(_07198_),
    .X(_07199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09378_ (.A1_N(_07104_),
    .A2_N(_07196_),
    .B1(\design_top.MEM[14][15] ),
    .B2(_07199_),
    .X(_05268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09379_ (.A1_N(_07110_),
    .A2_N(_07196_),
    .B1(\design_top.MEM[14][14] ),
    .B2(_07199_),
    .X(_05267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09380_ (.A1_N(_07111_),
    .A2_N(_07196_),
    .B1(\design_top.MEM[14][13] ),
    .B2(_07199_),
    .X(_05266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09381_ (.A1_N(_07112_),
    .A2_N(_07196_),
    .B1(\design_top.MEM[14][12] ),
    .B2(_07199_),
    .X(_05265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09382_ (.A1_N(_07113_),
    .A2_N(_07196_),
    .B1(\design_top.MEM[14][11] ),
    .B2(_07199_),
    .X(_05264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09383_ (.A1_N(_07114_),
    .A2_N(_07195_),
    .B1(\design_top.MEM[14][10] ),
    .B2(_07198_),
    .X(_05263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09384_ (.A1_N(_07115_),
    .A2_N(_07195_),
    .B1(\design_top.MEM[14][9] ),
    .B2(_07198_),
    .X(_05262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09385_ (.A1_N(_07116_),
    .A2_N(_07195_),
    .B1(\design_top.MEM[14][8] ),
    .B2(_07198_),
    .X(_05261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09386_ (.A(_06943_),
    .X(_07200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09387_ (.A(_07200_),
    .B(_07194_),
    .X(_07201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09388_ (.A(_07201_),
    .X(_07202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09389_ (.A1(_07197_),
    .A2(_07184_),
    .B1(_07201_),
    .X(_07203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09390_ (.A(_07203_),
    .X(_07204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09391_ (.A1_N(_07136_),
    .A2_N(_07202_),
    .B1(\design_top.MEM[14][23] ),
    .B2(_07204_),
    .X(_05260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09392_ (.A1_N(_07141_),
    .A2_N(_07202_),
    .B1(\design_top.MEM[14][22] ),
    .B2(_07204_),
    .X(_05259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09393_ (.A1_N(_07142_),
    .A2_N(_07202_),
    .B1(\design_top.MEM[14][21] ),
    .B2(_07204_),
    .X(_05258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09394_ (.A1_N(_07143_),
    .A2_N(_07202_),
    .B1(\design_top.MEM[14][20] ),
    .B2(_07204_),
    .X(_05257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09395_ (.A1_N(_07144_),
    .A2_N(_07202_),
    .B1(\design_top.MEM[14][19] ),
    .B2(_07204_),
    .X(_05256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09396_ (.A1_N(_07145_),
    .A2_N(_07201_),
    .B1(\design_top.MEM[14][18] ),
    .B2(_07203_),
    .X(_05255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09397_ (.A1_N(_07146_),
    .A2_N(_07201_),
    .B1(\design_top.MEM[14][17] ),
    .B2(_07203_),
    .X(_05254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09398_ (.A1_N(_07147_),
    .A2_N(_07201_),
    .B1(\design_top.MEM[14][16] ),
    .B2(_07203_),
    .X(_05253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09399_ (.A(_06845_),
    .X(_07205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09400_ (.A(_07205_),
    .B(_07194_),
    .X(_07206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09401_ (.A(_07206_),
    .X(_07207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09402_ (.A1(_07197_),
    .A2(_07184_),
    .B1(_07206_),
    .X(_07208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09403_ (.A(_07208_),
    .X(_07209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09404_ (.A1_N(_07122_),
    .A2_N(_07207_),
    .B1(\design_top.MEM[14][31] ),
    .B2(_07209_),
    .X(_05252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09405_ (.A(_06656_),
    .X(_07210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09406_ (.A1_N(_07210_),
    .A2_N(_07207_),
    .B1(\design_top.MEM[14][30] ),
    .B2(_07209_),
    .X(_05251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09407_ (.A(_06874_),
    .X(_07211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09408_ (.A1_N(_07211_),
    .A2_N(_07207_),
    .B1(\design_top.MEM[14][29] ),
    .B2(_07209_),
    .X(_05250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09409_ (.A(_06877_),
    .X(_07212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09410_ (.A1_N(_07212_),
    .A2_N(_07207_),
    .B1(\design_top.MEM[14][28] ),
    .B2(_07209_),
    .X(_05249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09411_ (.A(_06880_),
    .X(_07213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09412_ (.A1_N(_07213_),
    .A2_N(_07207_),
    .B1(\design_top.MEM[14][27] ),
    .B2(_07209_),
    .X(_05248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09413_ (.A(_06883_),
    .X(_07214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09414_ (.A1_N(_07214_),
    .A2_N(_07206_),
    .B1(\design_top.MEM[14][26] ),
    .B2(_07208_),
    .X(_05247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09415_ (.A(_06886_),
    .X(_07215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09416_ (.A1_N(_07215_),
    .A2_N(_07206_),
    .B1(\design_top.MEM[14][25] ),
    .B2(_07208_),
    .X(_05246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09417_ (.A(_06889_),
    .X(_07216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09418_ (.A1_N(_07216_),
    .A2_N(_07206_),
    .B1(\design_top.MEM[14][24] ),
    .B2(_07208_),
    .X(_05245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09419_ (.A(_06909_),
    .X(_07217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09420_ (.A(_07043_),
    .B(_07178_),
    .X(_07218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09421_ (.A(_07193_),
    .B(_07218_),
    .X(_07219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09422_ (.A(_07219_),
    .X(_07220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09423_ (.A(_07183_),
    .X(_07221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09424_ (.A1(_07084_),
    .A2(_07221_),
    .B1(_07219_),
    .X(_07222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09425_ (.A(_07222_),
    .X(_07223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09426_ (.A1_N(_07217_),
    .A2_N(_07220_),
    .B1(\design_top.MEM[15][15] ),
    .B2(_07223_),
    .X(_05244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09427_ (.A(_06919_),
    .X(_07224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09428_ (.A1_N(_07224_),
    .A2_N(_07220_),
    .B1(\design_top.MEM[15][14] ),
    .B2(_07223_),
    .X(_05243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09429_ (.A(_06922_),
    .X(_07225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09430_ (.A1_N(_07225_),
    .A2_N(_07220_),
    .B1(\design_top.MEM[15][13] ),
    .B2(_07223_),
    .X(_05242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09431_ (.A(_06925_),
    .X(_07226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09432_ (.A1_N(_07226_),
    .A2_N(_07220_),
    .B1(\design_top.MEM[15][12] ),
    .B2(_07223_),
    .X(_05241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09433_ (.A(_06928_),
    .X(_07227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09434_ (.A1_N(_07227_),
    .A2_N(_07220_),
    .B1(\design_top.MEM[15][11] ),
    .B2(_07223_),
    .X(_05240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09435_ (.A(_06931_),
    .X(_07228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09436_ (.A1_N(_07228_),
    .A2_N(_07219_),
    .B1(\design_top.MEM[15][10] ),
    .B2(_07222_),
    .X(_05239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09437_ (.A(_06934_),
    .X(_07229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09438_ (.A1_N(_07229_),
    .A2_N(_07219_),
    .B1(\design_top.MEM[15][9] ),
    .B2(_07222_),
    .X(_05238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09439_ (.A(_06937_),
    .X(_07230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09440_ (.A1_N(_07230_),
    .A2_N(_07219_),
    .B1(\design_top.MEM[15][8] ),
    .B2(_07222_),
    .X(_05237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09441_ (.A(_06940_),
    .X(_07231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09442_ (.A(_07200_),
    .B(_07218_),
    .X(_07232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09443_ (.A(_07232_),
    .X(_07233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09444_ (.A1(_07084_),
    .A2(_07221_),
    .B1(_07232_),
    .X(_07234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09445_ (.A(_07234_),
    .X(_07235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09446_ (.A1_N(_07231_),
    .A2_N(_07233_),
    .B1(\design_top.MEM[15][23] ),
    .B2(_07235_),
    .X(_05236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09447_ (.A(_06950_),
    .X(_07236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09448_ (.A1_N(_07236_),
    .A2_N(_07233_),
    .B1(\design_top.MEM[15][22] ),
    .B2(_07235_),
    .X(_05235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09449_ (.A(_06953_),
    .X(_07237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09450_ (.A1_N(_07237_),
    .A2_N(_07233_),
    .B1(\design_top.MEM[15][21] ),
    .B2(_07235_),
    .X(_05234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09451_ (.A(_06956_),
    .X(_07238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09452_ (.A1_N(_07238_),
    .A2_N(_07233_),
    .B1(\design_top.MEM[15][20] ),
    .B2(_07235_),
    .X(_05233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09453_ (.A(_06959_),
    .X(_07239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09454_ (.A1_N(_07239_),
    .A2_N(_07233_),
    .B1(\design_top.MEM[15][19] ),
    .B2(_07235_),
    .X(_05232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09455_ (.A(_06962_),
    .X(_07240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09456_ (.A1_N(_07240_),
    .A2_N(_07232_),
    .B1(\design_top.MEM[15][18] ),
    .B2(_07234_),
    .X(_05231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09457_ (.A(_06965_),
    .X(_07241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09458_ (.A1_N(_07241_),
    .A2_N(_07232_),
    .B1(\design_top.MEM[15][17] ),
    .B2(_07234_),
    .X(_05230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09459_ (.A(_06968_),
    .X(_07242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09460_ (.A1_N(_07242_),
    .A2_N(_07232_),
    .B1(\design_top.MEM[15][16] ),
    .B2(_07234_),
    .X(_05229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09461_ (.A(_06892_),
    .X(_07243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09462_ (.A(_07205_),
    .B(_07218_),
    .X(_07244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09463_ (.A(_07244_),
    .X(_07245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09464_ (.A(_07048_),
    .X(_07246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09465_ (.A1(_07246_),
    .A2(_07221_),
    .B1(_07244_),
    .X(_07247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09466_ (.A(_07247_),
    .X(_07248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09467_ (.A1_N(_07243_),
    .A2_N(_07245_),
    .B1(\design_top.MEM[15][31] ),
    .B2(_07248_),
    .X(_05228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09468_ (.A1_N(_07210_),
    .A2_N(_07245_),
    .B1(\design_top.MEM[15][30] ),
    .B2(_07248_),
    .X(_05227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09469_ (.A1_N(_07211_),
    .A2_N(_07245_),
    .B1(\design_top.MEM[15][29] ),
    .B2(_07248_),
    .X(_05226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09470_ (.A1_N(_07212_),
    .A2_N(_07245_),
    .B1(\design_top.MEM[15][28] ),
    .B2(_07248_),
    .X(_05225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09471_ (.A1_N(_07213_),
    .A2_N(_07245_),
    .B1(\design_top.MEM[15][27] ),
    .B2(_07248_),
    .X(_05224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09472_ (.A1_N(_07214_),
    .A2_N(_07244_),
    .B1(\design_top.MEM[15][26] ),
    .B2(_07247_),
    .X(_05223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09473_ (.A1_N(_07215_),
    .A2_N(_07244_),
    .B1(\design_top.MEM[15][25] ),
    .B2(_07247_),
    .X(_05222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09474_ (.A1_N(_07216_),
    .A2_N(_07244_),
    .B1(\design_top.MEM[15][24] ),
    .B2(_07247_),
    .X(_05221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09475_ (.A(_02480_),
    .B(_01337_),
    .X(_07249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09476_ (.A(_01371_),
    .B(_07249_),
    .X(_07250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09477_ (.A(_06985_),
    .B(_07250_),
    .X(_07251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09478_ (.A(_07193_),
    .B(_07251_),
    .X(_07252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09479_ (.A(_07252_),
    .X(_07253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _09480_ (.A(_07064_),
    .B(wbs_adr_i[1]),
    .C(wbs_adr_i[0]),
    .X(_07254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09481_ (.A(_07254_),
    .X(_07255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09482_ (.A(_07255_),
    .X(_07256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09483_ (.A1(_07151_),
    .A2(_07256_),
    .B1(_07252_),
    .X(_07257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09484_ (.A(_07257_),
    .X(_07258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09485_ (.A1_N(_07217_),
    .A2_N(_07253_),
    .B1(\design_top.MEM[16][15] ),
    .B2(_07258_),
    .X(_05220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09486_ (.A1_N(_07224_),
    .A2_N(_07253_),
    .B1(\design_top.MEM[16][14] ),
    .B2(_07258_),
    .X(_05219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09487_ (.A1_N(_07225_),
    .A2_N(_07253_),
    .B1(\design_top.MEM[16][13] ),
    .B2(_07258_),
    .X(_05218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09488_ (.A1_N(_07226_),
    .A2_N(_07253_),
    .B1(\design_top.MEM[16][12] ),
    .B2(_07258_),
    .X(_05217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09489_ (.A1_N(_07227_),
    .A2_N(_07253_),
    .B1(\design_top.MEM[16][11] ),
    .B2(_07258_),
    .X(_05216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09490_ (.A1_N(_07228_),
    .A2_N(_07252_),
    .B1(\design_top.MEM[16][10] ),
    .B2(_07257_),
    .X(_05215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09491_ (.A1_N(_07229_),
    .A2_N(_07252_),
    .B1(\design_top.MEM[16][9] ),
    .B2(_07257_),
    .X(_05214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09492_ (.A1_N(_07230_),
    .A2_N(_07252_),
    .B1(\design_top.MEM[16][8] ),
    .B2(_07257_),
    .X(_05213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09493_ (.A(_07205_),
    .B(_07251_),
    .X(_07259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09494_ (.A(_07259_),
    .X(_07260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09495_ (.A1(_07151_),
    .A2(_07256_),
    .B1(_07259_),
    .X(_07261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09496_ (.A(_07261_),
    .X(_07262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09497_ (.A1_N(_07243_),
    .A2_N(_07260_),
    .B1(\design_top.MEM[16][31] ),
    .B2(_07262_),
    .X(_05212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09498_ (.A1_N(_07210_),
    .A2_N(_07260_),
    .B1(\design_top.MEM[16][30] ),
    .B2(_07262_),
    .X(_05211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09499_ (.A1_N(_07211_),
    .A2_N(_07260_),
    .B1(\design_top.MEM[16][29] ),
    .B2(_07262_),
    .X(_05210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09500_ (.A1_N(_07212_),
    .A2_N(_07260_),
    .B1(\design_top.MEM[16][28] ),
    .B2(_07262_),
    .X(_05209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09501_ (.A1_N(_07213_),
    .A2_N(_07260_),
    .B1(\design_top.MEM[16][27] ),
    .B2(_07262_),
    .X(_05208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09502_ (.A1_N(_07214_),
    .A2_N(_07259_),
    .B1(\design_top.MEM[16][26] ),
    .B2(_07261_),
    .X(_05207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09503_ (.A1_N(_07215_),
    .A2_N(_07259_),
    .B1(\design_top.MEM[16][25] ),
    .B2(_07261_),
    .X(_05206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09504_ (.A1_N(_07216_),
    .A2_N(_07259_),
    .B1(\design_top.MEM[16][24] ),
    .B2(_07261_),
    .X(_05205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09505_ (.A(_07200_),
    .B(_07251_),
    .X(_07263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09506_ (.A(_07263_),
    .X(_07264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09507_ (.A1(_07151_),
    .A2(_07256_),
    .B1(_07263_),
    .X(_07265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09508_ (.A(_07265_),
    .X(_07266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09509_ (.A1_N(_07231_),
    .A2_N(_07264_),
    .B1(\design_top.MEM[16][23] ),
    .B2(_07266_),
    .X(_05204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09510_ (.A1_N(_07236_),
    .A2_N(_07264_),
    .B1(\design_top.MEM[16][22] ),
    .B2(_07266_),
    .X(_05203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09511_ (.A1_N(_07237_),
    .A2_N(_07264_),
    .B1(\design_top.MEM[16][21] ),
    .B2(_07266_),
    .X(_05202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09512_ (.A1_N(_07238_),
    .A2_N(_07264_),
    .B1(\design_top.MEM[16][20] ),
    .B2(_07266_),
    .X(_05201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09513_ (.A1_N(_07239_),
    .A2_N(_07264_),
    .B1(\design_top.MEM[16][19] ),
    .B2(_07266_),
    .X(_05200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09514_ (.A1_N(_07240_),
    .A2_N(_07263_),
    .B1(\design_top.MEM[16][18] ),
    .B2(_07265_),
    .X(_05199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09515_ (.A1_N(_07241_),
    .A2_N(_07263_),
    .B1(\design_top.MEM[16][17] ),
    .B2(_07265_),
    .X(_05198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09516_ (.A1_N(_07242_),
    .A2_N(_07263_),
    .B1(\design_top.MEM[16][16] ),
    .B2(_07265_),
    .X(_05197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09517_ (.A(_07154_),
    .B(_07250_),
    .X(_07267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09518_ (.A(_07193_),
    .B(_07267_),
    .X(_07268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09519_ (.A(_07268_),
    .X(_07269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09520_ (.A1(_07190_),
    .A2(_07256_),
    .B1(_07268_),
    .X(_07270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09521_ (.A(_07270_),
    .X(_07271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09522_ (.A1_N(_07217_),
    .A2_N(_07269_),
    .B1(\design_top.MEM[17][15] ),
    .B2(_07271_),
    .X(_05196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09523_ (.A1_N(_07224_),
    .A2_N(_07269_),
    .B1(\design_top.MEM[17][14] ),
    .B2(_07271_),
    .X(_05195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09524_ (.A1_N(_07225_),
    .A2_N(_07269_),
    .B1(\design_top.MEM[17][13] ),
    .B2(_07271_),
    .X(_05194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09525_ (.A1_N(_07226_),
    .A2_N(_07269_),
    .B1(\design_top.MEM[17][12] ),
    .B2(_07271_),
    .X(_05193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09526_ (.A1_N(_07227_),
    .A2_N(_07269_),
    .B1(\design_top.MEM[17][11] ),
    .B2(_07271_),
    .X(_05192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09527_ (.A1_N(_07228_),
    .A2_N(_07268_),
    .B1(\design_top.MEM[17][10] ),
    .B2(_07270_),
    .X(_05191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09528_ (.A1_N(_07229_),
    .A2_N(_07268_),
    .B1(\design_top.MEM[17][9] ),
    .B2(_07270_),
    .X(_05190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09529_ (.A1_N(_07230_),
    .A2_N(_07268_),
    .B1(\design_top.MEM[17][8] ),
    .B2(_07270_),
    .X(_05189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09530_ (.A(_07200_),
    .B(_07267_),
    .X(_07272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09531_ (.A(_07272_),
    .X(_07273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09532_ (.A1(_07190_),
    .A2(_07256_),
    .B1(_07272_),
    .X(_07274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09533_ (.A(_07274_),
    .X(_07275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09534_ (.A1_N(_07231_),
    .A2_N(_07273_),
    .B1(\design_top.MEM[17][23] ),
    .B2(_07275_),
    .X(_05188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09535_ (.A1_N(_07236_),
    .A2_N(_07273_),
    .B1(\design_top.MEM[17][22] ),
    .B2(_07275_),
    .X(_05187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09536_ (.A1_N(_07237_),
    .A2_N(_07273_),
    .B1(\design_top.MEM[17][21] ),
    .B2(_07275_),
    .X(_05186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09537_ (.A1_N(_07238_),
    .A2_N(_07273_),
    .B1(\design_top.MEM[17][20] ),
    .B2(_07275_),
    .X(_05185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09538_ (.A1_N(_07239_),
    .A2_N(_07273_),
    .B1(\design_top.MEM[17][19] ),
    .B2(_07275_),
    .X(_05184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09539_ (.A1_N(_07240_),
    .A2_N(_07272_),
    .B1(\design_top.MEM[17][18] ),
    .B2(_07274_),
    .X(_05183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09540_ (.A1_N(_07241_),
    .A2_N(_07272_),
    .B1(\design_top.MEM[17][17] ),
    .B2(_07274_),
    .X(_05182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09541_ (.A1_N(_07242_),
    .A2_N(_07272_),
    .B1(\design_top.MEM[17][16] ),
    .B2(_07274_),
    .X(_05181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09542_ (.A(_07205_),
    .B(_07267_),
    .X(_07276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09543_ (.A(_07276_),
    .X(_07277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09544_ (.A(_07255_),
    .X(_07278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09545_ (.A1(_07190_),
    .A2(_07278_),
    .B1(_07276_),
    .X(_07279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09546_ (.A(_07279_),
    .X(_07280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09547_ (.A1_N(_07243_),
    .A2_N(_07277_),
    .B1(\design_top.MEM[17][31] ),
    .B2(_07280_),
    .X(_05180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09548_ (.A1_N(_07210_),
    .A2_N(_07277_),
    .B1(\design_top.MEM[17][30] ),
    .B2(_07280_),
    .X(_05179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09549_ (.A1_N(_07211_),
    .A2_N(_07277_),
    .B1(\design_top.MEM[17][29] ),
    .B2(_07280_),
    .X(_05178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09550_ (.A1_N(_07212_),
    .A2_N(_07277_),
    .B1(\design_top.MEM[17][28] ),
    .B2(_07280_),
    .X(_05177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09551_ (.A1_N(_07213_),
    .A2_N(_07277_),
    .B1(\design_top.MEM[17][27] ),
    .B2(_07280_),
    .X(_05176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09552_ (.A1_N(_07214_),
    .A2_N(_07276_),
    .B1(\design_top.MEM[17][26] ),
    .B2(_07279_),
    .X(_05175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09553_ (.A1_N(_07215_),
    .A2_N(_07276_),
    .B1(\design_top.MEM[17][25] ),
    .B2(_07279_),
    .X(_05174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09554_ (.A1_N(_07216_),
    .A2_N(_07276_),
    .B1(\design_top.MEM[17][24] ),
    .B2(_07279_),
    .X(_05173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09555_ (.A(_06970_),
    .B(_07250_),
    .X(_07281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09556_ (.A(_07193_),
    .B(_07281_),
    .X(_07282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09557_ (.A(_07282_),
    .X(_07283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09558_ (.A1(_07197_),
    .A2(_07278_),
    .B1(_07282_),
    .X(_07284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09559_ (.A(_07284_),
    .X(_07285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09560_ (.A1_N(_07217_),
    .A2_N(_07283_),
    .B1(\design_top.MEM[18][15] ),
    .B2(_07285_),
    .X(_05172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09561_ (.A1_N(_07224_),
    .A2_N(_07283_),
    .B1(\design_top.MEM[18][14] ),
    .B2(_07285_),
    .X(_05171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09562_ (.A1_N(_07225_),
    .A2_N(_07283_),
    .B1(\design_top.MEM[18][13] ),
    .B2(_07285_),
    .X(_05170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09563_ (.A1_N(_07226_),
    .A2_N(_07283_),
    .B1(\design_top.MEM[18][12] ),
    .B2(_07285_),
    .X(_05169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09564_ (.A1_N(_07227_),
    .A2_N(_07283_),
    .B1(\design_top.MEM[18][11] ),
    .B2(_07285_),
    .X(_05168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09565_ (.A1_N(_07228_),
    .A2_N(_07282_),
    .B1(\design_top.MEM[18][10] ),
    .B2(_07284_),
    .X(_05167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09566_ (.A1_N(_07229_),
    .A2_N(_07282_),
    .B1(\design_top.MEM[18][9] ),
    .B2(_07284_),
    .X(_05166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09567_ (.A1_N(_07230_),
    .A2_N(_07282_),
    .B1(\design_top.MEM[18][8] ),
    .B2(_07284_),
    .X(_05165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09568_ (.A(_07200_),
    .B(_07281_),
    .X(_07286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09569_ (.A(_07286_),
    .X(_07287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09570_ (.A1(_07197_),
    .A2(_07278_),
    .B1(_07286_),
    .X(_07288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09571_ (.A(_07288_),
    .X(_07289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09572_ (.A1_N(_07231_),
    .A2_N(_07287_),
    .B1(\design_top.MEM[18][23] ),
    .B2(_07289_),
    .X(_05164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09573_ (.A1_N(_07236_),
    .A2_N(_07287_),
    .B1(\design_top.MEM[18][22] ),
    .B2(_07289_),
    .X(_05163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09574_ (.A1_N(_07237_),
    .A2_N(_07287_),
    .B1(\design_top.MEM[18][21] ),
    .B2(_07289_),
    .X(_05162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09575_ (.A1_N(_07238_),
    .A2_N(_07287_),
    .B1(\design_top.MEM[18][20] ),
    .B2(_07289_),
    .X(_05161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09576_ (.A1_N(_07239_),
    .A2_N(_07287_),
    .B1(\design_top.MEM[18][19] ),
    .B2(_07289_),
    .X(_05160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09577_ (.A1_N(_07240_),
    .A2_N(_07286_),
    .B1(\design_top.MEM[18][18] ),
    .B2(_07288_),
    .X(_05159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09578_ (.A1_N(_07241_),
    .A2_N(_07286_),
    .B1(\design_top.MEM[18][17] ),
    .B2(_07288_),
    .X(_05158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09579_ (.A1_N(_07242_),
    .A2_N(_07286_),
    .B1(\design_top.MEM[18][16] ),
    .B2(_07288_),
    .X(_05157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09580_ (.A(_07205_),
    .B(_07281_),
    .X(_07290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09581_ (.A(_07290_),
    .X(_07291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09582_ (.A(_06977_),
    .X(_07292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09583_ (.A1(_07292_),
    .A2(_07278_),
    .B1(_07290_),
    .X(_07293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09584_ (.A(_07293_),
    .X(_07294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09585_ (.A1_N(_07243_),
    .A2_N(_07291_),
    .B1(\design_top.MEM[18][31] ),
    .B2(_07294_),
    .X(_05156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09586_ (.A1_N(_07210_),
    .A2_N(_07291_),
    .B1(\design_top.MEM[18][30] ),
    .B2(_07294_),
    .X(_05155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09587_ (.A1_N(_07211_),
    .A2_N(_07291_),
    .B1(\design_top.MEM[18][29] ),
    .B2(_07294_),
    .X(_05154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09588_ (.A1_N(_07212_),
    .A2_N(_07291_),
    .B1(\design_top.MEM[18][28] ),
    .B2(_07294_),
    .X(_05153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09589_ (.A1_N(_07213_),
    .A2_N(_07291_),
    .B1(\design_top.MEM[18][27] ),
    .B2(_07294_),
    .X(_05152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09590_ (.A1_N(_07214_),
    .A2_N(_07290_),
    .B1(\design_top.MEM[18][26] ),
    .B2(_07293_),
    .X(_05151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09591_ (.A1_N(_07215_),
    .A2_N(_07290_),
    .B1(\design_top.MEM[18][25] ),
    .B2(_07293_),
    .X(_05150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09592_ (.A1_N(_07216_),
    .A2_N(_07290_),
    .B1(\design_top.MEM[18][24] ),
    .B2(_07293_),
    .X(_05149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09593_ (.A(_06911_),
    .X(_07295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09594_ (.A(_07043_),
    .B(_07250_),
    .X(_07296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09595_ (.A(_07295_),
    .B(_07296_),
    .X(_07297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09596_ (.A(_07297_),
    .X(_07298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09597_ (.A1(_07246_),
    .A2(_07278_),
    .B1(_07297_),
    .X(_07299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09598_ (.A(_07299_),
    .X(_07300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09599_ (.A1_N(_07217_),
    .A2_N(_07298_),
    .B1(\design_top.MEM[19][15] ),
    .B2(_07300_),
    .X(_05148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09600_ (.A1_N(_07224_),
    .A2_N(_07298_),
    .B1(\design_top.MEM[19][14] ),
    .B2(_07300_),
    .X(_05147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09601_ (.A1_N(_07225_),
    .A2_N(_07298_),
    .B1(\design_top.MEM[19][13] ),
    .B2(_07300_),
    .X(_05146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09602_ (.A1_N(_07226_),
    .A2_N(_07298_),
    .B1(\design_top.MEM[19][12] ),
    .B2(_07300_),
    .X(_05145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09603_ (.A1_N(_07227_),
    .A2_N(_07298_),
    .B1(\design_top.MEM[19][11] ),
    .B2(_07300_),
    .X(_05144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09604_ (.A1_N(_07228_),
    .A2_N(_07297_),
    .B1(\design_top.MEM[19][10] ),
    .B2(_07299_),
    .X(_05143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09605_ (.A1_N(_07229_),
    .A2_N(_07297_),
    .B1(\design_top.MEM[19][9] ),
    .B2(_07299_),
    .X(_05142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09606_ (.A1_N(_07230_),
    .A2_N(_07297_),
    .B1(\design_top.MEM[19][8] ),
    .B2(_07299_),
    .X(_05141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09607_ (.A(_06942_),
    .X(_07301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09608_ (.A(_07301_),
    .B(_07296_),
    .X(_07302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09609_ (.A(_07302_),
    .X(_07303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09610_ (.A1(_07246_),
    .A2(_07255_),
    .B1(_07302_),
    .X(_07304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09611_ (.A(_07304_),
    .X(_07305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09612_ (.A1_N(_07231_),
    .A2_N(_07303_),
    .B1(\design_top.MEM[19][23] ),
    .B2(_07305_),
    .X(_05140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09613_ (.A1_N(_07236_),
    .A2_N(_07303_),
    .B1(\design_top.MEM[19][22] ),
    .B2(_07305_),
    .X(_05139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09614_ (.A1_N(_07237_),
    .A2_N(_07303_),
    .B1(\design_top.MEM[19][21] ),
    .B2(_07305_),
    .X(_05138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09615_ (.A1_N(_07238_),
    .A2_N(_07303_),
    .B1(\design_top.MEM[19][20] ),
    .B2(_07305_),
    .X(_05137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09616_ (.A1_N(_07239_),
    .A2_N(_07303_),
    .B1(\design_top.MEM[19][19] ),
    .B2(_07305_),
    .X(_05136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09617_ (.A1_N(_07240_),
    .A2_N(_07302_),
    .B1(\design_top.MEM[19][18] ),
    .B2(_07304_),
    .X(_05135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09618_ (.A1_N(_07241_),
    .A2_N(_07302_),
    .B1(\design_top.MEM[19][17] ),
    .B2(_07304_),
    .X(_05134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09619_ (.A1_N(_07242_),
    .A2_N(_07302_),
    .B1(\design_top.MEM[19][16] ),
    .B2(_07304_),
    .X(_05133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09620_ (.A(_06844_),
    .X(_07306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09621_ (.A(_07306_),
    .B(_07296_),
    .X(_07307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09622_ (.A(_07307_),
    .X(_07308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09623_ (.A1(_07246_),
    .A2(_07255_),
    .B1(_07307_),
    .X(_07309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09624_ (.A(_07309_),
    .X(_07310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09625_ (.A1_N(_07243_),
    .A2_N(_07308_),
    .B1(\design_top.MEM[19][31] ),
    .B2(_07310_),
    .X(_05132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09626_ (.A(_06655_),
    .X(_07311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09627_ (.A1_N(_07311_),
    .A2_N(_07308_),
    .B1(\design_top.MEM[19][30] ),
    .B2(_07310_),
    .X(_05131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09628_ (.A(_06873_),
    .X(_07312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09629_ (.A1_N(_07312_),
    .A2_N(_07308_),
    .B1(\design_top.MEM[19][29] ),
    .B2(_07310_),
    .X(_05130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09630_ (.A(_06876_),
    .X(_07313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09631_ (.A1_N(_07313_),
    .A2_N(_07308_),
    .B1(\design_top.MEM[19][28] ),
    .B2(_07310_),
    .X(_05129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09632_ (.A(_06879_),
    .X(_07314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09633_ (.A1_N(_07314_),
    .A2_N(_07308_),
    .B1(\design_top.MEM[19][27] ),
    .B2(_07310_),
    .X(_05128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09634_ (.A(_06882_),
    .X(_07315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09635_ (.A1_N(_07315_),
    .A2_N(_07307_),
    .B1(\design_top.MEM[19][26] ),
    .B2(_07309_),
    .X(_05127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09636_ (.A(_06885_),
    .X(_07316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09637_ (.A1_N(_07316_),
    .A2_N(_07307_),
    .B1(\design_top.MEM[19][25] ),
    .B2(_07309_),
    .X(_05126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09638_ (.A(_06888_),
    .X(_07317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09639_ (.A1_N(_07317_),
    .A2_N(_07307_),
    .B1(\design_top.MEM[19][24] ),
    .B2(_07309_),
    .X(_05125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09640_ (.A(_06908_),
    .X(_07318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09641_ (.A(_07154_),
    .B(_06896_),
    .X(_07319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09642_ (.A(_07295_),
    .B(_07319_),
    .X(_07320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09643_ (.A(_07320_),
    .X(_07321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09644_ (.A1(_07190_),
    .A2(_06905_),
    .B1(_07320_),
    .X(_07322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09645_ (.A(_07322_),
    .X(_07323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09646_ (.A1_N(_07318_),
    .A2_N(_07321_),
    .B1(\design_top.MEM[1][15] ),
    .B2(_07323_),
    .X(_05124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09647_ (.A(_06918_),
    .X(_07324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09648_ (.A1_N(_07324_),
    .A2_N(_07321_),
    .B1(\design_top.MEM[1][14] ),
    .B2(_07323_),
    .X(_05123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09649_ (.A(_06921_),
    .X(_07325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09650_ (.A1_N(_07325_),
    .A2_N(_07321_),
    .B1(\design_top.MEM[1][13] ),
    .B2(_07323_),
    .X(_05122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09651_ (.A(_06924_),
    .X(_07326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09652_ (.A1_N(_07326_),
    .A2_N(_07321_),
    .B1(\design_top.MEM[1][12] ),
    .B2(_07323_),
    .X(_05121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09653_ (.A(_06927_),
    .X(_07327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09654_ (.A1_N(_07327_),
    .A2_N(_07321_),
    .B1(\design_top.MEM[1][11] ),
    .B2(_07323_),
    .X(_05120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09655_ (.A(_06930_),
    .X(_07328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09656_ (.A1_N(_07328_),
    .A2_N(_07320_),
    .B1(\design_top.MEM[1][10] ),
    .B2(_07322_),
    .X(_05119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09657_ (.A(_06933_),
    .X(_07329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09658_ (.A1_N(_07329_),
    .A2_N(_07320_),
    .B1(\design_top.MEM[1][9] ),
    .B2(_07322_),
    .X(_05118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09659_ (.A(_06936_),
    .X(_07330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09660_ (.A1_N(_07330_),
    .A2_N(_07320_),
    .B1(\design_top.MEM[1][8] ),
    .B2(_07322_),
    .X(_05117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09661_ (.A(_06939_),
    .X(_07331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09662_ (.A(_07301_),
    .B(_07319_),
    .X(_07332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09663_ (.A(_07332_),
    .X(_07333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09664_ (.A(_07189_),
    .X(_07334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09665_ (.A1(_07334_),
    .A2(_06904_),
    .B1(_07332_),
    .X(_07335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09666_ (.A(_07335_),
    .X(_07336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09667_ (.A1_N(_07331_),
    .A2_N(_07333_),
    .B1(\design_top.MEM[1][23] ),
    .B2(_07336_),
    .X(_05116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09668_ (.A(_06949_),
    .X(_07337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09669_ (.A1_N(_07337_),
    .A2_N(_07333_),
    .B1(\design_top.MEM[1][22] ),
    .B2(_07336_),
    .X(_05115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09670_ (.A(_06952_),
    .X(_07338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09671_ (.A1_N(_07338_),
    .A2_N(_07333_),
    .B1(\design_top.MEM[1][21] ),
    .B2(_07336_),
    .X(_05114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09672_ (.A(_06955_),
    .X(_07339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09673_ (.A1_N(_07339_),
    .A2_N(_07333_),
    .B1(\design_top.MEM[1][20] ),
    .B2(_07336_),
    .X(_05113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09674_ (.A(_06958_),
    .X(_07340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09675_ (.A1_N(_07340_),
    .A2_N(_07333_),
    .B1(\design_top.MEM[1][19] ),
    .B2(_07336_),
    .X(_05112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09676_ (.A(_06961_),
    .X(_07341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09677_ (.A1_N(_07341_),
    .A2_N(_07332_),
    .B1(\design_top.MEM[1][18] ),
    .B2(_07335_),
    .X(_05111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09678_ (.A(_06964_),
    .X(_07342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09679_ (.A1_N(_07342_),
    .A2_N(_07332_),
    .B1(\design_top.MEM[1][17] ),
    .B2(_07335_),
    .X(_05110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09680_ (.A(_06967_),
    .X(_07343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09681_ (.A1_N(_07343_),
    .A2_N(_07332_),
    .B1(\design_top.MEM[1][16] ),
    .B2(_07335_),
    .X(_05109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09682_ (.A(_06891_),
    .X(_07344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09683_ (.A(_07306_),
    .B(_07319_),
    .X(_07345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09684_ (.A(_07345_),
    .X(_07346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09685_ (.A1(_07334_),
    .A2(_06904_),
    .B1(_07345_),
    .X(_07347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09686_ (.A(_07347_),
    .X(_07348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09687_ (.A1_N(_07344_),
    .A2_N(_07346_),
    .B1(\design_top.MEM[1][31] ),
    .B2(_07348_),
    .X(_05108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09688_ (.A1_N(_07311_),
    .A2_N(_07346_),
    .B1(\design_top.MEM[1][30] ),
    .B2(_07348_),
    .X(_05107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09689_ (.A1_N(_07312_),
    .A2_N(_07346_),
    .B1(\design_top.MEM[1][29] ),
    .B2(_07348_),
    .X(_05106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09690_ (.A1_N(_07313_),
    .A2_N(_07346_),
    .B1(\design_top.MEM[1][28] ),
    .B2(_07348_),
    .X(_05105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09691_ (.A1_N(_07314_),
    .A2_N(_07346_),
    .B1(\design_top.MEM[1][27] ),
    .B2(_07348_),
    .X(_05104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09692_ (.A1_N(_07315_),
    .A2_N(_07345_),
    .B1(\design_top.MEM[1][26] ),
    .B2(_07347_),
    .X(_05103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09693_ (.A1_N(_07316_),
    .A2_N(_07345_),
    .B1(\design_top.MEM[1][25] ),
    .B2(_07347_),
    .X(_05102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09694_ (.A1_N(_07317_),
    .A2_N(_07345_),
    .B1(\design_top.MEM[1][24] ),
    .B2(_07347_),
    .X(_05101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09695_ (.A(_07306_),
    .B(_07169_),
    .X(_07349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09696_ (.A(_07349_),
    .X(_07350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09697_ (.A1(_07292_),
    .A2(_07166_),
    .B1(_07349_),
    .X(_07351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09698_ (.A(_07351_),
    .X(_07352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09699_ (.A1_N(_07344_),
    .A2_N(_07350_),
    .B1(\design_top.MEM[6][31] ),
    .B2(_07352_),
    .X(_05100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09700_ (.A1_N(_07311_),
    .A2_N(_07350_),
    .B1(\design_top.MEM[6][30] ),
    .B2(_07352_),
    .X(_05099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09701_ (.A1_N(_07312_),
    .A2_N(_07350_),
    .B1(\design_top.MEM[6][29] ),
    .B2(_07352_),
    .X(_05098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09702_ (.A1_N(_07313_),
    .A2_N(_07350_),
    .B1(\design_top.MEM[6][28] ),
    .B2(_07352_),
    .X(_05097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09703_ (.A1_N(_07314_),
    .A2_N(_07350_),
    .B1(\design_top.MEM[6][27] ),
    .B2(_07352_),
    .X(_05096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09704_ (.A1_N(_07315_),
    .A2_N(_07349_),
    .B1(\design_top.MEM[6][26] ),
    .B2(_07351_),
    .X(_05095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09705_ (.A1_N(_07316_),
    .A2_N(_07349_),
    .B1(\design_top.MEM[6][25] ),
    .B2(_07351_),
    .X(_05094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09706_ (.A1_N(_07317_),
    .A2_N(_07349_),
    .B1(\design_top.MEM[6][24] ),
    .B2(_07351_),
    .X(_05093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09707_ (.A(_07042_),
    .B(_07127_),
    .X(_07353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09708_ (.A(_07295_),
    .B(_07353_),
    .X(_07354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09709_ (.A(_07354_),
    .X(_07355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09710_ (.A1(_07246_),
    .A2(_07166_),
    .B1(_07354_),
    .X(_07356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09711_ (.A(_07356_),
    .X(_07357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09712_ (.A1_N(_07318_),
    .A2_N(_07355_),
    .B1(\design_top.MEM[7][15] ),
    .B2(_07357_),
    .X(_05092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09713_ (.A1_N(_07324_),
    .A2_N(_07355_),
    .B1(\design_top.MEM[7][14] ),
    .B2(_07357_),
    .X(_05091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09714_ (.A1_N(_07325_),
    .A2_N(_07355_),
    .B1(\design_top.MEM[7][13] ),
    .B2(_07357_),
    .X(_05090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09715_ (.A1_N(_07326_),
    .A2_N(_07355_),
    .B1(\design_top.MEM[7][12] ),
    .B2(_07357_),
    .X(_05089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09716_ (.A1_N(_07327_),
    .A2_N(_07355_),
    .B1(\design_top.MEM[7][11] ),
    .B2(_07357_),
    .X(_05088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09717_ (.A1_N(_07328_),
    .A2_N(_07354_),
    .B1(\design_top.MEM[7][10] ),
    .B2(_07356_),
    .X(_05087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09718_ (.A1_N(_07329_),
    .A2_N(_07354_),
    .B1(\design_top.MEM[7][9] ),
    .B2(_07356_),
    .X(_05086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09719_ (.A1_N(_07330_),
    .A2_N(_07354_),
    .B1(\design_top.MEM[7][8] ),
    .B2(_07356_),
    .X(_05085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09720_ (.A(_07306_),
    .B(_07353_),
    .X(_07358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09721_ (.A(_07358_),
    .X(_07359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09722_ (.A(_07048_),
    .X(_07360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09723_ (.A1(_07360_),
    .A2(_07132_),
    .B1(_07358_),
    .X(_07361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09724_ (.A(_07361_),
    .X(_07362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09725_ (.A1_N(_07344_),
    .A2_N(_07359_),
    .B1(\design_top.MEM[7][31] ),
    .B2(_07362_),
    .X(_05084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09726_ (.A1_N(_07311_),
    .A2_N(_07359_),
    .B1(\design_top.MEM[7][30] ),
    .B2(_07362_),
    .X(_05083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09727_ (.A1_N(_07312_),
    .A2_N(_07359_),
    .B1(\design_top.MEM[7][29] ),
    .B2(_07362_),
    .X(_05082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09728_ (.A1_N(_07313_),
    .A2_N(_07359_),
    .B1(\design_top.MEM[7][28] ),
    .B2(_07362_),
    .X(_05081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09729_ (.A1_N(_07314_),
    .A2_N(_07359_),
    .B1(\design_top.MEM[7][27] ),
    .B2(_07362_),
    .X(_05080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09730_ (.A1_N(_07315_),
    .A2_N(_07358_),
    .B1(\design_top.MEM[7][26] ),
    .B2(_07361_),
    .X(_05079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09731_ (.A1_N(_07316_),
    .A2_N(_07358_),
    .B1(\design_top.MEM[7][25] ),
    .B2(_07361_),
    .X(_05078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09732_ (.A1_N(_07317_),
    .A2_N(_07358_),
    .B1(\design_top.MEM[7][24] ),
    .B2(_07361_),
    .X(_05077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09733_ (.A(_01333_),
    .B(_07249_),
    .X(_07363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09734_ (.A(_06985_),
    .B(_07363_),
    .X(_07364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09735_ (.A(_07295_),
    .B(_07364_),
    .X(_07365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09736_ (.A(_07365_),
    .X(_07366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _09737_ (.A(_07064_),
    .B(wbs_adr_i[1]),
    .C(_07065_),
    .X(_07367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09738_ (.A(_07367_),
    .X(_07368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09739_ (.A(_07368_),
    .X(_07369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09740_ (.A1(_07151_),
    .A2(_07369_),
    .B1(_07365_),
    .X(_07370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09741_ (.A(_07370_),
    .X(_07371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09742_ (.A1_N(_07318_),
    .A2_N(_07366_),
    .B1(\design_top.MEM[20][15] ),
    .B2(_07371_),
    .X(_05076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09743_ (.A1_N(_07324_),
    .A2_N(_07366_),
    .B1(\design_top.MEM[20][14] ),
    .B2(_07371_),
    .X(_05075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09744_ (.A1_N(_07325_),
    .A2_N(_07366_),
    .B1(\design_top.MEM[20][13] ),
    .B2(_07371_),
    .X(_05074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09745_ (.A1_N(_07326_),
    .A2_N(_07366_),
    .B1(\design_top.MEM[20][12] ),
    .B2(_07371_),
    .X(_05073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09746_ (.A1_N(_07327_),
    .A2_N(_07366_),
    .B1(\design_top.MEM[20][11] ),
    .B2(_07371_),
    .X(_05072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09747_ (.A1_N(_07328_),
    .A2_N(_07365_),
    .B1(\design_top.MEM[20][10] ),
    .B2(_07370_),
    .X(_05071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09748_ (.A1_N(_07329_),
    .A2_N(_07365_),
    .B1(\design_top.MEM[20][9] ),
    .B2(_07370_),
    .X(_05070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09749_ (.A1_N(_07330_),
    .A2_N(_07365_),
    .B1(\design_top.MEM[20][8] ),
    .B2(_07370_),
    .X(_05069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09750_ (.A(_07301_),
    .B(_07364_),
    .X(_07372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09751_ (.A(_07372_),
    .X(_07373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09752_ (.A(_07150_),
    .X(_07374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09753_ (.A1(_07374_),
    .A2(_07369_),
    .B1(_07372_),
    .X(_07375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09754_ (.A(_07375_),
    .X(_07376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09755_ (.A1_N(_07331_),
    .A2_N(_07373_),
    .B1(\design_top.MEM[20][23] ),
    .B2(_07376_),
    .X(_05068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09756_ (.A1_N(_07337_),
    .A2_N(_07373_),
    .B1(\design_top.MEM[20][22] ),
    .B2(_07376_),
    .X(_05067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09757_ (.A1_N(_07338_),
    .A2_N(_07373_),
    .B1(\design_top.MEM[20][21] ),
    .B2(_07376_),
    .X(_05066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09758_ (.A1_N(_07339_),
    .A2_N(_07373_),
    .B1(\design_top.MEM[20][20] ),
    .B2(_07376_),
    .X(_05065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09759_ (.A1_N(_07340_),
    .A2_N(_07373_),
    .B1(\design_top.MEM[20][19] ),
    .B2(_07376_),
    .X(_05064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09760_ (.A1_N(_07341_),
    .A2_N(_07372_),
    .B1(\design_top.MEM[20][18] ),
    .B2(_07375_),
    .X(_05063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09761_ (.A1_N(_07342_),
    .A2_N(_07372_),
    .B1(\design_top.MEM[20][17] ),
    .B2(_07375_),
    .X(_05062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09762_ (.A1_N(_07343_),
    .A2_N(_07372_),
    .B1(\design_top.MEM[20][16] ),
    .B2(_07375_),
    .X(_05061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09763_ (.A(_07306_),
    .B(_07364_),
    .X(_07377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09764_ (.A(_07377_),
    .X(_07378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09765_ (.A1(_07374_),
    .A2(_07369_),
    .B1(_07377_),
    .X(_07379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09766_ (.A(_07379_),
    .X(_07380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09767_ (.A1_N(_07344_),
    .A2_N(_07378_),
    .B1(\design_top.MEM[20][31] ),
    .B2(_07380_),
    .X(_05060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09768_ (.A1_N(_07311_),
    .A2_N(_07378_),
    .B1(\design_top.MEM[20][30] ),
    .B2(_07380_),
    .X(_05059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09769_ (.A1_N(_07312_),
    .A2_N(_07378_),
    .B1(\design_top.MEM[20][29] ),
    .B2(_07380_),
    .X(_05058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09770_ (.A1_N(_07313_),
    .A2_N(_07378_),
    .B1(\design_top.MEM[20][28] ),
    .B2(_07380_),
    .X(_05057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09771_ (.A1_N(_07314_),
    .A2_N(_07378_),
    .B1(\design_top.MEM[20][27] ),
    .B2(_07380_),
    .X(_05056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09772_ (.A1_N(_07315_),
    .A2_N(_07377_),
    .B1(\design_top.MEM[20][26] ),
    .B2(_07379_),
    .X(_05055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09773_ (.A1_N(_07316_),
    .A2_N(_07377_),
    .B1(\design_top.MEM[20][25] ),
    .B2(_07379_),
    .X(_05054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09774_ (.A1_N(_07317_),
    .A2_N(_07377_),
    .B1(\design_top.MEM[20][24] ),
    .B2(_07379_),
    .X(_05053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09775_ (.A(_06851_),
    .B(_07363_),
    .X(_07381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09776_ (.A(_07295_),
    .B(_07381_),
    .X(_07382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09777_ (.A(_07382_),
    .X(_07383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09778_ (.A1(_07334_),
    .A2(_07369_),
    .B1(_07382_),
    .X(_07384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09779_ (.A(_07384_),
    .X(_07385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09780_ (.A1_N(_07318_),
    .A2_N(_07383_),
    .B1(\design_top.MEM[21][15] ),
    .B2(_07385_),
    .X(_05052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09781_ (.A1_N(_07324_),
    .A2_N(_07383_),
    .B1(\design_top.MEM[21][14] ),
    .B2(_07385_),
    .X(_05051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09782_ (.A1_N(_07325_),
    .A2_N(_07383_),
    .B1(\design_top.MEM[21][13] ),
    .B2(_07385_),
    .X(_05050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09783_ (.A1_N(_07326_),
    .A2_N(_07383_),
    .B1(\design_top.MEM[21][12] ),
    .B2(_07385_),
    .X(_05049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09784_ (.A1_N(_07327_),
    .A2_N(_07383_),
    .B1(\design_top.MEM[21][11] ),
    .B2(_07385_),
    .X(_05048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09785_ (.A1_N(_07328_),
    .A2_N(_07382_),
    .B1(\design_top.MEM[21][10] ),
    .B2(_07384_),
    .X(_05047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09786_ (.A1_N(_07329_),
    .A2_N(_07382_),
    .B1(\design_top.MEM[21][9] ),
    .B2(_07384_),
    .X(_05046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09787_ (.A1_N(_07330_),
    .A2_N(_07382_),
    .B1(\design_top.MEM[21][8] ),
    .B2(_07384_),
    .X(_05045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09788_ (.A(_07301_),
    .B(_07381_),
    .X(_07386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09789_ (.A(_07386_),
    .X(_07387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09790_ (.A1(_07334_),
    .A2(_07369_),
    .B1(_07386_),
    .X(_07388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09791_ (.A(_07388_),
    .X(_07389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09792_ (.A1_N(_07331_),
    .A2_N(_07387_),
    .B1(\design_top.MEM[21][23] ),
    .B2(_07389_),
    .X(_05044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09793_ (.A1_N(_07337_),
    .A2_N(_07387_),
    .B1(\design_top.MEM[21][22] ),
    .B2(_07389_),
    .X(_05043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09794_ (.A1_N(_07338_),
    .A2_N(_07387_),
    .B1(\design_top.MEM[21][21] ),
    .B2(_07389_),
    .X(_05042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09795_ (.A1_N(_07339_),
    .A2_N(_07387_),
    .B1(\design_top.MEM[21][20] ),
    .B2(_07389_),
    .X(_05041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09796_ (.A1_N(_07340_),
    .A2_N(_07387_),
    .B1(\design_top.MEM[21][19] ),
    .B2(_07389_),
    .X(_05040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09797_ (.A1_N(_07341_),
    .A2_N(_07386_),
    .B1(\design_top.MEM[21][18] ),
    .B2(_07388_),
    .X(_05039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09798_ (.A1_N(_07342_),
    .A2_N(_07386_),
    .B1(\design_top.MEM[21][17] ),
    .B2(_07388_),
    .X(_05038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09799_ (.A1_N(_07343_),
    .A2_N(_07386_),
    .B1(\design_top.MEM[21][16] ),
    .B2(_07388_),
    .X(_05037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09800_ (.A(_06844_),
    .X(_07390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09801_ (.A(_07390_),
    .B(_07381_),
    .X(_07391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09802_ (.A(_07391_),
    .X(_07392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09803_ (.A(_07368_),
    .X(_07393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09804_ (.A1(_07334_),
    .A2(_07393_),
    .B1(_07391_),
    .X(_07394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09805_ (.A(_07394_),
    .X(_07395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09806_ (.A1_N(_07344_),
    .A2_N(_07392_),
    .B1(\design_top.MEM[21][31] ),
    .B2(_07395_),
    .X(_05036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09807_ (.A(_06655_),
    .X(_07396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09808_ (.A1_N(_07396_),
    .A2_N(_07392_),
    .B1(\design_top.MEM[21][30] ),
    .B2(_07395_),
    .X(_05035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09809_ (.A(_06873_),
    .X(_07397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09810_ (.A1_N(_07397_),
    .A2_N(_07392_),
    .B1(\design_top.MEM[21][29] ),
    .B2(_07395_),
    .X(_05034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09811_ (.A(_06876_),
    .X(_07398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09812_ (.A1_N(_07398_),
    .A2_N(_07392_),
    .B1(\design_top.MEM[21][28] ),
    .B2(_07395_),
    .X(_05033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09813_ (.A(_06879_),
    .X(_07399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09814_ (.A1_N(_07399_),
    .A2_N(_07392_),
    .B1(\design_top.MEM[21][27] ),
    .B2(_07395_),
    .X(_05032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09815_ (.A(_06882_),
    .X(_07400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09816_ (.A1_N(_07400_),
    .A2_N(_07391_),
    .B1(\design_top.MEM[21][26] ),
    .B2(_07394_),
    .X(_05031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09817_ (.A(_06885_),
    .X(_07401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09818_ (.A1_N(_07401_),
    .A2_N(_07391_),
    .B1(\design_top.MEM[21][25] ),
    .B2(_07394_),
    .X(_05030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09819_ (.A(_06888_),
    .X(_07402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09820_ (.A1_N(_07402_),
    .A2_N(_07391_),
    .B1(\design_top.MEM[21][24] ),
    .B2(_07394_),
    .X(_05029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09821_ (.A(_06911_),
    .X(_07403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09822_ (.A(_06970_),
    .B(_07363_),
    .X(_07404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09823_ (.A(_07403_),
    .B(_07404_),
    .X(_07405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09824_ (.A(_07405_),
    .X(_07406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09825_ (.A1(_07292_),
    .A2(_07393_),
    .B1(_07405_),
    .X(_07407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09826_ (.A(_07407_),
    .X(_07408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09827_ (.A1_N(_07318_),
    .A2_N(_07406_),
    .B1(\design_top.MEM[22][15] ),
    .B2(_07408_),
    .X(_05028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09828_ (.A1_N(_07324_),
    .A2_N(_07406_),
    .B1(\design_top.MEM[22][14] ),
    .B2(_07408_),
    .X(_05027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09829_ (.A1_N(_07325_),
    .A2_N(_07406_),
    .B1(\design_top.MEM[22][13] ),
    .B2(_07408_),
    .X(_05026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09830_ (.A1_N(_07326_),
    .A2_N(_07406_),
    .B1(\design_top.MEM[22][12] ),
    .B2(_07408_),
    .X(_05025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09831_ (.A1_N(_07327_),
    .A2_N(_07406_),
    .B1(\design_top.MEM[22][11] ),
    .B2(_07408_),
    .X(_05024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09832_ (.A1_N(_07328_),
    .A2_N(_07405_),
    .B1(\design_top.MEM[22][10] ),
    .B2(_07407_),
    .X(_05023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09833_ (.A1_N(_07329_),
    .A2_N(_07405_),
    .B1(\design_top.MEM[22][9] ),
    .B2(_07407_),
    .X(_05022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09834_ (.A1_N(_07330_),
    .A2_N(_07405_),
    .B1(\design_top.MEM[22][8] ),
    .B2(_07407_),
    .X(_05021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09835_ (.A(_07301_),
    .B(_07353_),
    .X(_07409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09836_ (.A(_07409_),
    .X(_07410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09837_ (.A1(_07360_),
    .A2(_07132_),
    .B1(_07409_),
    .X(_07411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09838_ (.A(_07411_),
    .X(_07412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09839_ (.A1_N(_07331_),
    .A2_N(_07410_),
    .B1(\design_top.MEM[7][23] ),
    .B2(_07412_),
    .X(_05020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09840_ (.A1_N(_07337_),
    .A2_N(_07410_),
    .B1(\design_top.MEM[7][22] ),
    .B2(_07412_),
    .X(_05019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09841_ (.A1_N(_07338_),
    .A2_N(_07410_),
    .B1(\design_top.MEM[7][21] ),
    .B2(_07412_),
    .X(_05018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09842_ (.A1_N(_07339_),
    .A2_N(_07410_),
    .B1(\design_top.MEM[7][20] ),
    .B2(_07412_),
    .X(_05017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09843_ (.A1_N(_07340_),
    .A2_N(_07410_),
    .B1(\design_top.MEM[7][19] ),
    .B2(_07412_),
    .X(_05016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09844_ (.A1_N(_07341_),
    .A2_N(_07409_),
    .B1(\design_top.MEM[7][18] ),
    .B2(_07411_),
    .X(_05015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09845_ (.A1_N(_07342_),
    .A2_N(_07409_),
    .B1(\design_top.MEM[7][17] ),
    .B2(_07411_),
    .X(_05014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09846_ (.A1_N(_07343_),
    .A2_N(_07409_),
    .B1(\design_top.MEM[7][16] ),
    .B2(_07411_),
    .X(_05013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09847_ (.A(_06908_),
    .X(_07413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09848_ (.A(_06857_),
    .B(_06985_),
    .X(_07414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09849_ (.A(_07403_),
    .B(_07414_),
    .X(_07415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09850_ (.A(_07415_),
    .X(_07416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09851_ (.A1(_06975_),
    .A2(_06901_),
    .B1(_07415_),
    .X(_07417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09852_ (.A(_07417_),
    .X(_07418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09853_ (.A1_N(_07413_),
    .A2_N(_07416_),
    .B1(\design_top.MEM[8][15] ),
    .B2(_07418_),
    .X(_05012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09854_ (.A(_06918_),
    .X(_07419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09855_ (.A1_N(_07419_),
    .A2_N(_07416_),
    .B1(\design_top.MEM[8][14] ),
    .B2(_07418_),
    .X(_05011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09856_ (.A(_06921_),
    .X(_07420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09857_ (.A1_N(_07420_),
    .A2_N(_07416_),
    .B1(\design_top.MEM[8][13] ),
    .B2(_07418_),
    .X(_05010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09858_ (.A(_06924_),
    .X(_07421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09859_ (.A1_N(_07421_),
    .A2_N(_07416_),
    .B1(\design_top.MEM[8][12] ),
    .B2(_07418_),
    .X(_05009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09860_ (.A(_06927_),
    .X(_07422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09861_ (.A1_N(_07422_),
    .A2_N(_07416_),
    .B1(\design_top.MEM[8][11] ),
    .B2(_07418_),
    .X(_05008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09862_ (.A(_06930_),
    .X(_07423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09863_ (.A1_N(_07423_),
    .A2_N(_07415_),
    .B1(\design_top.MEM[8][10] ),
    .B2(_07417_),
    .X(_05007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09864_ (.A(_06933_),
    .X(_07424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09865_ (.A1_N(_07424_),
    .A2_N(_07415_),
    .B1(\design_top.MEM[8][9] ),
    .B2(_07417_),
    .X(_05006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09866_ (.A(_06936_),
    .X(_07425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09867_ (.A1_N(_07425_),
    .A2_N(_07415_),
    .B1(\design_top.MEM[8][8] ),
    .B2(_07417_),
    .X(_05005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09868_ (.A(_06942_),
    .X(_07426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09869_ (.A(_07426_),
    .B(_07414_),
    .X(_07427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09870_ (.A(_07427_),
    .X(_07428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09871_ (.A1(_06870_),
    .A2(_06901_),
    .B1(_07427_),
    .X(_07429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09872_ (.A(_07429_),
    .X(_07430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09873_ (.A1_N(_07331_),
    .A2_N(_07428_),
    .B1(\design_top.MEM[8][23] ),
    .B2(_07430_),
    .X(_05004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09874_ (.A1_N(_07337_),
    .A2_N(_07428_),
    .B1(\design_top.MEM[8][22] ),
    .B2(_07430_),
    .X(_05003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09875_ (.A1_N(_07338_),
    .A2_N(_07428_),
    .B1(\design_top.MEM[8][21] ),
    .B2(_07430_),
    .X(_05002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09876_ (.A1_N(_07339_),
    .A2_N(_07428_),
    .B1(\design_top.MEM[8][20] ),
    .B2(_07430_),
    .X(_05001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09877_ (.A1_N(_07340_),
    .A2_N(_07428_),
    .B1(\design_top.MEM[8][19] ),
    .B2(_07430_),
    .X(_05000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09878_ (.A1_N(_07341_),
    .A2_N(_07427_),
    .B1(\design_top.MEM[8][18] ),
    .B2(_07429_),
    .X(_04999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09879_ (.A1_N(_07342_),
    .A2_N(_07427_),
    .B1(\design_top.MEM[8][17] ),
    .B2(_07429_),
    .X(_04998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09880_ (.A1_N(_07343_),
    .A2_N(_07427_),
    .B1(\design_top.MEM[8][16] ),
    .B2(_07429_),
    .X(_04997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09881_ (.A(_06891_),
    .X(_07431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09882_ (.A(_07390_),
    .B(_07414_),
    .X(_07432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09883_ (.A(_07432_),
    .X(_07433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09884_ (.A1(_06870_),
    .A2(_06901_),
    .B1(_07432_),
    .X(_07434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09885_ (.A(_07434_),
    .X(_07435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09886_ (.A1_N(_07431_),
    .A2_N(_07433_),
    .B1(\design_top.MEM[8][31] ),
    .B2(_07435_),
    .X(_04996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09887_ (.A1_N(_07396_),
    .A2_N(_07433_),
    .B1(\design_top.MEM[8][30] ),
    .B2(_07435_),
    .X(_04995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09888_ (.A1_N(_07397_),
    .A2_N(_07433_),
    .B1(\design_top.MEM[8][29] ),
    .B2(_07435_),
    .X(_04994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09889_ (.A1_N(_07398_),
    .A2_N(_07433_),
    .B1(\design_top.MEM[8][28] ),
    .B2(_07435_),
    .X(_04993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09890_ (.A1_N(_07399_),
    .A2_N(_07433_),
    .B1(\design_top.MEM[8][27] ),
    .B2(_07435_),
    .X(_04992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09891_ (.A1_N(_07400_),
    .A2_N(_07432_),
    .B1(\design_top.MEM[8][26] ),
    .B2(_07434_),
    .X(_04991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09892_ (.A1_N(_07401_),
    .A2_N(_07432_),
    .B1(\design_top.MEM[8][25] ),
    .B2(_07434_),
    .X(_04990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09893_ (.A1_N(_07402_),
    .A2_N(_07432_),
    .B1(\design_top.MEM[8][24] ),
    .B2(_07434_),
    .X(_04989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09894_ (.A(_06939_),
    .X(_07436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09895_ (.A(_07042_),
    .B(_07363_),
    .X(_07437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09896_ (.A(_07426_),
    .B(_07437_),
    .X(_07438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09897_ (.A(_07438_),
    .X(_07439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09898_ (.A1(_07360_),
    .A2(_07393_),
    .B1(_07438_),
    .X(_07440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09899_ (.A(_07440_),
    .X(_07441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09900_ (.A1_N(_07436_),
    .A2_N(_07439_),
    .B1(\design_top.MEM[23][23] ),
    .B2(_07441_),
    .X(_04988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09901_ (.A(_06949_),
    .X(_07442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09902_ (.A1_N(_07442_),
    .A2_N(_07439_),
    .B1(\design_top.MEM[23][22] ),
    .B2(_07441_),
    .X(_04987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09903_ (.A(_06952_),
    .X(_07443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09904_ (.A1_N(_07443_),
    .A2_N(_07439_),
    .B1(\design_top.MEM[23][21] ),
    .B2(_07441_),
    .X(_04986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09905_ (.A(_06955_),
    .X(_07444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09906_ (.A1_N(_07444_),
    .A2_N(_07439_),
    .B1(\design_top.MEM[23][20] ),
    .B2(_07441_),
    .X(_04985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09907_ (.A(_06958_),
    .X(_07445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09908_ (.A1_N(_07445_),
    .A2_N(_07439_),
    .B1(\design_top.MEM[23][19] ),
    .B2(_07441_),
    .X(_04984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09909_ (.A(_06961_),
    .X(_07446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09910_ (.A1_N(_07446_),
    .A2_N(_07438_),
    .B1(\design_top.MEM[23][18] ),
    .B2(_07440_),
    .X(_04983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09911_ (.A(_06964_),
    .X(_07447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09912_ (.A1_N(_07447_),
    .A2_N(_07438_),
    .B1(\design_top.MEM[23][17] ),
    .B2(_07440_),
    .X(_04982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09913_ (.A(_06967_),
    .X(_07448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09914_ (.A1_N(_07448_),
    .A2_N(_07438_),
    .B1(\design_top.MEM[23][16] ),
    .B2(_07440_),
    .X(_04981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09915_ (.A(_06858_),
    .B(_06913_),
    .X(_07449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09916_ (.A(_07449_),
    .X(_07450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09917_ (.A(_07189_),
    .X(_07451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09918_ (.A1(_07451_),
    .A2(_06869_),
    .B1(_07449_),
    .X(_07452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09919_ (.A(_07452_),
    .X(_07453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09920_ (.A1_N(_07413_),
    .A2_N(_07450_),
    .B1(\design_top.MEM[9][15] ),
    .B2(_07453_),
    .X(_04980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09921_ (.A1_N(_07419_),
    .A2_N(_07450_),
    .B1(\design_top.MEM[9][14] ),
    .B2(_07453_),
    .X(_04979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09922_ (.A1_N(_07420_),
    .A2_N(_07450_),
    .B1(\design_top.MEM[9][13] ),
    .B2(_07453_),
    .X(_04978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09923_ (.A1_N(_07421_),
    .A2_N(_07450_),
    .B1(\design_top.MEM[9][12] ),
    .B2(_07453_),
    .X(_04977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09924_ (.A1_N(_07422_),
    .A2_N(_07450_),
    .B1(\design_top.MEM[9][11] ),
    .B2(_07453_),
    .X(_04976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09925_ (.A1_N(_07423_),
    .A2_N(_07449_),
    .B1(\design_top.MEM[9][10] ),
    .B2(_07452_),
    .X(_04975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09926_ (.A1_N(_07424_),
    .A2_N(_07449_),
    .B1(\design_top.MEM[9][9] ),
    .B2(_07452_),
    .X(_04974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09927_ (.A1_N(_07425_),
    .A2_N(_07449_),
    .B1(\design_top.MEM[9][8] ),
    .B2(_07452_),
    .X(_04973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09928_ (.A(_07390_),
    .B(_07437_),
    .X(_07454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09929_ (.A(_07454_),
    .X(_07455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09930_ (.A1(_07360_),
    .A2(_07393_),
    .B1(_07454_),
    .X(_07456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09931_ (.A(_07456_),
    .X(_07457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09932_ (.A1_N(_07431_),
    .A2_N(_07455_),
    .B1(\design_top.MEM[23][31] ),
    .B2(_07457_),
    .X(_04972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09933_ (.A1_N(_07396_),
    .A2_N(_07455_),
    .B1(\design_top.MEM[23][30] ),
    .B2(_07457_),
    .X(_04971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09934_ (.A1_N(_07397_),
    .A2_N(_07455_),
    .B1(\design_top.MEM[23][29] ),
    .B2(_07457_),
    .X(_04970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09935_ (.A1_N(_07398_),
    .A2_N(_07455_),
    .B1(\design_top.MEM[23][28] ),
    .B2(_07457_),
    .X(_04969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09936_ (.A1_N(_07399_),
    .A2_N(_07455_),
    .B1(\design_top.MEM[23][27] ),
    .B2(_07457_),
    .X(_04968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09937_ (.A1_N(_07400_),
    .A2_N(_07454_),
    .B1(\design_top.MEM[23][26] ),
    .B2(_07456_),
    .X(_04967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09938_ (.A1_N(_07401_),
    .A2_N(_07454_),
    .B1(\design_top.MEM[23][25] ),
    .B2(_07456_),
    .X(_04966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09939_ (.A1_N(_07402_),
    .A2_N(_07454_),
    .B1(\design_top.MEM[23][24] ),
    .B2(_07456_),
    .X(_04965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09940_ (.A(_01371_),
    .B(_07058_),
    .X(_07458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09941_ (.A(_06894_),
    .B(_07458_),
    .X(_07459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09942_ (.A(_07403_),
    .B(_07459_),
    .X(_07460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09943_ (.A(_07460_),
    .X(_07461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _09944_ (.A(_07064_),
    .B(_06867_),
    .C(wbs_adr_i[0]),
    .X(_07462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09945_ (.A(_07462_),
    .X(_07463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09946_ (.A(_07463_),
    .X(_07464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09947_ (.A1(_07374_),
    .A2(_07464_),
    .B1(_07460_),
    .X(_07465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09948_ (.A(_07465_),
    .X(_07466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09949_ (.A1_N(_07413_),
    .A2_N(_07461_),
    .B1(\design_top.MEM[24][15] ),
    .B2(_07466_),
    .X(_04964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09950_ (.A1_N(_07419_),
    .A2_N(_07461_),
    .B1(\design_top.MEM[24][14] ),
    .B2(_07466_),
    .X(_04963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09951_ (.A1_N(_07420_),
    .A2_N(_07461_),
    .B1(\design_top.MEM[24][13] ),
    .B2(_07466_),
    .X(_04962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09952_ (.A1_N(_07421_),
    .A2_N(_07461_),
    .B1(\design_top.MEM[24][12] ),
    .B2(_07466_),
    .X(_04961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09953_ (.A1_N(_07422_),
    .A2_N(_07461_),
    .B1(\design_top.MEM[24][11] ),
    .B2(_07466_),
    .X(_04960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09954_ (.A1_N(_07423_),
    .A2_N(_07460_),
    .B1(\design_top.MEM[24][10] ),
    .B2(_07465_),
    .X(_04959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09955_ (.A1_N(_07424_),
    .A2_N(_07460_),
    .B1(\design_top.MEM[24][9] ),
    .B2(_07465_),
    .X(_04958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09956_ (.A1_N(_07425_),
    .A2_N(_07460_),
    .B1(\design_top.MEM[24][8] ),
    .B2(_07465_),
    .X(_04957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09957_ (.A(_06858_),
    .B(_06944_),
    .X(_07467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09958_ (.A(_07467_),
    .X(_07468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09959_ (.A1(_07451_),
    .A2(_06869_),
    .B1(_07467_),
    .X(_07469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09960_ (.A(_07469_),
    .X(_07470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09961_ (.A1_N(_07436_),
    .A2_N(_07468_),
    .B1(\design_top.MEM[9][23] ),
    .B2(_07470_),
    .X(_04956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09962_ (.A1_N(_07442_),
    .A2_N(_07468_),
    .B1(\design_top.MEM[9][22] ),
    .B2(_07470_),
    .X(_04955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09963_ (.A1_N(_07443_),
    .A2_N(_07468_),
    .B1(\design_top.MEM[9][21] ),
    .B2(_07470_),
    .X(_04954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09964_ (.A1_N(_07444_),
    .A2_N(_07468_),
    .B1(\design_top.MEM[9][20] ),
    .B2(_07470_),
    .X(_04953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09965_ (.A1_N(_07445_),
    .A2_N(_07468_),
    .B1(\design_top.MEM[9][19] ),
    .B2(_07470_),
    .X(_04952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09966_ (.A1_N(_07446_),
    .A2_N(_07467_),
    .B1(\design_top.MEM[9][18] ),
    .B2(_07469_),
    .X(_04951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09967_ (.A1_N(_07447_),
    .A2_N(_07467_),
    .B1(\design_top.MEM[9][17] ),
    .B2(_07469_),
    .X(_04950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09968_ (.A1_N(_07448_),
    .A2_N(_07467_),
    .B1(\design_top.MEM[9][16] ),
    .B2(_07469_),
    .X(_04949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09969_ (.A(_07426_),
    .B(_07459_),
    .X(_07471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09970_ (.A(_07471_),
    .X(_07472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09971_ (.A1(_07374_),
    .A2(_07464_),
    .B1(_07471_),
    .X(_07473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09972_ (.A(_07473_),
    .X(_07474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09973_ (.A1_N(_07436_),
    .A2_N(_07472_),
    .B1(\design_top.MEM[24][23] ),
    .B2(_07474_),
    .X(_04948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09974_ (.A1_N(_07442_),
    .A2_N(_07472_),
    .B1(\design_top.MEM[24][22] ),
    .B2(_07474_),
    .X(_04947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09975_ (.A1_N(_07443_),
    .A2_N(_07472_),
    .B1(\design_top.MEM[24][21] ),
    .B2(_07474_),
    .X(_04946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09976_ (.A1_N(_07444_),
    .A2_N(_07472_),
    .B1(\design_top.MEM[24][20] ),
    .B2(_07474_),
    .X(_04945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09977_ (.A1_N(_07445_),
    .A2_N(_07472_),
    .B1(\design_top.MEM[24][19] ),
    .B2(_07474_),
    .X(_04944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09978_ (.A1_N(_07446_),
    .A2_N(_07471_),
    .B1(\design_top.MEM[24][18] ),
    .B2(_07473_),
    .X(_04943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09979_ (.A1_N(_07447_),
    .A2_N(_07471_),
    .B1(\design_top.MEM[24][17] ),
    .B2(_07473_),
    .X(_04942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09980_ (.A1_N(_07448_),
    .A2_N(_07471_),
    .B1(\design_top.MEM[24][16] ),
    .B2(_07473_),
    .X(_04941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09981_ (.A(_07390_),
    .B(_07459_),
    .X(_07475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09982_ (.A(_07475_),
    .X(_07476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09983_ (.A1(_07374_),
    .A2(_07464_),
    .B1(_07475_),
    .X(_07477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09984_ (.A(_07477_),
    .X(_07478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09985_ (.A1_N(_07431_),
    .A2_N(_07476_),
    .B1(\design_top.MEM[24][31] ),
    .B2(_07478_),
    .X(_04940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09986_ (.A1_N(_07396_),
    .A2_N(_07476_),
    .B1(\design_top.MEM[24][30] ),
    .B2(_07478_),
    .X(_04939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09987_ (.A1_N(_07397_),
    .A2_N(_07476_),
    .B1(\design_top.MEM[24][29] ),
    .B2(_07478_),
    .X(_04938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09988_ (.A1_N(_07398_),
    .A2_N(_07476_),
    .B1(\design_top.MEM[24][28] ),
    .B2(_07478_),
    .X(_04937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09989_ (.A1_N(_07399_),
    .A2_N(_07476_),
    .B1(\design_top.MEM[24][27] ),
    .B2(_07478_),
    .X(_04936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09990_ (.A1_N(_07400_),
    .A2_N(_07475_),
    .B1(\design_top.MEM[24][26] ),
    .B2(_07477_),
    .X(_04935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09991_ (.A1_N(_07401_),
    .A2_N(_07475_),
    .B1(\design_top.MEM[24][25] ),
    .B2(_07477_),
    .X(_04934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09992_ (.A1_N(_07402_),
    .A2_N(_07475_),
    .B1(\design_top.MEM[24][24] ),
    .B2(_07477_),
    .X(_04933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09993_ (.A(_06851_),
    .B(_07458_),
    .X(_07479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _09994_ (.A(_07403_),
    .B(_07479_),
    .X(_07480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09995_ (.A(_07480_),
    .X(_07481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _09996_ (.A1(_07451_),
    .A2(_07464_),
    .B1(_07480_),
    .X(_07482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _09997_ (.A(_07482_),
    .X(_07483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09998_ (.A1_N(_07413_),
    .A2_N(_07481_),
    .B1(\design_top.MEM[25][15] ),
    .B2(_07483_),
    .X(_04932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _09999_ (.A1_N(_07419_),
    .A2_N(_07481_),
    .B1(\design_top.MEM[25][14] ),
    .B2(_07483_),
    .X(_04931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10000_ (.A1_N(_07420_),
    .A2_N(_07481_),
    .B1(\design_top.MEM[25][13] ),
    .B2(_07483_),
    .X(_04930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10001_ (.A1_N(_07421_),
    .A2_N(_07481_),
    .B1(\design_top.MEM[25][12] ),
    .B2(_07483_),
    .X(_04929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10002_ (.A1_N(_07422_),
    .A2_N(_07481_),
    .B1(\design_top.MEM[25][11] ),
    .B2(_07483_),
    .X(_04928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10003_ (.A1_N(_07423_),
    .A2_N(_07480_),
    .B1(\design_top.MEM[25][10] ),
    .B2(_07482_),
    .X(_04927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10004_ (.A1_N(_07424_),
    .A2_N(_07480_),
    .B1(\design_top.MEM[25][9] ),
    .B2(_07482_),
    .X(_04926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10005_ (.A1_N(_07425_),
    .A2_N(_07480_),
    .B1(\design_top.MEM[25][8] ),
    .B2(_07482_),
    .X(_04925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10006_ (.A(_07426_),
    .B(_07479_),
    .X(_07484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10007_ (.A(_07484_),
    .X(_07485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10008_ (.A1(_07451_),
    .A2(_07464_),
    .B1(_07484_),
    .X(_07486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10009_ (.A(_07486_),
    .X(_07487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10010_ (.A1_N(_07436_),
    .A2_N(_07485_),
    .B1(\design_top.MEM[25][23] ),
    .B2(_07487_),
    .X(_04924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10011_ (.A1_N(_07442_),
    .A2_N(_07485_),
    .B1(\design_top.MEM[25][22] ),
    .B2(_07487_),
    .X(_04923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10012_ (.A1_N(_07443_),
    .A2_N(_07485_),
    .B1(\design_top.MEM[25][21] ),
    .B2(_07487_),
    .X(_04922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10013_ (.A1_N(_07444_),
    .A2_N(_07485_),
    .B1(\design_top.MEM[25][20] ),
    .B2(_07487_),
    .X(_04921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10014_ (.A1_N(_07445_),
    .A2_N(_07485_),
    .B1(\design_top.MEM[25][19] ),
    .B2(_07487_),
    .X(_04920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10015_ (.A1_N(_07446_),
    .A2_N(_07484_),
    .B1(\design_top.MEM[25][18] ),
    .B2(_07486_),
    .X(_04919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10016_ (.A1_N(_07447_),
    .A2_N(_07484_),
    .B1(\design_top.MEM[25][17] ),
    .B2(_07486_),
    .X(_04918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10017_ (.A1_N(_07448_),
    .A2_N(_07484_),
    .B1(\design_top.MEM[25][16] ),
    .B2(_07486_),
    .X(_04917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10018_ (.A(_07390_),
    .B(_07479_),
    .X(_07488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10019_ (.A(_07488_),
    .X(_07489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10020_ (.A(_07463_),
    .X(_07490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10021_ (.A1(_07451_),
    .A2(_07490_),
    .B1(_07488_),
    .X(_07491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10022_ (.A(_07491_),
    .X(_07492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10023_ (.A1_N(_07431_),
    .A2_N(_07489_),
    .B1(\design_top.MEM[25][31] ),
    .B2(_07492_),
    .X(_04916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10024_ (.A1_N(_07396_),
    .A2_N(_07489_),
    .B1(\design_top.MEM[25][30] ),
    .B2(_07492_),
    .X(_04915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10025_ (.A1_N(_07397_),
    .A2_N(_07489_),
    .B1(\design_top.MEM[25][29] ),
    .B2(_07492_),
    .X(_04914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10026_ (.A1_N(_07398_),
    .A2_N(_07489_),
    .B1(\design_top.MEM[25][28] ),
    .B2(_07492_),
    .X(_04913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10027_ (.A1_N(_07399_),
    .A2_N(_07489_),
    .B1(\design_top.MEM[25][27] ),
    .B2(_07492_),
    .X(_04912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10028_ (.A1_N(_07400_),
    .A2_N(_07488_),
    .B1(\design_top.MEM[25][26] ),
    .B2(_07491_),
    .X(_04911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10029_ (.A1_N(_07401_),
    .A2_N(_07488_),
    .B1(\design_top.MEM[25][25] ),
    .B2(_07491_),
    .X(_04910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10030_ (.A1_N(_07402_),
    .A2_N(_07488_),
    .B1(\design_top.MEM[25][24] ),
    .B2(_07491_),
    .X(_04909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10031_ (.A(_06970_),
    .B(_07458_),
    .X(_07493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10032_ (.A(_07403_),
    .B(_07493_),
    .X(_07494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10033_ (.A(_07494_),
    .X(_07495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10034_ (.A1(_07292_),
    .A2(_07490_),
    .B1(_07494_),
    .X(_07496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10035_ (.A(_07496_),
    .X(_07497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10036_ (.A1_N(_07413_),
    .A2_N(_07495_),
    .B1(\design_top.MEM[26][15] ),
    .B2(_07497_),
    .X(_04908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10037_ (.A1_N(_07419_),
    .A2_N(_07495_),
    .B1(\design_top.MEM[26][14] ),
    .B2(_07497_),
    .X(_04907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10038_ (.A1_N(_07420_),
    .A2_N(_07495_),
    .B1(\design_top.MEM[26][13] ),
    .B2(_07497_),
    .X(_04906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10039_ (.A1_N(_07421_),
    .A2_N(_07495_),
    .B1(\design_top.MEM[26][12] ),
    .B2(_07497_),
    .X(_04905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10040_ (.A1_N(_07422_),
    .A2_N(_07495_),
    .B1(\design_top.MEM[26][11] ),
    .B2(_07497_),
    .X(_04904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10041_ (.A1_N(_07423_),
    .A2_N(_07494_),
    .B1(\design_top.MEM[26][10] ),
    .B2(_07496_),
    .X(_04903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10042_ (.A1_N(_07424_),
    .A2_N(_07494_),
    .B1(\design_top.MEM[26][9] ),
    .B2(_07496_),
    .X(_04902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10043_ (.A1_N(_07425_),
    .A2_N(_07494_),
    .B1(\design_top.MEM[26][8] ),
    .B2(_07496_),
    .X(_04901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10044_ (.A(_07426_),
    .B(_07404_),
    .X(_07498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10045_ (.A(_07498_),
    .X(_07499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10046_ (.A1(_07292_),
    .A2(_07393_),
    .B1(_07498_),
    .X(_07500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10047_ (.A(_07500_),
    .X(_07501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10048_ (.A1_N(_07436_),
    .A2_N(_07499_),
    .B1(\design_top.MEM[22][23] ),
    .B2(_07501_),
    .X(_04900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10049_ (.A1_N(_07442_),
    .A2_N(_07499_),
    .B1(\design_top.MEM[22][22] ),
    .B2(_07501_),
    .X(_04899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10050_ (.A1_N(_07443_),
    .A2_N(_07499_),
    .B1(\design_top.MEM[22][21] ),
    .B2(_07501_),
    .X(_04898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10051_ (.A1_N(_07444_),
    .A2_N(_07499_),
    .B1(\design_top.MEM[22][20] ),
    .B2(_07501_),
    .X(_04897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10052_ (.A1_N(_07445_),
    .A2_N(_07499_),
    .B1(\design_top.MEM[22][19] ),
    .B2(_07501_),
    .X(_04896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10053_ (.A1_N(_07446_),
    .A2_N(_07498_),
    .B1(\design_top.MEM[22][18] ),
    .B2(_07500_),
    .X(_04895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10054_ (.A1_N(_07447_),
    .A2_N(_07498_),
    .B1(\design_top.MEM[22][17] ),
    .B2(_07500_),
    .X(_04894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10055_ (.A1_N(_07448_),
    .A2_N(_07498_),
    .B1(\design_top.MEM[22][16] ),
    .B2(_07500_),
    .X(_04893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10056_ (.A(_06844_),
    .X(_07502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10057_ (.A(_07502_),
    .B(_07404_),
    .X(_07503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10058_ (.A(_07503_),
    .X(_07504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10059_ (.A1(_06978_),
    .A2(_07368_),
    .B1(_07503_),
    .X(_07505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10060_ (.A(_07505_),
    .X(_07506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10061_ (.A1_N(_07431_),
    .A2_N(_07504_),
    .B1(\design_top.MEM[22][31] ),
    .B2(_07506_),
    .X(_04892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10062_ (.A(_06655_),
    .X(_07507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10063_ (.A1_N(_07507_),
    .A2_N(_07504_),
    .B1(\design_top.MEM[22][30] ),
    .B2(_07506_),
    .X(_04891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10064_ (.A(_06873_),
    .X(_07508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10065_ (.A1_N(_07508_),
    .A2_N(_07504_),
    .B1(\design_top.MEM[22][29] ),
    .B2(_07506_),
    .X(_04890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10066_ (.A(_06876_),
    .X(_07509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10067_ (.A1_N(_07509_),
    .A2_N(_07504_),
    .B1(\design_top.MEM[22][28] ),
    .B2(_07506_),
    .X(_04889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10068_ (.A(_06879_),
    .X(_07510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10069_ (.A1_N(_07510_),
    .A2_N(_07504_),
    .B1(\design_top.MEM[22][27] ),
    .B2(_07506_),
    .X(_04888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10070_ (.A(_06882_),
    .X(_07511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10071_ (.A1_N(_07511_),
    .A2_N(_07503_),
    .B1(\design_top.MEM[22][26] ),
    .B2(_07505_),
    .X(_04887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10072_ (.A(_06885_),
    .X(_07512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10073_ (.A1_N(_07512_),
    .A2_N(_07503_),
    .B1(\design_top.MEM[22][25] ),
    .B2(_07505_),
    .X(_04886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10074_ (.A(_06888_),
    .X(_07513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10075_ (.A1_N(_07513_),
    .A2_N(_07503_),
    .B1(\design_top.MEM[22][24] ),
    .B2(_07505_),
    .X(_04885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10076_ (.A(_06939_),
    .X(_07514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10077_ (.A(_06942_),
    .X(_07515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10078_ (.A(_07515_),
    .B(_07493_),
    .X(_07516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10079_ (.A(_07516_),
    .X(_07517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10080_ (.A1(_06978_),
    .A2(_07490_),
    .B1(_07516_),
    .X(_07518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10081_ (.A(_07518_),
    .X(_07519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10082_ (.A1_N(_07514_),
    .A2_N(_07517_),
    .B1(\design_top.MEM[26][23] ),
    .B2(_07519_),
    .X(_04884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10083_ (.A(_06949_),
    .X(_07520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10084_ (.A1_N(_07520_),
    .A2_N(_07517_),
    .B1(\design_top.MEM[26][22] ),
    .B2(_07519_),
    .X(_04883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10085_ (.A(_06952_),
    .X(_07521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10086_ (.A1_N(_07521_),
    .A2_N(_07517_),
    .B1(\design_top.MEM[26][21] ),
    .B2(_07519_),
    .X(_04882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10087_ (.A(_06955_),
    .X(_07522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10088_ (.A1_N(_07522_),
    .A2_N(_07517_),
    .B1(\design_top.MEM[26][20] ),
    .B2(_07519_),
    .X(_04881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10089_ (.A(_06958_),
    .X(_07523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10090_ (.A1_N(_07523_),
    .A2_N(_07517_),
    .B1(\design_top.MEM[26][19] ),
    .B2(_07519_),
    .X(_04880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10091_ (.A(_06961_),
    .X(_07524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10092_ (.A1_N(_07524_),
    .A2_N(_07516_),
    .B1(\design_top.MEM[26][18] ),
    .B2(_07518_),
    .X(_04879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10093_ (.A(_06964_),
    .X(_07525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10094_ (.A1_N(_07525_),
    .A2_N(_07516_),
    .B1(\design_top.MEM[26][17] ),
    .B2(_07518_),
    .X(_04878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10095_ (.A(_06967_),
    .X(_07526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10096_ (.A1_N(_07526_),
    .A2_N(_07516_),
    .B1(\design_top.MEM[26][16] ),
    .B2(_07518_),
    .X(_04877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10097_ (.A(_06891_),
    .X(_07527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10098_ (.A(_07502_),
    .B(_07493_),
    .X(_07528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10099_ (.A(_07528_),
    .X(_07529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10100_ (.A1(_06978_),
    .A2(_07490_),
    .B1(_07528_),
    .X(_07530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10101_ (.A(_07530_),
    .X(_07531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10102_ (.A1_N(_07527_),
    .A2_N(_07529_),
    .B1(\design_top.MEM[26][31] ),
    .B2(_07531_),
    .X(_04876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10103_ (.A1_N(_07507_),
    .A2_N(_07529_),
    .B1(\design_top.MEM[26][30] ),
    .B2(_07531_),
    .X(_04875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10104_ (.A1_N(_07508_),
    .A2_N(_07529_),
    .B1(\design_top.MEM[26][29] ),
    .B2(_07531_),
    .X(_04874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10105_ (.A1_N(_07509_),
    .A2_N(_07529_),
    .B1(\design_top.MEM[26][28] ),
    .B2(_07531_),
    .X(_04873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10106_ (.A1_N(_07510_),
    .A2_N(_07529_),
    .B1(\design_top.MEM[26][27] ),
    .B2(_07531_),
    .X(_04872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10107_ (.A1_N(_07511_),
    .A2_N(_07528_),
    .B1(\design_top.MEM[26][26] ),
    .B2(_07530_),
    .X(_04871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10108_ (.A1_N(_07512_),
    .A2_N(_07528_),
    .B1(\design_top.MEM[26][25] ),
    .B2(_07530_),
    .X(_04870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10109_ (.A1_N(_07513_),
    .A2_N(_07528_),
    .B1(\design_top.MEM[26][24] ),
    .B2(_07530_),
    .X(_04869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10110_ (.A(_06908_),
    .X(_07532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10111_ (.A(_06911_),
    .X(_07533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10112_ (.A(_07042_),
    .B(_07458_),
    .X(_07534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10113_ (.A(_07533_),
    .B(_07534_),
    .X(_07535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10114_ (.A(_07535_),
    .X(_07536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10115_ (.A1(_07360_),
    .A2(_07490_),
    .B1(_07535_),
    .X(_07537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10116_ (.A(_07537_),
    .X(_07538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10117_ (.A1_N(_07532_),
    .A2_N(_07536_),
    .B1(\design_top.MEM[27][15] ),
    .B2(_07538_),
    .X(_04868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10118_ (.A(_06918_),
    .X(_07539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10119_ (.A1_N(_07539_),
    .A2_N(_07536_),
    .B1(\design_top.MEM[27][14] ),
    .B2(_07538_),
    .X(_04867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10120_ (.A(_06921_),
    .X(_07540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10121_ (.A1_N(_07540_),
    .A2_N(_07536_),
    .B1(\design_top.MEM[27][13] ),
    .B2(_07538_),
    .X(_04866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10122_ (.A(_06924_),
    .X(_07541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10123_ (.A1_N(_07541_),
    .A2_N(_07536_),
    .B1(\design_top.MEM[27][12] ),
    .B2(_07538_),
    .X(_04865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10124_ (.A(_06927_),
    .X(_07542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10125_ (.A1_N(_07542_),
    .A2_N(_07536_),
    .B1(\design_top.MEM[27][11] ),
    .B2(_07538_),
    .X(_04864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10126_ (.A(_06930_),
    .X(_07543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10127_ (.A1_N(_07543_),
    .A2_N(_07535_),
    .B1(\design_top.MEM[27][10] ),
    .B2(_07537_),
    .X(_04863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10128_ (.A(_06933_),
    .X(_07544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10129_ (.A1_N(_07544_),
    .A2_N(_07535_),
    .B1(\design_top.MEM[27][9] ),
    .B2(_07537_),
    .X(_04862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10130_ (.A(_06936_),
    .X(_07545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10131_ (.A1_N(_07545_),
    .A2_N(_07535_),
    .B1(\design_top.MEM[27][8] ),
    .B2(_07537_),
    .X(_04861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10132_ (.A(_07515_),
    .B(_07534_),
    .X(_07546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10133_ (.A(_07546_),
    .X(_07547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10134_ (.A1(_07049_),
    .A2(_07463_),
    .B1(_07546_),
    .X(_07548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10135_ (.A(_07548_),
    .X(_07549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10136_ (.A1_N(_07514_),
    .A2_N(_07547_),
    .B1(\design_top.MEM[27][23] ),
    .B2(_07549_),
    .X(_04860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10137_ (.A1_N(_07520_),
    .A2_N(_07547_),
    .B1(\design_top.MEM[27][22] ),
    .B2(_07549_),
    .X(_04859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10138_ (.A1_N(_07521_),
    .A2_N(_07547_),
    .B1(\design_top.MEM[27][21] ),
    .B2(_07549_),
    .X(_04858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10139_ (.A1_N(_07522_),
    .A2_N(_07547_),
    .B1(\design_top.MEM[27][20] ),
    .B2(_07549_),
    .X(_04857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10140_ (.A1_N(_07523_),
    .A2_N(_07547_),
    .B1(\design_top.MEM[27][19] ),
    .B2(_07549_),
    .X(_04856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10141_ (.A1_N(_07524_),
    .A2_N(_07546_),
    .B1(\design_top.MEM[27][18] ),
    .B2(_07548_),
    .X(_04855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10142_ (.A1_N(_07525_),
    .A2_N(_07546_),
    .B1(\design_top.MEM[27][17] ),
    .B2(_07548_),
    .X(_04854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10143_ (.A1_N(_07526_),
    .A2_N(_07546_),
    .B1(\design_top.MEM[27][16] ),
    .B2(_07548_),
    .X(_04853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10144_ (.A(_07502_),
    .B(_07534_),
    .X(_07550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10145_ (.A(_07550_),
    .X(_07551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10146_ (.A1(_07049_),
    .A2(_07463_),
    .B1(_07550_),
    .X(_07552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10147_ (.A(_07552_),
    .X(_07553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10148_ (.A1_N(_07527_),
    .A2_N(_07551_),
    .B1(\design_top.MEM[27][31] ),
    .B2(_07553_),
    .X(_04852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10149_ (.A1_N(_07507_),
    .A2_N(_07551_),
    .B1(\design_top.MEM[27][30] ),
    .B2(_07553_),
    .X(_04851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10150_ (.A1_N(_07508_),
    .A2_N(_07551_),
    .B1(\design_top.MEM[27][29] ),
    .B2(_07553_),
    .X(_04850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10151_ (.A1_N(_07509_),
    .A2_N(_07551_),
    .B1(\design_top.MEM[27][28] ),
    .B2(_07553_),
    .X(_04849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10152_ (.A1_N(_07510_),
    .A2_N(_07551_),
    .B1(\design_top.MEM[27][27] ),
    .B2(_07553_),
    .X(_04848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10153_ (.A1_N(_07511_),
    .A2_N(_07550_),
    .B1(\design_top.MEM[27][26] ),
    .B2(_07552_),
    .X(_04847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10154_ (.A1_N(_07512_),
    .A2_N(_07550_),
    .B1(\design_top.MEM[27][25] ),
    .B2(_07552_),
    .X(_04846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10155_ (.A1_N(_07513_),
    .A2_N(_07550_),
    .B1(\design_top.MEM[27][24] ),
    .B2(_07552_),
    .X(_04845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10156_ (.A(_06894_),
    .B(_07059_),
    .X(_07554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10157_ (.A(_07533_),
    .B(_07554_),
    .X(_07555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10158_ (.A(_07555_),
    .X(_07556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10159_ (.A(_07150_),
    .X(_07557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10160_ (.A1(_07557_),
    .A2(_07094_),
    .B1(_07555_),
    .X(_07558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10161_ (.A(_07558_),
    .X(_07559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10162_ (.A1_N(_07532_),
    .A2_N(_07556_),
    .B1(\design_top.MEM[28][15] ),
    .B2(_07559_),
    .X(_04844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10163_ (.A1_N(_07539_),
    .A2_N(_07556_),
    .B1(\design_top.MEM[28][14] ),
    .B2(_07559_),
    .X(_04843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10164_ (.A1_N(_07540_),
    .A2_N(_07556_),
    .B1(\design_top.MEM[28][13] ),
    .B2(_07559_),
    .X(_04842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10165_ (.A1_N(_07541_),
    .A2_N(_07556_),
    .B1(\design_top.MEM[28][12] ),
    .B2(_07559_),
    .X(_04841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10166_ (.A1_N(_07542_),
    .A2_N(_07556_),
    .B1(\design_top.MEM[28][11] ),
    .B2(_07559_),
    .X(_04840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10167_ (.A1_N(_07543_),
    .A2_N(_07555_),
    .B1(\design_top.MEM[28][10] ),
    .B2(_07558_),
    .X(_04839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10168_ (.A1_N(_07544_),
    .A2_N(_07555_),
    .B1(\design_top.MEM[28][9] ),
    .B2(_07558_),
    .X(_04838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10169_ (.A1_N(_07545_),
    .A2_N(_07555_),
    .B1(\design_top.MEM[28][8] ),
    .B2(_07558_),
    .X(_04837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10170_ (.A(_07515_),
    .B(_07554_),
    .X(_07560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10171_ (.A(_07560_),
    .X(_07561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10172_ (.A1(_07557_),
    .A2(_07094_),
    .B1(_07560_),
    .X(_07562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10173_ (.A(_07562_),
    .X(_07563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10174_ (.A1_N(_07514_),
    .A2_N(_07561_),
    .B1(\design_top.MEM[28][23] ),
    .B2(_07563_),
    .X(_04836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10175_ (.A1_N(_07520_),
    .A2_N(_07561_),
    .B1(\design_top.MEM[28][22] ),
    .B2(_07563_),
    .X(_04835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10176_ (.A1_N(_07521_),
    .A2_N(_07561_),
    .B1(\design_top.MEM[28][21] ),
    .B2(_07563_),
    .X(_04834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10177_ (.A1_N(_07522_),
    .A2_N(_07561_),
    .B1(\design_top.MEM[28][20] ),
    .B2(_07563_),
    .X(_04833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10178_ (.A1_N(_07523_),
    .A2_N(_07561_),
    .B1(\design_top.MEM[28][19] ),
    .B2(_07563_),
    .X(_04832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10179_ (.A1_N(_07524_),
    .A2_N(_07560_),
    .B1(\design_top.MEM[28][18] ),
    .B2(_07562_),
    .X(_04831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10180_ (.A1_N(_07525_),
    .A2_N(_07560_),
    .B1(\design_top.MEM[28][17] ),
    .B2(_07562_),
    .X(_04830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10181_ (.A1_N(_07526_),
    .A2_N(_07560_),
    .B1(\design_top.MEM[28][16] ),
    .B2(_07562_),
    .X(_04829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10182_ (.A(_07502_),
    .B(_07554_),
    .X(_07564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10183_ (.A(_07564_),
    .X(_07565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10184_ (.A1(_07557_),
    .A2(_07094_),
    .B1(_07564_),
    .X(_07566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10185_ (.A(_07566_),
    .X(_07567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10186_ (.A1_N(_07527_),
    .A2_N(_07565_),
    .B1(\design_top.MEM[28][31] ),
    .B2(_07567_),
    .X(_04828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10187_ (.A1_N(_07507_),
    .A2_N(_07565_),
    .B1(\design_top.MEM[28][30] ),
    .B2(_07567_),
    .X(_04827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10188_ (.A1_N(_07508_),
    .A2_N(_07565_),
    .B1(\design_top.MEM[28][29] ),
    .B2(_07567_),
    .X(_04826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10189_ (.A1_N(_07509_),
    .A2_N(_07565_),
    .B1(\design_top.MEM[28][28] ),
    .B2(_07567_),
    .X(_04825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10190_ (.A1_N(_07510_),
    .A2_N(_07565_),
    .B1(\design_top.MEM[28][27] ),
    .B2(_07567_),
    .X(_04824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10191_ (.A1_N(_07511_),
    .A2_N(_07564_),
    .B1(\design_top.MEM[28][26] ),
    .B2(_07566_),
    .X(_04823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10192_ (.A1_N(_07512_),
    .A2_N(_07564_),
    .B1(\design_top.MEM[28][25] ),
    .B2(_07566_),
    .X(_04822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10193_ (.A1_N(_07513_),
    .A2_N(_07564_),
    .B1(\design_top.MEM[28][24] ),
    .B2(_07566_),
    .X(_04821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10194_ (.A(_06851_),
    .B(_07059_),
    .X(_07568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10195_ (.A(_07533_),
    .B(_07568_),
    .X(_07569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10196_ (.A(_07569_),
    .X(_07570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10197_ (.A1(_06865_),
    .A2(_07094_),
    .B1(_07569_),
    .X(_07571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10198_ (.A(_07571_),
    .X(_07572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10199_ (.A1_N(_07532_),
    .A2_N(_07570_),
    .B1(\design_top.MEM[29][15] ),
    .B2(_07572_),
    .X(_04820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10200_ (.A1_N(_07539_),
    .A2_N(_07570_),
    .B1(\design_top.MEM[29][14] ),
    .B2(_07572_),
    .X(_04819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10201_ (.A1_N(_07540_),
    .A2_N(_07570_),
    .B1(\design_top.MEM[29][13] ),
    .B2(_07572_),
    .X(_04818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10202_ (.A1_N(_07541_),
    .A2_N(_07570_),
    .B1(\design_top.MEM[29][12] ),
    .B2(_07572_),
    .X(_04817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10203_ (.A1_N(_07542_),
    .A2_N(_07570_),
    .B1(\design_top.MEM[29][11] ),
    .B2(_07572_),
    .X(_04816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10204_ (.A1_N(_07543_),
    .A2_N(_07569_),
    .B1(\design_top.MEM[29][10] ),
    .B2(_07571_),
    .X(_04815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10205_ (.A1_N(_07544_),
    .A2_N(_07569_),
    .B1(\design_top.MEM[29][9] ),
    .B2(_07571_),
    .X(_04814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10206_ (.A1_N(_07545_),
    .A2_N(_07569_),
    .B1(\design_top.MEM[29][8] ),
    .B2(_07571_),
    .X(_04813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10207_ (.A(_07533_),
    .B(_07437_),
    .X(_07573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10208_ (.A(_07573_),
    .X(_07574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10209_ (.A1(_07049_),
    .A2(_07368_),
    .B1(_07573_),
    .X(_07575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10210_ (.A(_07575_),
    .X(_07576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10211_ (.A1_N(_07532_),
    .A2_N(_07574_),
    .B1(\design_top.MEM[23][15] ),
    .B2(_07576_),
    .X(_04812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10212_ (.A1_N(_07539_),
    .A2_N(_07574_),
    .B1(\design_top.MEM[23][14] ),
    .B2(_07576_),
    .X(_04811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10213_ (.A1_N(_07540_),
    .A2_N(_07574_),
    .B1(\design_top.MEM[23][13] ),
    .B2(_07576_),
    .X(_04810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10214_ (.A1_N(_07541_),
    .A2_N(_07574_),
    .B1(\design_top.MEM[23][12] ),
    .B2(_07576_),
    .X(_04809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10215_ (.A1_N(_07542_),
    .A2_N(_07574_),
    .B1(\design_top.MEM[23][11] ),
    .B2(_07576_),
    .X(_04808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10216_ (.A1_N(_07543_),
    .A2_N(_07573_),
    .B1(\design_top.MEM[23][10] ),
    .B2(_07575_),
    .X(_04807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10217_ (.A1_N(_07544_),
    .A2_N(_07573_),
    .B1(\design_top.MEM[23][9] ),
    .B2(_07575_),
    .X(_04806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10218_ (.A1_N(_07545_),
    .A2_N(_07573_),
    .B1(\design_top.MEM[23][8] ),
    .B2(_07575_),
    .X(_04805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10219_ (.A(_07515_),
    .B(_07568_),
    .X(_07577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10220_ (.A(_07577_),
    .X(_07578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10221_ (.A1(_06865_),
    .A2(_07067_),
    .B1(_07577_),
    .X(_07579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10222_ (.A(_07579_),
    .X(_07580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10223_ (.A1_N(_07514_),
    .A2_N(_07578_),
    .B1(\design_top.MEM[29][23] ),
    .B2(_07580_),
    .X(_04804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10224_ (.A1_N(_07520_),
    .A2_N(_07578_),
    .B1(\design_top.MEM[29][22] ),
    .B2(_07580_),
    .X(_04803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10225_ (.A1_N(_07521_),
    .A2_N(_07578_),
    .B1(\design_top.MEM[29][21] ),
    .B2(_07580_),
    .X(_04802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10226_ (.A1_N(_07522_),
    .A2_N(_07578_),
    .B1(\design_top.MEM[29][20] ),
    .B2(_07580_),
    .X(_04801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10227_ (.A1_N(_07523_),
    .A2_N(_07578_),
    .B1(\design_top.MEM[29][19] ),
    .B2(_07580_),
    .X(_04800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10228_ (.A1_N(_07524_),
    .A2_N(_07577_),
    .B1(\design_top.MEM[29][18] ),
    .B2(_07579_),
    .X(_04799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10229_ (.A1_N(_07525_),
    .A2_N(_07577_),
    .B1(\design_top.MEM[29][17] ),
    .B2(_07579_),
    .X(_04798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10230_ (.A1_N(_07526_),
    .A2_N(_07577_),
    .B1(\design_top.MEM[29][16] ),
    .B2(_07579_),
    .X(_04797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10231_ (.A(_07502_),
    .B(_07568_),
    .X(_07581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10232_ (.A(_07581_),
    .X(_07582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10233_ (.A1(_06865_),
    .A2(_07067_),
    .B1(_07581_),
    .X(_07583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10234_ (.A(_07583_),
    .X(_07584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10235_ (.A1_N(_07527_),
    .A2_N(_07582_),
    .B1(\design_top.MEM[29][31] ),
    .B2(_07584_),
    .X(_04796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10236_ (.A1_N(_07507_),
    .A2_N(_07582_),
    .B1(\design_top.MEM[29][30] ),
    .B2(_07584_),
    .X(_04795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10237_ (.A1_N(_07508_),
    .A2_N(_07582_),
    .B1(\design_top.MEM[29][29] ),
    .B2(_07584_),
    .X(_04794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10238_ (.A1_N(_07509_),
    .A2_N(_07582_),
    .B1(\design_top.MEM[29][28] ),
    .B2(_07584_),
    .X(_04793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10239_ (.A1_N(_07510_),
    .A2_N(_07582_),
    .B1(\design_top.MEM[29][27] ),
    .B2(_07584_),
    .X(_04792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10240_ (.A1_N(_07511_),
    .A2_N(_07581_),
    .B1(\design_top.MEM[29][26] ),
    .B2(_07583_),
    .X(_04791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10241_ (.A1_N(_07512_),
    .A2_N(_07581_),
    .B1(\design_top.MEM[29][25] ),
    .B2(_07583_),
    .X(_04790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10242_ (.A1_N(_07513_),
    .A2_N(_07581_),
    .B1(\design_top.MEM[29][24] ),
    .B2(_07583_),
    .X(_04789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10243_ (.A(_07533_),
    .B(_07052_),
    .X(_07585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10244_ (.A(_07585_),
    .X(_07586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10245_ (.A1(_07055_),
    .A2(_07039_),
    .B1(_07585_),
    .X(_07587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10246_ (.A(_07587_),
    .X(_07588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10247_ (.A1_N(_07532_),
    .A2_N(_07586_),
    .B1(\design_top.MEM[2][15] ),
    .B2(_07588_),
    .X(_04788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10248_ (.A1_N(_07539_),
    .A2_N(_07586_),
    .B1(\design_top.MEM[2][14] ),
    .B2(_07588_),
    .X(_04787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10249_ (.A1_N(_07540_),
    .A2_N(_07586_),
    .B1(\design_top.MEM[2][13] ),
    .B2(_07588_),
    .X(_04786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10250_ (.A1_N(_07541_),
    .A2_N(_07586_),
    .B1(\design_top.MEM[2][12] ),
    .B2(_07588_),
    .X(_04785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10251_ (.A1_N(_07542_),
    .A2_N(_07586_),
    .B1(\design_top.MEM[2][11] ),
    .B2(_07588_),
    .X(_04784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10252_ (.A1_N(_07543_),
    .A2_N(_07585_),
    .B1(\design_top.MEM[2][10] ),
    .B2(_07587_),
    .X(_04783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10253_ (.A1_N(_07544_),
    .A2_N(_07585_),
    .B1(\design_top.MEM[2][9] ),
    .B2(_07587_),
    .X(_04782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10254_ (.A1_N(_07545_),
    .A2_N(_07585_),
    .B1(\design_top.MEM[2][8] ),
    .B2(_07587_),
    .X(_04781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10255_ (.A(_07515_),
    .B(_07052_),
    .X(_07589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10256_ (.A(_07589_),
    .X(_07590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10257_ (.A1(_06905_),
    .A2(_07039_),
    .B1(_07589_),
    .X(_07591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10258_ (.A(_07591_),
    .X(_07592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10259_ (.A1_N(_07514_),
    .A2_N(_07590_),
    .B1(\design_top.MEM[2][23] ),
    .B2(_07592_),
    .X(_04780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10260_ (.A1_N(_07520_),
    .A2_N(_07590_),
    .B1(\design_top.MEM[2][22] ),
    .B2(_07592_),
    .X(_04779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10261_ (.A1_N(_07521_),
    .A2_N(_07590_),
    .B1(\design_top.MEM[2][21] ),
    .B2(_07592_),
    .X(_04778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10262_ (.A1_N(_07522_),
    .A2_N(_07590_),
    .B1(\design_top.MEM[2][20] ),
    .B2(_07592_),
    .X(_04777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10263_ (.A1_N(_07523_),
    .A2_N(_07590_),
    .B1(\design_top.MEM[2][19] ),
    .B2(_07592_),
    .X(_04776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10264_ (.A1_N(_07524_),
    .A2_N(_07589_),
    .B1(\design_top.MEM[2][18] ),
    .B2(_07591_),
    .X(_04775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10265_ (.A1_N(_07525_),
    .A2_N(_07589_),
    .B1(\design_top.MEM[2][17] ),
    .B2(_07591_),
    .X(_04774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10266_ (.A1_N(_07526_),
    .A2_N(_07589_),
    .B1(\design_top.MEM[2][16] ),
    .B2(_07591_),
    .X(_04773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10267_ (.A(_06912_),
    .B(_07179_),
    .X(_07593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10268_ (.A(_07593_),
    .X(_07594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10269_ (.A1(_06865_),
    .A2(_07221_),
    .B1(_07593_),
    .X(_07595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10270_ (.A(_07595_),
    .X(_07596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10271_ (.A1_N(_06909_),
    .A2_N(_07594_),
    .B1(\design_top.MEM[13][15] ),
    .B2(_07596_),
    .X(_04772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10272_ (.A1_N(_06919_),
    .A2_N(_07594_),
    .B1(\design_top.MEM[13][14] ),
    .B2(_07596_),
    .X(_04771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10273_ (.A1_N(_06922_),
    .A2_N(_07594_),
    .B1(\design_top.MEM[13][13] ),
    .B2(_07596_),
    .X(_04770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10274_ (.A1_N(_06925_),
    .A2_N(_07594_),
    .B1(\design_top.MEM[13][12] ),
    .B2(_07596_),
    .X(_04769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10275_ (.A1_N(_06928_),
    .A2_N(_07594_),
    .B1(\design_top.MEM[13][11] ),
    .B2(_07596_),
    .X(_04768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10276_ (.A1_N(_06931_),
    .A2_N(_07593_),
    .B1(\design_top.MEM[13][10] ),
    .B2(_07595_),
    .X(_04767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10277_ (.A1_N(_06934_),
    .A2_N(_07593_),
    .B1(\design_top.MEM[13][9] ),
    .B2(_07595_),
    .X(_04766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10278_ (.A1_N(_06937_),
    .A2_N(_07593_),
    .B1(\design_top.MEM[13][8] ),
    .B2(_07595_),
    .X(_04765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10279_ (.A(_06943_),
    .B(_07044_),
    .X(_07597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10280_ (.A(_07597_),
    .X(_07598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10281_ (.A1(_06870_),
    .A2(_07083_),
    .B1(_07597_),
    .X(_07599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10282_ (.A(_07599_),
    .X(_07600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10283_ (.A1_N(_06940_),
    .A2_N(_07598_),
    .B1(\design_top.MEM[11][23] ),
    .B2(_07600_),
    .X(_04764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10284_ (.A1_N(_06950_),
    .A2_N(_07598_),
    .B1(\design_top.MEM[11][22] ),
    .B2(_07600_),
    .X(_04763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10285_ (.A1_N(_06953_),
    .A2_N(_07598_),
    .B1(\design_top.MEM[11][21] ),
    .B2(_07600_),
    .X(_04762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10286_ (.A1_N(_06956_),
    .A2_N(_07598_),
    .B1(\design_top.MEM[11][20] ),
    .B2(_07600_),
    .X(_04761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10287_ (.A1_N(_06959_),
    .A2_N(_07598_),
    .B1(\design_top.MEM[11][19] ),
    .B2(_07600_),
    .X(_04760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10288_ (.A1_N(_06962_),
    .A2_N(_07597_),
    .B1(\design_top.MEM[11][18] ),
    .B2(_07599_),
    .X(_04759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10289_ (.A1_N(_06965_),
    .A2_N(_07597_),
    .B1(\design_top.MEM[11][17] ),
    .B2(_07599_),
    .X(_04758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10290_ (.A1_N(_06968_),
    .A2_N(_07597_),
    .B1(\design_top.MEM[11][16] ),
    .B2(_07599_),
    .X(_04757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _10291_ (.A1(_00802_),
    .A2(_06782_),
    .A3(_06981_),
    .B1(_06783_),
    .B2(_06784_),
    .X(_07601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10292_ (.A(_06982_),
    .B(_07601_),
    .X(_01381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _10293_ (.A(_07042_),
    .B(_01381_),
    .C(_06987_),
    .X(_07602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10294_ (.A(_07602_),
    .Y(_07603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10295_ (.A(_07603_),
    .X(_07604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10296_ (.A(_07604_),
    .X(_07605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10297_ (.A(_07602_),
    .X(_07606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10298_ (.A1(\design_top.IOMUX[3][31] ),
    .A2(_07605_),
    .B1(\design_top.DATAO[31] ),
    .B2(_07606_),
    .C1(_07032_),
    .X(_04756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10299_ (.A(_07604_),
    .X(_07607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10300_ (.A(_07602_),
    .X(_07608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10301_ (.A(_07608_),
    .X(_07609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10302_ (.A1(\design_top.IOMUX[3][30] ),
    .A2(_07607_),
    .B1(\design_top.DATAO[30] ),
    .B2(_07609_),
    .C1(_07032_),
    .X(_04755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10303_ (.A1(\design_top.IOMUX[3][29] ),
    .A2(_07607_),
    .B1(\design_top.DATAO[29] ),
    .B2(_07609_),
    .C1(_07032_),
    .X(_04754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10304_ (.A1(\design_top.IOMUX[3][28] ),
    .A2(_07607_),
    .B1(\design_top.DATAO[28] ),
    .B2(_07609_),
    .C1(_07032_),
    .X(_04753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10305_ (.A(_07031_),
    .X(_07610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10306_ (.A1(\design_top.IOMUX[3][27] ),
    .A2(_07607_),
    .B1(\design_top.DATAO[27] ),
    .B2(_07609_),
    .C1(_07610_),
    .X(_04752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10307_ (.A1(\design_top.IOMUX[3][26] ),
    .A2(_07607_),
    .B1(\design_top.DATAO[26] ),
    .B2(_07609_),
    .C1(_07610_),
    .X(_04751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10308_ (.A(_07604_),
    .X(_07611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10309_ (.A(_07608_),
    .X(_07612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10310_ (.A1(\design_top.IOMUX[3][25] ),
    .A2(_07611_),
    .B1(\design_top.DATAO[25] ),
    .B2(_07612_),
    .C1(_07610_),
    .X(_04750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10311_ (.A1(\design_top.IOMUX[3][24] ),
    .A2(_07611_),
    .B1(\design_top.DATAO[24] ),
    .B2(_07612_),
    .C1(_07610_),
    .X(_04749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10312_ (.A1(\design_top.IOMUX[3][23] ),
    .A2(_07611_),
    .B1(\design_top.DATAO[23] ),
    .B2(_07612_),
    .C1(_07610_),
    .X(_04748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10313_ (.A(_07031_),
    .X(_07613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10314_ (.A1(\design_top.IOMUX[3][22] ),
    .A2(_07611_),
    .B1(\design_top.DATAO[22] ),
    .B2(_07612_),
    .C1(_07613_),
    .X(_04747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10315_ (.A1(\design_top.IOMUX[3][21] ),
    .A2(_07611_),
    .B1(\design_top.DATAO[21] ),
    .B2(_07612_),
    .C1(_07613_),
    .X(_04746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10316_ (.A(_07603_),
    .X(_07614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10317_ (.A(_07608_),
    .X(_07615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10318_ (.A1(\design_top.IOMUX[3][20] ),
    .A2(_07614_),
    .B1(\design_top.DATAO[20] ),
    .B2(_07615_),
    .C1(_07613_),
    .X(_04745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10319_ (.A1(\design_top.IOMUX[3][19] ),
    .A2(_07614_),
    .B1(\design_top.DATAO[19] ),
    .B2(_07615_),
    .C1(_07613_),
    .X(_04744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10320_ (.A1(\design_top.IOMUX[3][18] ),
    .A2(_07614_),
    .B1(\design_top.DATAO[18] ),
    .B2(_07615_),
    .C1(_07613_),
    .X(_04743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10321_ (.A(_06991_),
    .X(_07616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10322_ (.A1(\design_top.IOMUX[3][17] ),
    .A2(_07614_),
    .B1(\design_top.DATAO[17] ),
    .B2(_07615_),
    .C1(_07616_),
    .X(_04742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10323_ (.A1(\design_top.IOMUX[3][16] ),
    .A2(_07614_),
    .B1(\design_top.DATAO[16] ),
    .B2(_07615_),
    .C1(_07616_),
    .X(_04741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10324_ (.A(_07603_),
    .X(_07617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10325_ (.A(_07602_),
    .X(_07618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10326_ (.A1(\design_top.IOMUX[3][15] ),
    .A2(_07617_),
    .B1(\design_top.DATAO[15] ),
    .B2(_07618_),
    .C1(_07616_),
    .X(_04740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10327_ (.A1(\design_top.IOMUX[3][14] ),
    .A2(_07617_),
    .B1(\design_top.DATAO[14] ),
    .B2(_07618_),
    .C1(_07616_),
    .X(_04739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10328_ (.A1(\design_top.IOMUX[3][13] ),
    .A2(_07617_),
    .B1(\design_top.DATAO[13] ),
    .B2(_07618_),
    .C1(_07616_),
    .X(_04738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10329_ (.A(_06991_),
    .X(_07619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10330_ (.A1(\design_top.IOMUX[3][12] ),
    .A2(_07617_),
    .B1(\design_top.DATAO[12] ),
    .B2(_07618_),
    .C1(_07619_),
    .X(_04737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10331_ (.A1(\design_top.IOMUX[3][11] ),
    .A2(_07617_),
    .B1(\design_top.DATAO[11] ),
    .B2(_07618_),
    .C1(_07619_),
    .X(_04736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10332_ (.A(_07603_),
    .X(_07620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10333_ (.A(_07602_),
    .X(_07621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10334_ (.A1(\design_top.IOMUX[3][10] ),
    .A2(_07620_),
    .B1(\design_top.DATAO[10] ),
    .B2(_07621_),
    .C1(_07619_),
    .X(_04735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10335_ (.A1(\design_top.IOMUX[3][9] ),
    .A2(_07620_),
    .B1(\design_top.DATAO[9] ),
    .B2(_07621_),
    .C1(_07619_),
    .X(_04734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10336_ (.A1(\design_top.IOMUX[3][8] ),
    .A2(_07620_),
    .B1(\design_top.DATAO[8] ),
    .B2(_07621_),
    .C1(_07619_),
    .X(_04733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10337_ (.A(_06991_),
    .X(_07622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10338_ (.A1(\design_top.IOMUX[3][7] ),
    .A2(_07620_),
    .B1(\design_top.DATAO[7] ),
    .B2(_07621_),
    .C1(_07622_),
    .X(_04732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10339_ (.A(\design_top.IRES[7] ),
    .X(_07623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10340_ (.A(_07623_),
    .X(_07624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a221o_2 _10341_ (.A1(\design_top.DATAO[6] ),
    .A2(_07605_),
    .B1(\design_top.IOMUX[3][6] ),
    .B2(_07606_),
    .C1(_07624_),
    .X(_04731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a221o_2 _10342_ (.A1(\design_top.DATAO[5] ),
    .A2(_07605_),
    .B1(\design_top.IOMUX[3][5] ),
    .B2(_07606_),
    .C1(_07624_),
    .X(_04730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10343_ (.A1(\design_top.IOMUX[3][4] ),
    .A2(_07620_),
    .B1(\design_top.DATAO[4] ),
    .B2(_07621_),
    .C1(_07622_),
    .X(_04729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10344_ (.A1(\design_top.IOMUX[3][3] ),
    .A2(_07604_),
    .B1(\design_top.DATAO[3] ),
    .B2(_07608_),
    .C1(_07622_),
    .X(_04728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10345_ (.A1(\design_top.IOMUX[3][2] ),
    .A2(_07604_),
    .B1(\design_top.DATAO[2] ),
    .B2(_07608_),
    .C1(_07622_),
    .X(_04727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a221o_2 _10346_ (.A1(\design_top.DATAO[1] ),
    .A2(_07605_),
    .B1(\design_top.IOMUX[3][1] ),
    .B2(_07606_),
    .C1(_07623_),
    .X(_04726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a221o_2 _10347_ (.A1(\design_top.DATAO[0] ),
    .A2(_07605_),
    .B1(\design_top.IOMUX[3][0] ),
    .B2(_07606_),
    .C1(_07623_),
    .X(_04725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10348_ (.A(_06845_),
    .B(_07044_),
    .X(_07625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10349_ (.A(_07625_),
    .X(_07626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10350_ (.A1(_06870_),
    .A2(_07083_),
    .B1(_07625_),
    .X(_07627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10351_ (.A(_07627_),
    .X(_07628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10352_ (.A1_N(_07527_),
    .A2_N(_07626_),
    .B1(\design_top.MEM[11][31] ),
    .B2(_07628_),
    .X(_04724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10353_ (.A1_N(_06656_),
    .A2_N(_07626_),
    .B1(\design_top.MEM[11][30] ),
    .B2(_07628_),
    .X(_04723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10354_ (.A1_N(_06874_),
    .A2_N(_07626_),
    .B1(\design_top.MEM[11][29] ),
    .B2(_07628_),
    .X(_04722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10355_ (.A1_N(_06877_),
    .A2_N(_07626_),
    .B1(\design_top.MEM[11][28] ),
    .B2(_07628_),
    .X(_04721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10356_ (.A1_N(_06880_),
    .A2_N(_07626_),
    .B1(\design_top.MEM[11][27] ),
    .B2(_07628_),
    .X(_04720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10357_ (.A1_N(_06883_),
    .A2_N(_07625_),
    .B1(\design_top.MEM[11][26] ),
    .B2(_07627_),
    .X(_04719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10358_ (.A1_N(_06886_),
    .A2_N(_07625_),
    .B1(\design_top.MEM[11][25] ),
    .B2(_07627_),
    .X(_04718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10359_ (.A1_N(_06889_),
    .A2_N(_07625_),
    .B1(\design_top.MEM[11][24] ),
    .B2(_07627_),
    .X(_04717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10360_ (.A(_06894_),
    .B(_07178_),
    .X(_07629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10361_ (.A(_06912_),
    .B(_07629_),
    .X(_07630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10362_ (.A(_07630_),
    .X(_07631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10363_ (.A1(_07557_),
    .A2(_07221_),
    .B1(_07630_),
    .X(_07632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10364_ (.A(_07632_),
    .X(_07633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10365_ (.A1_N(_06909_),
    .A2_N(_07631_),
    .B1(\design_top.MEM[12][15] ),
    .B2(_07633_),
    .X(_04716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10366_ (.A1_N(_06919_),
    .A2_N(_07631_),
    .B1(\design_top.MEM[12][14] ),
    .B2(_07633_),
    .X(_04715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10367_ (.A1_N(_06922_),
    .A2_N(_07631_),
    .B1(\design_top.MEM[12][13] ),
    .B2(_07633_),
    .X(_04714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10368_ (.A1_N(_06925_),
    .A2_N(_07631_),
    .B1(\design_top.MEM[12][12] ),
    .B2(_07633_),
    .X(_04713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10369_ (.A1_N(_06928_),
    .A2_N(_07631_),
    .B1(\design_top.MEM[12][11] ),
    .B2(_07633_),
    .X(_04712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10370_ (.A1_N(_06931_),
    .A2_N(_07630_),
    .B1(\design_top.MEM[12][10] ),
    .B2(_07632_),
    .X(_04711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10371_ (.A1_N(_06934_),
    .A2_N(_07630_),
    .B1(\design_top.MEM[12][9] ),
    .B2(_07632_),
    .X(_04710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10372_ (.A1_N(_06937_),
    .A2_N(_07630_),
    .B1(\design_top.MEM[12][8] ),
    .B2(_07632_),
    .X(_04709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10373_ (.A(_06845_),
    .B(_07629_),
    .X(_07634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10374_ (.A(_07634_),
    .X(_07635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10375_ (.A1(_07557_),
    .A2(_07183_),
    .B1(_07634_),
    .X(_07636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10376_ (.A(_07636_),
    .X(_07637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10377_ (.A1_N(_06892_),
    .A2_N(_07635_),
    .B1(\design_top.MEM[12][31] ),
    .B2(_07637_),
    .X(_04708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10378_ (.A1_N(_06656_),
    .A2_N(_07635_),
    .B1(\design_top.MEM[12][30] ),
    .B2(_07637_),
    .X(_04707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10379_ (.A1_N(_06874_),
    .A2_N(_07635_),
    .B1(\design_top.MEM[12][29] ),
    .B2(_07637_),
    .X(_04706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10380_ (.A1_N(_06877_),
    .A2_N(_07635_),
    .B1(\design_top.MEM[12][28] ),
    .B2(_07637_),
    .X(_04705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10381_ (.A1_N(_06880_),
    .A2_N(_07635_),
    .B1(\design_top.MEM[12][27] ),
    .B2(_07637_),
    .X(_04704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10382_ (.A1_N(_06883_),
    .A2_N(_07634_),
    .B1(\design_top.MEM[12][26] ),
    .B2(_07636_),
    .X(_04703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10383_ (.A1_N(_06886_),
    .A2_N(_07634_),
    .B1(\design_top.MEM[12][25] ),
    .B2(_07636_),
    .X(_04702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10384_ (.A1_N(_06889_),
    .A2_N(_07634_),
    .B1(\design_top.MEM[12][24] ),
    .B2(_07636_),
    .X(_04701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10385_ (.A(\design_top.core0.XRES ),
    .X(_07638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10386_ (.A(_07638_),
    .X(_07639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10387_ (.A(\design_top.IDATA[31] ),
    .Y(_07640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10388_ (.A(_06662_),
    .X(_07641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10389_ (.A(_07641_),
    .X(_07642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10390_ (.A(_01420_),
    .Y(_07643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _10391_ (.A(_01421_),
    .B(_07643_),
    .C(_01422_),
    .X(_07644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10392_ (.A(io_out[21]),
    .B(io_out[20]),
    .Y(_07645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _10393_ (.A(io_out[23]),
    .B(_07645_),
    .C_N(io_out[22]),
    .X(_07646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10394_ (.A(_07644_),
    .B(_07646_),
    .Y(_07647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10395_ (.A(_01421_),
    .Y(_07648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _10396_ (.A(_07648_),
    .B(_07643_),
    .C(_01422_),
    .X(_07649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10397_ (.A(_07646_),
    .B(_07649_),
    .Y(_07650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10398_ (.A(_07647_),
    .B(_07650_),
    .X(_07651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10399_ (.A(_07651_),
    .Y(_07652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10400_ (.A(_07652_),
    .X(_00643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10401_ (.A(\design_top.core0.UIMM[31] ),
    .Y(_07653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10402_ (.A(_06661_),
    .X(_07654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10403_ (.A(_07654_),
    .X(_07655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10404_ (.A(_07655_),
    .X(_07656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _10405_ (.A1(_07640_),
    .A2(_07642_),
    .A3(_00643_),
    .B1(_07653_),
    .B2(_07656_),
    .X(_07657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10406_ (.A(_07639_),
    .B(_07657_),
    .Y(_04700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10407_ (.A(_06662_),
    .X(_07658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10408_ (.A(_07658_),
    .X(_07659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10409_ (.A(_07659_),
    .X(_07660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10410_ (.A(_07660_),
    .X(\design_top.HLT ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10411_ (.A(\design_top.IDATA[30] ),
    .Y(_07661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10412_ (.A(\design_top.core0.UIMM[30] ),
    .Y(_07662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10413_ (.A(_07655_),
    .X(_07663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _10414_ (.A1(_07661_),
    .A2(_07642_),
    .A3(_00643_),
    .B1(_07662_),
    .B2(_07663_),
    .X(_07664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10415_ (.A(_07639_),
    .B(_07664_),
    .Y(_04699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10416_ (.A(_07659_),
    .X(_07665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10417_ (.A(_00701_),
    .Y(_07666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10418_ (.A(_06662_),
    .B(_07652_),
    .X(_07667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10419_ (.A(_07667_),
    .X(_07668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _10420_ (.A1_N(\design_top.core0.UIMM[29] ),
    .A2_N(_07665_),
    .B1(_07666_),
    .B2(_07668_),
    .X(_07669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10421_ (.A(_07639_),
    .B(_07669_),
    .Y(_04698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10422_ (.A(_00697_),
    .Y(_07670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _10423_ (.A1_N(\design_top.core0.UIMM[28] ),
    .A2_N(_07665_),
    .B1(_07670_),
    .B2(_07668_),
    .X(_07671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10424_ (.A(_07639_),
    .B(_07671_),
    .Y(_04697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10425_ (.A(_00693_),
    .Y(_07672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _10426_ (.A1_N(\design_top.core0.UIMM[27] ),
    .A2_N(_07665_),
    .B1(_07672_),
    .B2(_07668_),
    .X(_07673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10427_ (.A(_07639_),
    .B(_07673_),
    .Y(_04696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10428_ (.A(_07638_),
    .X(_07674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10429_ (.A(_07658_),
    .X(_07675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10430_ (.A(_07675_),
    .X(_07676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10431_ (.A(_00689_),
    .Y(_07677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _10432_ (.A1_N(\design_top.core0.UIMM[26] ),
    .A2_N(_07676_),
    .B1(_07677_),
    .B2(_07668_),
    .X(_07678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10433_ (.A(_07674_),
    .B(_07678_),
    .Y(_04695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10434_ (.A(_00685_),
    .Y(_07679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _10435_ (.A1_N(\design_top.core0.UIMM[25] ),
    .A2_N(_07676_),
    .B1(_07679_),
    .B2(_07668_),
    .X(_07680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10436_ (.A(_07674_),
    .B(_07680_),
    .Y(_04694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10437_ (.A(_00681_),
    .Y(_07681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _10438_ (.A1_N(\design_top.core0.UIMM[24] ),
    .A2_N(_07676_),
    .B1(_07681_),
    .B2(_07667_),
    .X(_07682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10439_ (.A(_07674_),
    .B(_07682_),
    .Y(_04693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10440_ (.A(\design_top.IDATA[23] ),
    .Y(_07683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10441_ (.A(\design_top.core0.UIMM[23] ),
    .Y(_07684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _10442_ (.A1(_07683_),
    .A2(_07642_),
    .A3(_00643_),
    .B1(_07684_),
    .B2(_07663_),
    .X(_07685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10443_ (.A(_07674_),
    .B(_07685_),
    .Y(_04692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10444_ (.A(\design_top.IDATA[22] ),
    .Y(_07686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10445_ (.A(_07641_),
    .X(_07687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10446_ (.A(\design_top.core0.UIMM[22] ),
    .Y(_07688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _10447_ (.A1(_07686_),
    .A2(_07687_),
    .A3(_07652_),
    .B1(_07688_),
    .B2(_07663_),
    .X(_07689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10448_ (.A(_07674_),
    .B(_07689_),
    .Y(_04691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10449_ (.A(_07638_),
    .X(_07690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10450_ (.A(\design_top.IDATA[21] ),
    .Y(_07691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10451_ (.A(\design_top.core0.UIMM[21] ),
    .Y(_07692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _10452_ (.A1(_07691_),
    .A2(_07687_),
    .A3(_07652_),
    .B1(_07692_),
    .B2(_07663_),
    .X(_07693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10453_ (.A(_07690_),
    .B(_07693_),
    .Y(_04690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10454_ (.A(_00761_),
    .Y(_07694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _10455_ (.A(io_out[23]),
    .B(io_out[22]),
    .C(_07645_),
    .X(_07695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31ai_2 _10456_ (.A1(_07648_),
    .A2(_01420_),
    .A3(_07695_),
    .B1(_07654_),
    .Y(_07696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10457_ (.A(_07696_),
    .X(_07697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _10458_ (.A1_N(\design_top.core0.UIMM[20] ),
    .A2_N(_07676_),
    .B1(_07694_),
    .B2(_07697_),
    .X(_07698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10459_ (.A(_07690_),
    .B(_07698_),
    .Y(_04689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10460_ (.A(_00759_),
    .Y(_07699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _10461_ (.A1_N(\design_top.core0.UIMM[19] ),
    .A2_N(_07676_),
    .B1(_07699_),
    .B2(_07697_),
    .X(_07700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10462_ (.A(_07690_),
    .B(_07700_),
    .Y(_04688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10463_ (.A(_07675_),
    .X(_07701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10464_ (.A(_00757_),
    .Y(_07702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _10465_ (.A1_N(\design_top.core0.UIMM[18] ),
    .A2_N(_07701_),
    .B1(_07702_),
    .B2(_07697_),
    .X(_07703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10466_ (.A(_07690_),
    .B(_07703_),
    .Y(_04687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10467_ (.A(_00755_),
    .Y(_07704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _10468_ (.A1_N(\design_top.core0.UIMM[17] ),
    .A2_N(_07701_),
    .B1(_07704_),
    .B2(_07697_),
    .X(_07705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10469_ (.A(_07690_),
    .B(_07705_),
    .Y(_04686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10470_ (.A(_07638_),
    .X(_07706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10471_ (.A(_00753_),
    .Y(_07707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _10472_ (.A1_N(\design_top.core0.UIMM[16] ),
    .A2_N(_07701_),
    .B1(_07707_),
    .B2(_07697_),
    .X(_07708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10473_ (.A(_07706_),
    .B(_07708_),
    .Y(_04685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10474_ (.A(_00751_),
    .Y(_07709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _10475_ (.A1_N(\design_top.core0.UIMM[15] ),
    .A2_N(_07701_),
    .B1(_07709_),
    .B2(_07696_),
    .X(_07710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10476_ (.A(_07706_),
    .B(_07710_),
    .Y(_04684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10477_ (.A(_00749_),
    .Y(_07711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _10478_ (.A1_N(\design_top.core0.UIMM[14] ),
    .A2_N(_07701_),
    .B1(_07711_),
    .B2(_07696_),
    .X(_07712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10479_ (.A(_07706_),
    .B(_07712_),
    .Y(_04683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10480_ (.A(_00747_),
    .Y(_07713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _10481_ (.A1_N(\design_top.core0.UIMM[13] ),
    .A2_N(_07660_),
    .B1(_07713_),
    .B2(_07696_),
    .X(_07714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10482_ (.A(_07706_),
    .B(_07714_),
    .Y(_04682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10483_ (.A(_00745_),
    .Y(_07715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10484_ (.A(_01422_),
    .Y(_07716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and4b_2 _10485_ (.A_N(_07695_),
    .B(_07643_),
    .C(_07716_),
    .D(_01421_),
    .X(_00010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10486_ (.A(_07658_),
    .B(_00010_),
    .X(_07717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _10487_ (.A1_N(\design_top.core0.UIMM[12] ),
    .A2_N(_07660_),
    .B1(_07715_),
    .B2(_07717_),
    .X(_07718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10488_ (.A(_07706_),
    .B(_07718_),
    .Y(_04681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10489_ (.A(_07687_),
    .X(_07719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10490_ (.A(_07655_),
    .X(_07720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10491_ (.A(\design_top.core0.XRES ),
    .Y(_07721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10492_ (.A(_07721_),
    .X(_07722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10493_ (.A(_07722_),
    .X(_07723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10494_ (.A1(_00049_),
    .A2(_07719_),
    .B1(\design_top.core0.SIMM[11] ),
    .B2(_07720_),
    .C1(_07723_),
    .X(_04680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10495_ (.A(_07722_),
    .X(_07724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10496_ (.A(_07724_),
    .X(_07725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10497_ (.A1(_00048_),
    .A2(_07719_),
    .B1(\design_top.core0.SIMM[10] ),
    .B2(_07720_),
    .C1(_07725_),
    .X(_04679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10498_ (.A(_07654_),
    .X(_07726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10499_ (.A(_07726_),
    .X(_07727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10500_ (.A(_07727_),
    .X(_07728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10501_ (.A1(_00077_),
    .A2(_07719_),
    .B1(_06748_),
    .B2(_07728_),
    .C1(_07725_),
    .X(_04678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10502_ (.A1(_00076_),
    .A2(_07719_),
    .B1(_06750_),
    .B2(_07728_),
    .C1(_07725_),
    .X(_04677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10503_ (.A(_07687_),
    .X(_07729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10504_ (.A1(_00075_),
    .A2(_07729_),
    .B1(_06763_),
    .B2(_07728_),
    .C1(_07725_),
    .X(_04676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10505_ (.A1(_00074_),
    .A2(_07729_),
    .B1(_06760_),
    .B2(_07728_),
    .C1(_07725_),
    .X(_04675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10506_ (.A(_07724_),
    .X(_07730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10507_ (.A1(_00073_),
    .A2(_07729_),
    .B1(_06767_),
    .B2(_07728_),
    .C1(_07730_),
    .X(_04674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10508_ (.A(_07727_),
    .X(_07731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10509_ (.A1(_00072_),
    .A2(_07729_),
    .B1(_06853_),
    .B2(_07731_),
    .C1(_07730_),
    .X(_04673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10510_ (.A1(_00071_),
    .A2(_07729_),
    .B1(_06847_),
    .B2(_07731_),
    .C1(_07730_),
    .X(_04672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10511_ (.A(_07641_),
    .X(_07732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10512_ (.A(_07732_),
    .X(_07733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10513_ (.A1(_00069_),
    .A2(_07733_),
    .B1(_06792_),
    .B2(_07731_),
    .C1(_07730_),
    .X(_04671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10514_ (.A1(_00058_),
    .A2(_07733_),
    .B1(_06780_),
    .B2(_07731_),
    .C1(_07730_),
    .X(_04670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10515_ (.A(_07724_),
    .X(_07734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10516_ (.A1(_00047_),
    .A2(_07733_),
    .B1(\design_top.core0.SIMM[0] ),
    .B2(_07731_),
    .C1(_07734_),
    .X(_04669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10517_ (.A(_07638_),
    .X(_07735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10518_ (.A1(_07640_),
    .A2(_07660_),
    .B1(_00763_),
    .B2(_07656_),
    .X(_07736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10519_ (.A(_07735_),
    .B(_07736_),
    .Y(_04668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10520_ (.A(_07727_),
    .X(_07737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10521_ (.A1(_00070_),
    .A2(_07733_),
    .B1(\design_top.core0.SIMM[30] ),
    .B2(_07737_),
    .C1(_07734_),
    .X(_04667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10522_ (.A1(_00068_),
    .A2(_07733_),
    .B1(_06668_),
    .B2(_07737_),
    .C1(_07734_),
    .X(_04666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10523_ (.A(_07732_),
    .X(_07738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10524_ (.A1(_00067_),
    .A2(_07738_),
    .B1(_06674_),
    .B2(_07737_),
    .C1(_07734_),
    .X(_04665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10525_ (.A1(_00066_),
    .A2(_07738_),
    .B1(\design_top.core0.SIMM[27] ),
    .B2(_07737_),
    .C1(_07734_),
    .X(_04664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10526_ (.A(_07724_),
    .X(_07739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10527_ (.A1(_00065_),
    .A2(_07738_),
    .B1(\design_top.core0.SIMM[26] ),
    .B2(_07737_),
    .C1(_07739_),
    .X(_04663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10528_ (.A(_07654_),
    .X(_07740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10529_ (.A(_07740_),
    .X(_07741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10530_ (.A1(_00064_),
    .A2(_07738_),
    .B1(_06683_),
    .B2(_07741_),
    .C1(_07739_),
    .X(_04662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10531_ (.A1(_00063_),
    .A2(_07738_),
    .B1(_06685_),
    .B2(_07741_),
    .C1(_07739_),
    .X(_04661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10532_ (.A(_07732_),
    .X(_07742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10533_ (.A(\design_top.core0.SIMM[23] ),
    .X(_07743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10534_ (.A1(_00062_),
    .A2(_07742_),
    .B1(_07743_),
    .B2(_07741_),
    .C1(_07739_),
    .X(_04660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10535_ (.A1(_00061_),
    .A2(_07742_),
    .B1(_06699_),
    .B2(_07741_),
    .C1(_07739_),
    .X(_04659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10536_ (.A(_07724_),
    .X(_07744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10537_ (.A1(_00060_),
    .A2(_07742_),
    .B1(_06820_),
    .B2(_07741_),
    .C1(_07744_),
    .X(_04658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10538_ (.A(_07740_),
    .X(_07745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10539_ (.A1(_00059_),
    .A2(_07742_),
    .B1(_06690_),
    .B2(_07745_),
    .C1(_07744_),
    .X(_04657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10540_ (.A1(_00057_),
    .A2(_07742_),
    .B1(\design_top.core0.SIMM[19] ),
    .B2(_07745_),
    .C1(_07744_),
    .X(_04656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10541_ (.A(_07732_),
    .X(_07746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10542_ (.A1(_00056_),
    .A2(_07746_),
    .B1(\design_top.core0.SIMM[18] ),
    .B2(_07745_),
    .C1(_07744_),
    .X(_04655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10543_ (.A1(_00055_),
    .A2(_07746_),
    .B1(_06714_),
    .B2(_07745_),
    .C1(_07744_),
    .X(_04654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10544_ (.A(_07722_),
    .X(_07747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10545_ (.A(_07747_),
    .X(_07748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10546_ (.A1(_00054_),
    .A2(_07746_),
    .B1(_06717_),
    .B2(_07745_),
    .C1(_07748_),
    .X(_04653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10547_ (.A(_07740_),
    .X(_07749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10548_ (.A1(_00053_),
    .A2(_07746_),
    .B1(_06808_),
    .B2(_07749_),
    .C1(_07748_),
    .X(_04652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10549_ (.A1(_00052_),
    .A2(_07746_),
    .B1(\design_top.core0.SIMM[14] ),
    .B2(_07749_),
    .C1(_07748_),
    .X(_04651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10550_ (.A(_07732_),
    .X(_07750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10551_ (.A1(_00051_),
    .A2(_07750_),
    .B1(_06730_),
    .B2(_07749_),
    .C1(_07748_),
    .X(_04650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10552_ (.A1(_00050_),
    .A2(_07750_),
    .B1(_06725_),
    .B2(_07749_),
    .C1(_07748_),
    .X(_04649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10553_ (.A(_07641_),
    .X(_07751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10554_ (.A(_07695_),
    .X(_07752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10555_ (.A(\design_top.core0.XRCC ),
    .Y(_07753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _10556_ (.A1(_07751_),
    .A2(_07752_),
    .A3(_07649_),
    .B1(_07753_),
    .B2(_07663_),
    .X(_07754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10557_ (.A(_07735_),
    .B(_07754_),
    .Y(_04648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10558_ (.A(\design_top.core0.XMCC ),
    .Y(_07755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10559_ (.A(_07726_),
    .X(_07756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _10560_ (.A1(_07751_),
    .A2(_07752_),
    .A3(_07644_),
    .B1(_07755_),
    .B2(_07756_),
    .X(_07757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10561_ (.A(_07735_),
    .B(_07757_),
    .Y(_04647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10562_ (.A(_07722_),
    .X(_07758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _10563_ (.A1(\design_top.core0.XSCC ),
    .A2(_07720_),
    .B1(_07758_),
    .C1(_07717_),
    .X(_04646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and4b_2 _10564_ (.A_N(_07752_),
    .B(_07716_),
    .C(_07648_),
    .D(_07643_),
    .X(_07759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10565_ (.A(_07758_),
    .X(_07760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10566_ (.A1(\design_top.HLT ),
    .A2(_07759_),
    .B1(_07760_),
    .X(_04645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _10567_ (.A(_07648_),
    .B(_01420_),
    .C(_07716_),
    .X(_07761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10568_ (.A(\design_top.core0.XBCC ),
    .Y(_07762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _10569_ (.A1(_07751_),
    .A2(_07752_),
    .A3(_07761_),
    .B1(_07762_),
    .B2(_07756_),
    .X(_07763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10570_ (.A(_07735_),
    .B(_07763_),
    .Y(_04644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10571_ (.A(_07752_),
    .B(_07761_),
    .Y(_00009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10572_ (.A(\design_top.core0.XJALR ),
    .Y(_07764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _10573_ (.A1(_07751_),
    .A2(_07761_),
    .A3(_07646_),
    .B1(_07764_),
    .B2(_07756_),
    .X(_07765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10574_ (.A(_07735_),
    .B(_07765_),
    .Y(_04643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10575_ (.A(_07655_),
    .X(_07766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10576_ (.A(_07687_),
    .X(_07767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and4bb_2 _10577_ (.A_N(_07761_),
    .B_N(_07645_),
    .C(io_out[23]),
    .D(io_out[22]),
    .X(_00008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10578_ (.A(_07747_),
    .X(_07768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10579_ (.A1(\design_top.core0.XJAL ),
    .A2(_07766_),
    .B1(_07767_),
    .B2(_00008_),
    .C1(_07768_),
    .X(_04642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10580_ (.A1(\design_top.core0.XAUIPC ),
    .A2(_07766_),
    .B1(_07767_),
    .B2(_07647_),
    .C1(_07768_),
    .X(_04641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10581_ (.A1(\design_top.core0.XLUI ),
    .A2(_07766_),
    .B1(_07719_),
    .B2(_07650_),
    .C1(_07768_),
    .X(_04640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10582_ (.A(\design_top.core0.XRES ),
    .X(_07769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10583_ (.A(\design_top.core0.FCT7[5] ),
    .Y(_07770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10584_ (.A1(_07661_),
    .A2(_07660_),
    .B1(_07770_),
    .B2(_07656_),
    .X(_07771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10585_ (.A(_07769_),
    .B(_07771_),
    .Y(_04639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10586_ (.A(_07675_),
    .X(_07772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22oi_2 _10587_ (.A1(\design_top.IDATA[23] ),
    .A2(_07766_),
    .B1(\design_top.core0.S2PTR[3] ),
    .B2(_07772_),
    .Y(_07773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10588_ (.A(_07769_),
    .B(_07773_),
    .Y(_04638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22oi_2 _10589_ (.A1(\design_top.IDATA[22] ),
    .A2(_07656_),
    .B1(\design_top.core0.S2PTR[2] ),
    .B2(_07665_),
    .Y(_07774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10590_ (.A(_07769_),
    .B(_07774_),
    .Y(_04637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22oi_2 _10591_ (.A1(\design_top.IDATA[21] ),
    .A2(_07656_),
    .B1(\design_top.core0.S2PTR[1] ),
    .B2(_07665_),
    .Y(_07775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10592_ (.A(_07769_),
    .B(_07775_),
    .Y(_04636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10593_ (.A1(\design_top.IDATA[20] ),
    .A2(_07750_),
    .B1(\design_top.core0.S2PTR[0] ),
    .B2(_07749_),
    .C1(_07768_),
    .X(_04635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10594_ (.A(_07740_),
    .X(_07776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10595_ (.A1(\design_top.IDATA[18] ),
    .A2(_07750_),
    .B1(\design_top.core0.S1PTR[3] ),
    .B2(_07776_),
    .C1(_07768_),
    .X(_04634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10596_ (.A(_07747_),
    .X(_07777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10597_ (.A1(\design_top.IDATA[17] ),
    .A2(_07750_),
    .B1(\design_top.core0.S1PTR[2] ),
    .B2(_07776_),
    .C1(_07777_),
    .X(_04633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10598_ (.A(_07641_),
    .X(_07778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10599_ (.A(_07778_),
    .X(_07779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10600_ (.A1(\design_top.IDATA[16] ),
    .A2(_07779_),
    .B1(\design_top.core0.S1PTR[1] ),
    .B2(_07776_),
    .C1(_07777_),
    .X(_04632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10601_ (.A1(\design_top.IDATA[15] ),
    .A2(_07779_),
    .B1(\design_top.core0.S1PTR[0] ),
    .B2(_07776_),
    .C1(_07777_),
    .X(_04631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10602_ (.A1(\design_top.IDATA[14] ),
    .A2(_07779_),
    .B1(\design_top.core0.FCT3[2] ),
    .B2(_07776_),
    .C1(_07777_),
    .X(_04630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10603_ (.A(\design_top.core0.FCT3[1] ),
    .X(_07780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10604_ (.A(_07740_),
    .X(_07781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10605_ (.A1(\design_top.IDATA[13] ),
    .A2(_07779_),
    .B1(_07780_),
    .B2(_07781_),
    .C1(_07777_),
    .X(_04629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10606_ (.A(_07747_),
    .X(_07782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10607_ (.A1(\design_top.IDATA[12] ),
    .A2(_07779_),
    .B1(\design_top.core0.FCT3[0] ),
    .B2(_07781_),
    .C1(_07782_),
    .X(_04628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10608_ (.A(_07778_),
    .X(_07783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10609_ (.A1(\design_top.IDATA[10] ),
    .A2(_07783_),
    .B1(\design_top.core0.XIDATA[10] ),
    .B2(_07781_),
    .C1(_07782_),
    .X(_04627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10610_ (.A1(\design_top.IDATA[9] ),
    .A2(_07783_),
    .B1(\design_top.core0.XIDATA[9] ),
    .B2(_07781_),
    .C1(_07782_),
    .X(_04626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10611_ (.A1(\design_top.IDATA[8] ),
    .A2(_07783_),
    .B1(\design_top.core0.XIDATA[8] ),
    .B2(_07781_),
    .C1(_07782_),
    .X(_04625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10612_ (.A(_07654_),
    .X(_07784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10613_ (.A(_07784_),
    .X(_07785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10614_ (.A1(\design_top.IDATA[7] ),
    .A2(_07783_),
    .B1(\design_top.core0.XIDATA[7] ),
    .B2(_07785_),
    .C1(_07782_),
    .X(_04624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10615_ (.A(_07747_),
    .X(_07786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10616_ (.A1(_00101_),
    .A2(_07783_),
    .B1(\design_top.IADDR[31] ),
    .B2(_07785_),
    .C1(_07786_),
    .X(_04623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10617_ (.A(_07778_),
    .X(_07787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10618_ (.A1(_00100_),
    .A2(_07787_),
    .B1(\design_top.IADDR[30] ),
    .B2(_07785_),
    .C1(_07786_),
    .X(_04622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10619_ (.A1(_00098_),
    .A2(_07787_),
    .B1(\design_top.IADDR[29] ),
    .B2(_07785_),
    .C1(_07786_),
    .X(_04621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10620_ (.A1(_00097_),
    .A2(_07787_),
    .B1(\design_top.IADDR[28] ),
    .B2(_07785_),
    .C1(_07786_),
    .X(_04620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10621_ (.A(_07784_),
    .X(_07788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10622_ (.A1(_00096_),
    .A2(_07787_),
    .B1(\design_top.IADDR[27] ),
    .B2(_07788_),
    .C1(_07786_),
    .X(_04619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10623_ (.A(_07722_),
    .X(_07789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10624_ (.A(_07789_),
    .X(_07790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10625_ (.A1(_00095_),
    .A2(_07787_),
    .B1(\design_top.IADDR[26] ),
    .B2(_07788_),
    .C1(_07790_),
    .X(_04618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10626_ (.A(_07778_),
    .X(_07791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10627_ (.A1(_00094_),
    .A2(_07791_),
    .B1(\design_top.IADDR[25] ),
    .B2(_07788_),
    .C1(_07790_),
    .X(_04617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10628_ (.A1(_00093_),
    .A2(_07791_),
    .B1(\design_top.IADDR[24] ),
    .B2(_07788_),
    .C1(_07790_),
    .X(_04616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10629_ (.A1(_00092_),
    .A2(_07791_),
    .B1(\design_top.IADDR[23] ),
    .B2(_07788_),
    .C1(_07790_),
    .X(_04615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10630_ (.A(_07784_),
    .X(_07792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10631_ (.A1(_00091_),
    .A2(_07791_),
    .B1(\design_top.IADDR[22] ),
    .B2(_07792_),
    .C1(_07790_),
    .X(_04614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10632_ (.A(_07789_),
    .X(_07793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10633_ (.A1(_00090_),
    .A2(_07791_),
    .B1(\design_top.IADDR[21] ),
    .B2(_07792_),
    .C1(_07793_),
    .X(_04613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10634_ (.A(_07778_),
    .X(_07794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10635_ (.A1(_00089_),
    .A2(_07794_),
    .B1(\design_top.IADDR[20] ),
    .B2(_07792_),
    .C1(_07793_),
    .X(_04612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10636_ (.A1(_00088_),
    .A2(_07794_),
    .B1(\design_top.IADDR[19] ),
    .B2(_07792_),
    .C1(_07793_),
    .X(_04611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10637_ (.A1(_00087_),
    .A2(_07794_),
    .B1(\design_top.IADDR[18] ),
    .B2(_07792_),
    .C1(_07793_),
    .X(_04610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10638_ (.A(_07784_),
    .X(_07795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10639_ (.A1(_00086_),
    .A2(_07794_),
    .B1(\design_top.IADDR[17] ),
    .B2(_07795_),
    .C1(_07793_),
    .X(_04609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10640_ (.A(_07789_),
    .X(_07796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10641_ (.A1(_00085_),
    .A2(_07794_),
    .B1(\design_top.IADDR[16] ),
    .B2(_07795_),
    .C1(_07796_),
    .X(_04608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10642_ (.A(_07675_),
    .X(_07797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10643_ (.A1(_00084_),
    .A2(_07797_),
    .B1(\design_top.IADDR[15] ),
    .B2(_07795_),
    .C1(_07796_),
    .X(_04607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10644_ (.A1(_00083_),
    .A2(_07797_),
    .B1(\design_top.IADDR[14] ),
    .B2(_07795_),
    .C1(_07796_),
    .X(_04606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10645_ (.A1(_00082_),
    .A2(_07797_),
    .B1(\design_top.IADDR[13] ),
    .B2(_07795_),
    .C1(_07796_),
    .X(_04605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10646_ (.A(_07784_),
    .X(_07798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10647_ (.A1(_00081_),
    .A2(_07797_),
    .B1(\design_top.IADDR[12] ),
    .B2(_07798_),
    .C1(_07796_),
    .X(_04604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10648_ (.A(_07789_),
    .X(_07799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10649_ (.A1(_00080_),
    .A2(_07797_),
    .B1(\design_top.IADDR[11] ),
    .B2(_07798_),
    .C1(_07799_),
    .X(_04603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10650_ (.A(_07675_),
    .X(_07800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10651_ (.A1(_00079_),
    .A2(_07800_),
    .B1(\design_top.IADDR[10] ),
    .B2(_07798_),
    .C1(_07799_),
    .X(_04602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10652_ (.A1(_00108_),
    .A2(_07800_),
    .B1(\design_top.IADDR[9] ),
    .B2(_07798_),
    .C1(_07799_),
    .X(_04601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10653_ (.A1(_00107_),
    .A2(_07800_),
    .B1(\design_top.IADDR[8] ),
    .B2(_07798_),
    .C1(_07799_),
    .X(_04600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10654_ (.A(_07655_),
    .X(_07801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10655_ (.A1(_00106_),
    .A2(_07800_),
    .B1(\design_top.IADDR[7] ),
    .B2(_07801_),
    .C1(_07799_),
    .X(_04599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10656_ (.A(_07789_),
    .X(_07802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10657_ (.A1(_00105_),
    .A2(_07800_),
    .B1(\design_top.IADDR[6] ),
    .B2(_07801_),
    .C1(_07802_),
    .X(_04598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10658_ (.A1(_00104_),
    .A2(_07772_),
    .B1(\design_top.IADDR[5] ),
    .B2(_07801_),
    .C1(_07802_),
    .X(_04597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10659_ (.A(\design_top.IADDR[4] ),
    .X(_07803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10660_ (.A1(_00103_),
    .A2(_07772_),
    .B1(_07803_),
    .B2(_07801_),
    .C1(_07802_),
    .X(_04596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10661_ (.A1(_00102_),
    .A2(_07772_),
    .B1(io_out[19]),
    .B2(_07801_),
    .C1(_07802_),
    .X(_04595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10662_ (.A1(_00099_),
    .A2(_07772_),
    .B1(io_out[18]),
    .B2(_07766_),
    .C1(_07802_),
    .X(_04594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10663_ (.A(_07756_),
    .X(_07804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _10664_ (.A1(_00011_),
    .A2(_07804_),
    .B1(_07769_),
    .X(_04593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _10665_ (.A(_07758_),
    .B(\design_top.core0.FLUSH[1] ),
    .C(_06659_),
    .X(_04592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10666_ (.A(_06943_),
    .B(_07629_),
    .X(_07805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10667_ (.A(_07805_),
    .X(_07806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10668_ (.A1(_06901_),
    .A2(_07183_),
    .B1(_07805_),
    .X(_07807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10669_ (.A(_07807_),
    .X(_07808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10670_ (.A1_N(_06940_),
    .A2_N(_07806_),
    .B1(\design_top.MEM[12][23] ),
    .B2(_07808_),
    .X(_04591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10671_ (.A1_N(_06950_),
    .A2_N(_07806_),
    .B1(\design_top.MEM[12][22] ),
    .B2(_07808_),
    .X(_04590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10672_ (.A1_N(_06953_),
    .A2_N(_07806_),
    .B1(\design_top.MEM[12][21] ),
    .B2(_07808_),
    .X(_04589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10673_ (.A1_N(_06956_),
    .A2_N(_07806_),
    .B1(\design_top.MEM[12][20] ),
    .B2(_07808_),
    .X(_04588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10674_ (.A1_N(_06959_),
    .A2_N(_07806_),
    .B1(\design_top.MEM[12][19] ),
    .B2(_07808_),
    .X(_04587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10675_ (.A1_N(_06962_),
    .A2_N(_07805_),
    .B1(\design_top.MEM[12][18] ),
    .B2(_07807_),
    .X(_04586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10676_ (.A1_N(_06965_),
    .A2_N(_07805_),
    .B1(\design_top.MEM[12][17] ),
    .B2(_07807_),
    .X(_04585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _10677_ (.A1_N(_06968_),
    .A2_N(_07805_),
    .B1(\design_top.MEM[12][16] ),
    .B2(_07807_),
    .X(_04584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10678_ (.A(\design_top.core0.FCT3[2] ),
    .Y(_07809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10679_ (.A(\design_top.core0.FCT3[1] ),
    .B(\design_top.core0.FCT3[0] ),
    .X(_07810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10680_ (.A(_07810_),
    .X(_01366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10681_ (.A1(_06787_),
    .A2(_00799_),
    .B1(_06786_),
    .B2(_00796_),
    .X(_07811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10682_ (.A(_01254_),
    .B(_07811_),
    .Y(_01605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10683_ (.A1(_01254_),
    .A2(_07811_),
    .B1(_01605_),
    .Y(_07812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10684_ (.A(_07812_),
    .X(_07813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10685_ (.A(_06764_),
    .B(_01190_),
    .Y(_01192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10686_ (.A1(_06764_),
    .A2(_01190_),
    .B1(_01192_),
    .Y(_07814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10687_ (.A(_07814_),
    .Y(_07815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10688_ (.A(_06768_),
    .B(_01216_),
    .Y(_01217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10689_ (.A1(_06768_),
    .A2(_01216_),
    .B1(_01217_),
    .Y(_07816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10690_ (.A(_07816_),
    .X(_07817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10691_ (.A(_01230_),
    .B(_06769_),
    .Y(_01780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10692_ (.A1(_01230_),
    .A2(_06769_),
    .B1(_01780_),
    .Y(_07818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10693_ (.A(_07818_),
    .Y(_07819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10694_ (.A(_06761_),
    .B(_01204_),
    .Y(_01868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10695_ (.A1(_06761_),
    .A2(_01204_),
    .B1(_01868_),
    .Y(_07820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10696_ (.A(_07820_),
    .Y(_07821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _10697_ (.A(_07815_),
    .B(_07817_),
    .C(_07819_),
    .D(_07821_),
    .X(_07822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10698_ (.A1(_06787_),
    .A2(_00817_),
    .B1(_06786_),
    .B2(_00814_),
    .X(_07823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10699_ (.A(_01238_),
    .B(_07823_),
    .Y(_01239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10700_ (.A1(_01238_),
    .A2(_07823_),
    .B1(_01239_),
    .Y(_07824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10701_ (.A(_07822_),
    .B(_07824_),
    .X(_07825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10702_ (.A(_06788_),
    .X(_07826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10703_ (.A(_01246_),
    .B(_07826_),
    .Y(_01247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10704_ (.A1(_01246_),
    .A2(_07826_),
    .B1(_01247_),
    .Y(_07827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10705_ (.A(_07827_),
    .X(_07828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10706_ (.A(_06726_),
    .B(_01122_),
    .Y(_02051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10707_ (.A1(_06726_),
    .A2(_01122_),
    .B1(_02051_),
    .Y(_07829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10708_ (.A(_07829_),
    .Y(_07830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10709_ (.A(_06805_),
    .B(_01108_),
    .Y(_01109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10710_ (.A1(_06805_),
    .A2(_01108_),
    .B1(_01109_),
    .Y(_07831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10711_ (.A(_06809_),
    .B(_01081_),
    .X(_07832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10712_ (.A(_06809_),
    .B(_01081_),
    .Y(_01083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10713_ (.A(_07832_),
    .B(_01083_),
    .Y(_01305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10714_ (.A(_01305_),
    .Y(_07833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10715_ (.A(_01088_),
    .B(_01095_),
    .Y(_02100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10716_ (.A1(_01088_),
    .A2(_01095_),
    .B1(_02100_),
    .Y(_07834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10717_ (.A(_07834_),
    .Y(_07835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _10718_ (.A(_07830_),
    .B(_07831_),
    .C(_07833_),
    .D(_07835_),
    .X(_07836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10719_ (.A(_01162_),
    .X(_07837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10720_ (.A1(_06786_),
    .A2(_01152_),
    .B1(_06787_),
    .B2(_01155_),
    .X(_07838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10721_ (.A(_01162_),
    .B(_07838_),
    .Y(_01163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10722_ (.A1(_07837_),
    .A2(_07838_),
    .B1(_01163_),
    .Y(_07839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10723_ (.A(_01141_),
    .X(_07840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10724_ (.A(_07840_),
    .B(_01148_),
    .Y(_02004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10725_ (.A1(_07840_),
    .A2(_01148_),
    .B1(_02004_),
    .Y(_07841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10726_ (.A(_07841_),
    .Y(_07842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10727_ (.A(_06754_),
    .B(_01134_),
    .Y(_01135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10728_ (.A1(_06754_),
    .A2(_01134_),
    .B1(_01135_),
    .Y(_07843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10729_ (.A(_06751_),
    .B(_01177_),
    .Y(_01956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10730_ (.A1(_06751_),
    .A2(_01177_),
    .B1(_01956_),
    .Y(_07844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10731_ (.A(_07844_),
    .Y(_07845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _10732_ (.A(_07842_),
    .B(_07843_),
    .C(_07845_),
    .X(_07846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _10733_ (.A(_07828_),
    .B(_07836_),
    .C(_07839_),
    .D(_07846_),
    .X(_07847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10734_ (.A(_01019_),
    .B(_01026_),
    .Y(_01027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10735_ (.A(_01019_),
    .B(_01026_),
    .Y(_02190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10736_ (.A(_02190_),
    .Y(_07848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10737_ (.A(_01027_),
    .B(_07848_),
    .X(_07849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10738_ (.A(_07849_),
    .Y(_07850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10739_ (.A(_01005_),
    .X(_07851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10740_ (.A(_07851_),
    .B(_01012_),
    .X(_07852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10741_ (.A(_07851_),
    .B(_01012_),
    .Y(_01014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10742_ (.A(_07852_),
    .B(_01014_),
    .Y(_01309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10743_ (.A(_01309_),
    .Y(_07853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10744_ (.A(_01068_),
    .B(_06718_),
    .Y(_02146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10745_ (.A1(_01068_),
    .A2(_06718_),
    .B1(_02146_),
    .Y(_01306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10746_ (.A(_01306_),
    .Y(_07854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10747_ (.A(_06716_),
    .B(_01054_),
    .Y(_01055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10748_ (.A1(_06716_),
    .A2(_01054_),
    .B1(_01055_),
    .Y(_07855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _10749_ (.A(_07850_),
    .B(_07853_),
    .C(_07854_),
    .D(_07855_),
    .X(_07856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10750_ (.A(_00897_),
    .X(_07857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10751_ (.A(_07857_),
    .B(_00904_),
    .Y(_00905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10752_ (.A1(_07857_),
    .A2(_00904_),
    .B1(_00905_),
    .Y(_07858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10753_ (.A(_00911_),
    .B(_00918_),
    .Y(_02362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10754_ (.A1(_00911_),
    .A2(_00918_),
    .B1(_02362_),
    .Y(_07859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10755_ (.A(_07859_),
    .Y(_07860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10756_ (.A(_06684_),
    .B(_00931_),
    .Y(_00932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10757_ (.A1(_06684_),
    .A2(_00931_),
    .B1(_00932_),
    .Y(_07861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10758_ (.A(_00945_),
    .B(_06686_),
    .Y(_02319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10759_ (.A1(_00945_),
    .A2(_06686_),
    .B1(_02319_),
    .Y(_07862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4b_2 _10760_ (.A(_07858_),
    .B(_07860_),
    .C(_07861_),
    .D_N(_07862_),
    .X(_07863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10761_ (.A(_06841_),
    .B(_00849_),
    .Y(_00850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10762_ (.A1(_06841_),
    .A2(_00849_),
    .B1(_00850_),
    .Y(_07864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10763_ (.A(_00870_),
    .B(_00877_),
    .Y(_00879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10764_ (.A1(_00870_),
    .A2(_00877_),
    .B1(_00879_),
    .Y(_01319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10765_ (.A(_01319_),
    .Y(_07865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10766_ (.A(_00884_),
    .B(_00891_),
    .Y(_00892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10767_ (.A1(_00884_),
    .A2(_00891_),
    .B1(_00892_),
    .Y(_07866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10768_ (.A(_00856_),
    .B(_00863_),
    .Y(_00865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10769_ (.A1(_00856_),
    .A2(_00863_),
    .B1(_00865_),
    .Y(_01320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10770_ (.A(_01320_),
    .Y(_07867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _10771_ (.A(_07864_),
    .B(_07865_),
    .C(_07866_),
    .D(_07867_),
    .X(_07868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10772_ (.A(_06702_),
    .B(_00958_),
    .X(_07869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10773_ (.A(_06702_),
    .B(_00958_),
    .Y(_00960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10774_ (.A(_07869_),
    .B(_00960_),
    .Y(_01313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10775_ (.A(_01313_),
    .Y(_07870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10776_ (.A(_06821_),
    .B(_00985_),
    .Y(_00986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10777_ (.A1(_06821_),
    .A2(_00985_),
    .B1(_00986_),
    .Y(_07871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10778_ (.A(_06691_),
    .B(_00999_),
    .Y(_02233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10779_ (.A1(_06691_),
    .A2(_00999_),
    .B1(_02233_),
    .Y(_07872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10780_ (.A(_07872_),
    .Y(_07873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10781_ (.A(_00965_),
    .B(_00972_),
    .Y(_02276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10782_ (.A1(_00965_),
    .A2(_00972_),
    .B1(_02276_),
    .Y(_07874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10783_ (.A(_07874_),
    .Y(_07875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _10784_ (.A(_07870_),
    .B(_07871_),
    .C(_07873_),
    .D(_07875_),
    .X(_07876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _10785_ (.A(_07856_),
    .B(_07863_),
    .C(_07868_),
    .D(_07876_),
    .X(_07877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _10786_ (.A(_07813_),
    .B(_07825_),
    .C(_07847_),
    .D(_07877_),
    .X(_07878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10787_ (.A(_01328_),
    .Y(_07879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _10788_ (.A1(_07809_),
    .A2(_01366_),
    .A3(_07878_),
    .B1(_07879_),
    .X(_07880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10789_ (.A1(\design_top.core0.XJALR ),
    .A2(\design_top.core0.XJAL ),
    .B1(_00786_),
    .X(_00822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _10790_ (.A1(\design_top.core0.XBCC ),
    .A2(_00786_),
    .A3(_07880_),
    .B1(_00822_),
    .X(_01518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10791_ (.A(_01518_),
    .Y(_01329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10792_ (.A(_07658_),
    .B(_01329_),
    .X(_07881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10793_ (.A(_07881_),
    .Y(_07882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10794_ (.A(_02469_),
    .Y(_07883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10795_ (.A1(io_out[17]),
    .A2(_07882_),
    .B1(_07883_),
    .B2(_07881_),
    .C1(_07758_),
    .X(_04583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10796_ (.A(_02468_),
    .Y(_07884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10797_ (.A1(io_out[16]),
    .A2(_07882_),
    .B1(_07884_),
    .B2(_07881_),
    .C1(_07758_),
    .X(_04582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10798_ (.A(\design_top.uart0.UART_RBAUD[1] ),
    .B(\design_top.uart0.UART_RBAUD[0] ),
    .X(_07885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _10799_ (.A(\design_top.uart0.UART_RBAUD[2] ),
    .B(_07885_),
    .C(\design_top.uart0.UART_RBAUD[3] ),
    .X(_07886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10800_ (.A(\design_top.uart0.UART_RBAUD[4] ),
    .B(_07886_),
    .X(_07887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10801_ (.A(\design_top.uart0.UART_RBAUD[5] ),
    .B(_07887_),
    .X(_07888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10802_ (.A(\design_top.uart0.UART_RBAUD[6] ),
    .B(_07888_),
    .X(_07889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10803_ (.A(\design_top.uart0.UART_RBAUD[7] ),
    .B(_07889_),
    .X(_07890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10804_ (.A(\design_top.uart0.UART_RBAUD[8] ),
    .B(_07890_),
    .X(_07891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10805_ (.A(\design_top.uart0.UART_RBAUD[9] ),
    .B(_07891_),
    .X(_07892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10806_ (.A(\design_top.uart0.UART_RBAUD[10] ),
    .B(_07892_),
    .X(_07893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10807_ (.A(\design_top.uart0.UART_RBAUD[11] ),
    .B(_07893_),
    .X(_07894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10808_ (.A(\design_top.uart0.UART_RBAUD[12] ),
    .B(_07894_),
    .X(_07895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10809_ (.A(\design_top.uart0.UART_RBAUD[13] ),
    .B(_07895_),
    .X(_07896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _10810_ (.A(\design_top.uart0.UART_RBAUD[14] ),
    .B(_07896_),
    .C(\design_top.uart0.UART_RBAUD[15] ),
    .X(_02591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10811_ (.A(_02591_),
    .Y(_07897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10812_ (.A(\design_top.uart0.UART_RSTATE[1] ),
    .Y(_07898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10813_ (.A(\design_top.uart0.UART_RSTATE[2] ),
    .Y(_07899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _10814_ (.A(_07898_),
    .B(\design_top.uart0.UART_RSTATE[0] ),
    .C(\design_top.uart0.UART_RSTATE[3] ),
    .D(_07899_),
    .X(_07900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10815_ (.A(_07900_),
    .Y(_01370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10816_ (.A(_07897_),
    .B(_01370_),
    .X(_07901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10817_ (.A(_07901_),
    .Y(_07902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _10818_ (.A1(\design_top.uart0.UART_RBAUD[14] ),
    .A2(_07896_),
    .B1(\design_top.uart0.UART_RBAUD[15] ),
    .C1(_07902_),
    .X(_04581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10819_ (.A(_07901_),
    .X(_07903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _10820_ (.A1_N(\design_top.uart0.UART_RBAUD[14] ),
    .A2_N(_07896_),
    .B1(\design_top.uart0.UART_RBAUD[14] ),
    .B2(_07896_),
    .Y(_07904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10821_ (.A(_07903_),
    .B(_07904_),
    .Y(_04580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10822_ (.A(\design_top.uart0.UART_RBAUD[13] ),
    .B(_07895_),
    .Y(_07905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10823_ (.A1(_07896_),
    .A2(_07905_),
    .B1(_07903_),
    .Y(_04579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10824_ (.A(\design_top.uart0.UART_RBAUD[12] ),
    .B(_07894_),
    .Y(_07906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10825_ (.A1(_07895_),
    .A2(_07906_),
    .B1(_07903_),
    .Y(_04578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10826_ (.A(\design_top.uart0.UART_RBAUD[11] ),
    .B(_07893_),
    .Y(_07907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10827_ (.A1(_07894_),
    .A2(_07907_),
    .B1(_07903_),
    .Y(_04577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10828_ (.A(\design_top.uart0.UART_RBAUD[10] ),
    .B(_07892_),
    .Y(_07908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10829_ (.A1(_07893_),
    .A2(_07908_),
    .B1(_07901_),
    .Y(_04576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10830_ (.A(_07891_),
    .Y(_07909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _10831_ (.A1(\design_top.uart0.UART_RBAUD[8] ),
    .A2(_07890_),
    .B1(_07909_),
    .C1(_07901_),
    .X(_04575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10832_ (.A(_07888_),
    .Y(_07910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _10833_ (.A1(\design_top.uart0.UART_RBAUD[5] ),
    .A2(_07887_),
    .B1(_07910_),
    .C1(_07901_),
    .X(_04574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10834_ (.A(_07886_),
    .Y(_07911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10835_ (.A1(\design_top.uart0.UART_RBAUD[2] ),
    .A2(_07885_),
    .B1(\design_top.uart0.UART_RBAUD[3] ),
    .X(_07912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10836_ (.A1(_07911_),
    .A2(_07912_),
    .B1(_07902_),
    .X(_04573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10837_ (.A(\design_top.uart0.UART_RBAUD[0] ),
    .B(_07903_),
    .Y(_04572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _10838_ (.A(\design_top.uart0.UART_XBAUD[1] ),
    .B(\design_top.uart0.UART_XBAUD[0] ),
    .C(\design_top.uart0.UART_XBAUD[2] ),
    .D(\design_top.uart0.UART_XBAUD[3] ),
    .X(_07913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10839_ (.A(\design_top.uart0.UART_XBAUD[4] ),
    .B(_07913_),
    .X(_07914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10840_ (.A(\design_top.uart0.UART_XBAUD[5] ),
    .B(_07914_),
    .X(_07915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10841_ (.A(\design_top.uart0.UART_XBAUD[6] ),
    .B(_07915_),
    .X(_07916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10842_ (.A(\design_top.uart0.UART_XBAUD[7] ),
    .B(_07916_),
    .X(_07917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10843_ (.A(\design_top.uart0.UART_XBAUD[8] ),
    .B(_07917_),
    .X(_07918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10844_ (.A(\design_top.uart0.UART_XBAUD[9] ),
    .B(_07918_),
    .X(_07919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10845_ (.A(\design_top.uart0.UART_XBAUD[10] ),
    .B(_07919_),
    .X(_07920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10846_ (.A(\design_top.uart0.UART_XBAUD[11] ),
    .B(_07920_),
    .X(_07921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10847_ (.A(\design_top.uart0.UART_XBAUD[12] ),
    .B(_07921_),
    .X(_07922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10848_ (.A(\design_top.uart0.UART_XBAUD[13] ),
    .B(_07922_),
    .X(_07923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10849_ (.A(\design_top.uart0.UART_XSTATE[1] ),
    .Y(_07924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10850_ (.A(\design_top.uart0.UART_XSTATE[2] ),
    .Y(_07925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _10851_ (.A(_07924_),
    .B(\design_top.uart0.UART_XSTATE[3] ),
    .C(_07925_),
    .X(_07926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _10852_ (.A(\design_top.uart0.UART_XBAUD[14] ),
    .B(_07923_),
    .C(\design_top.uart0.UART_XBAUD[15] ),
    .X(_07927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10853_ (.A(_07927_),
    .X(_00782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10854_ (.A1(\design_top.uart0.UART_XSTATE[0] ),
    .A2(_07926_),
    .B1(_00782_),
    .Y(_07928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10855_ (.A(_07928_),
    .Y(_07929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _10856_ (.A1(\design_top.uart0.UART_XBAUD[14] ),
    .A2(_07923_),
    .B1(\design_top.uart0.UART_XBAUD[15] ),
    .C1(_07929_),
    .X(_04571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10857_ (.A(_07928_),
    .X(_07930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10858_ (.A(_07930_),
    .X(_07931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _10859_ (.A1_N(\design_top.uart0.UART_XBAUD[14] ),
    .A2_N(_07923_),
    .B1(\design_top.uart0.UART_XBAUD[14] ),
    .B2(_07923_),
    .Y(_07932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10860_ (.A(_07931_),
    .B(_07932_),
    .Y(_04570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10861_ (.A(\design_top.uart0.UART_XBAUD[13] ),
    .B(_07922_),
    .Y(_07933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10862_ (.A1(_07923_),
    .A2(_07933_),
    .B1(_07931_),
    .Y(_04569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10863_ (.A(\design_top.uart0.UART_XBAUD[12] ),
    .B(_07921_),
    .Y(_07934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10864_ (.A1(_07922_),
    .A2(_07934_),
    .B1(_07931_),
    .Y(_04568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10865_ (.A(\design_top.uart0.UART_XBAUD[11] ),
    .B(_07920_),
    .Y(_07935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10866_ (.A(_07930_),
    .X(_07936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10867_ (.A1(_07921_),
    .A2(_07935_),
    .B1(_07936_),
    .Y(_04567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10868_ (.A(\design_top.uart0.UART_XBAUD[10] ),
    .B(_07919_),
    .Y(_07937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10869_ (.A1(_07920_),
    .A2(_07937_),
    .B1(_07936_),
    .Y(_04566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10870_ (.A(_07919_),
    .Y(_07938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _10871_ (.A1(\design_top.uart0.UART_XBAUD[9] ),
    .A2(_07918_),
    .B1(_07938_),
    .C1(_07936_),
    .X(_04565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10872_ (.A(_07918_),
    .Y(_07939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _10873_ (.A1(\design_top.uart0.UART_XBAUD[8] ),
    .A2(_07917_),
    .B1(_07939_),
    .C1(_07930_),
    .X(_04564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10874_ (.A(\design_top.uart0.UART_XBAUD[7] ),
    .B(_07916_),
    .Y(_07940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10875_ (.A1(_07917_),
    .A2(_07940_),
    .B1(_07936_),
    .Y(_04563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10876_ (.A(_07916_),
    .Y(_07941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _10877_ (.A1(\design_top.uart0.UART_XBAUD[6] ),
    .A2(_07915_),
    .B1(_07941_),
    .C1(_07930_),
    .X(_04562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10878_ (.A(_07915_),
    .Y(_07942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _10879_ (.A1(\design_top.uart0.UART_XBAUD[5] ),
    .A2(_07914_),
    .B1(_07942_),
    .C1(_07930_),
    .X(_04561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10880_ (.A(\design_top.uart0.UART_XBAUD[4] ),
    .B(_07913_),
    .Y(_07943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10881_ (.A1(_07914_),
    .A2(_07943_),
    .B1(_07936_),
    .Y(_04560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10882_ (.A(_07913_),
    .Y(_07944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10883_ (.A(\design_top.uart0.UART_XBAUD[1] ),
    .X(_07945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10884_ (.A(\design_top.uart0.UART_XBAUD[0] ),
    .X(_07946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _10885_ (.A1(_07945_),
    .A2(_07946_),
    .A3(\design_top.uart0.UART_XBAUD[2] ),
    .B1(\design_top.uart0.UART_XBAUD[3] ),
    .X(_07947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10886_ (.A1(_07944_),
    .A2(_07947_),
    .B1(_07929_),
    .X(_04559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10887_ (.A1(_07945_),
    .A2(\design_top.uart0.UART_XBAUD[0] ),
    .B1(\design_top.uart0.UART_XBAUD[2] ),
    .Y(_07948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o311a_2 _10888_ (.A1(_07945_),
    .A2(_07946_),
    .A3(\design_top.uart0.UART_XBAUD[2] ),
    .B1(_07948_),
    .C1(_07929_),
    .X(_07949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10889_ (.A(_07949_),
    .Y(_04558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _10890_ (.A1_N(_07945_),
    .A2_N(_07946_),
    .B1(_07945_),
    .B2(_07946_),
    .Y(_07950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10891_ (.A(_07931_),
    .B(_07950_),
    .Y(_04557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10892_ (.A(_07946_),
    .B(_07931_),
    .Y(_04556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10893_ (.A(_07760_),
    .B(_00007_),
    .X(_04555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10894_ (.A(_07760_),
    .B(_00006_),
    .X(_04554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10895_ (.A(_07760_),
    .B(_00005_),
    .X(_04553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10896_ (.A(_07760_),
    .B(_00004_),
    .X(_04552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _10897_ (.A(_07622_),
    .B(\design_top.DACK[1] ),
    .C(\design_top.DACK[0] ),
    .X(_04551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10898_ (.A(_06992_),
    .B(_00012_),
    .X(_04550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10899_ (.A(\design_top.uart0.UART_XSTATE[3] ),
    .Y(_07951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a41o_2 _10900_ (.A1(_07924_),
    .A2(\design_top.uart0.UART_XSTATE[0] ),
    .A3(_07951_),
    .A4(_07925_),
    .B1(_07623_),
    .X(_07952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10901_ (.A(\design_top.uart0.UART_XSTATE[0] ),
    .Y(_07953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _10902_ (.A(_07953_),
    .B(_00783_),
    .C(_07924_),
    .X(_07954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10903_ (.A(_07925_),
    .B(_07954_),
    .Y(_07955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _10904_ (.A1(_07953_),
    .A2(_00783_),
    .A3(_07926_),
    .B1(_07951_),
    .B2(_07955_),
    .X(_07956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10905_ (.A(_07952_),
    .B(_07956_),
    .Y(_04549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10906_ (.A1(_07925_),
    .A2(_07954_),
    .B1(_07955_),
    .Y(_07957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10907_ (.A(_07952_),
    .B(_07957_),
    .X(_04548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10908_ (.A(_07954_),
    .Y(_07958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10909_ (.A1(_07953_),
    .A2(_00783_),
    .B1(_07924_),
    .X(_07959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10910_ (.A(_07952_),
    .Y(_07960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10911_ (.A1(_07958_),
    .A2(_07959_),
    .B1(_07960_),
    .Y(_04547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10912_ (.A(_00783_),
    .Y(_07961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10913_ (.A1(_07953_),
    .A2(_00783_),
    .B1(\design_top.uart0.UART_XSTATE[0] ),
    .B2(_07961_),
    .C1(_07960_),
    .X(_04546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10914_ (.A(_07899_),
    .X(_07962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10915_ (.A(\design_top.uart0.UART_RSTATE[0] ),
    .Y(_07963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _10916_ (.A(_07963_),
    .B(_00785_),
    .C(_07898_),
    .X(_07964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10917_ (.A(\design_top.uart0.UART_RSTATE[3] ),
    .Y(_07965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10918_ (.A(_07965_),
    .X(_07966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10919_ (.A(\design_top.uart0.UART_RSTATE[1] ),
    .X(_07967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _10920_ (.A(_07967_),
    .B(_07963_),
    .C(\design_top.uart0.UART_RSTATE[3] ),
    .D(\design_top.uart0.UART_RSTATE[2] ),
    .X(_07968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10921_ (.A(_06991_),
    .B(_07968_),
    .Y(_07969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10922_ (.A(_07969_),
    .Y(_07970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10923_ (.A1(_07962_),
    .A2(_07964_),
    .B1(_07966_),
    .Y(_07971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o311a_2 _10924_ (.A1(_07962_),
    .A2(_07964_),
    .A3(_07966_),
    .B1(_07970_),
    .C1(_07971_),
    .X(_04545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10925_ (.A(\design_top.uart0.UART_RSTATE[2] ),
    .X(_07972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10926_ (.A(_07964_),
    .Y(_07973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _10927_ (.A1(_07962_),
    .A2(_07964_),
    .B1(_07972_),
    .B2(_07973_),
    .X(_07974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10928_ (.A(_07969_),
    .B(_07974_),
    .X(_04544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10929_ (.A(_07963_),
    .X(_07975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10930_ (.A(_07898_),
    .X(_07976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10931_ (.A1(_07975_),
    .A2(_00785_),
    .B1(_07976_),
    .X(_07977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10932_ (.A1(_07973_),
    .A2(_07977_),
    .B1(_07970_),
    .Y(_04543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10933_ (.A(\design_top.uart0.UART_RSTATE[0] ),
    .X(_07978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10934_ (.A(_00785_),
    .Y(_07979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _10935_ (.A1(_07975_),
    .A2(_00785_),
    .B1(_07978_),
    .B2(_07979_),
    .C1(_07970_),
    .X(_04542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10936_ (.A(_07892_),
    .Y(_07980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10937_ (.A(\design_top.uart0.UART_RBAUD[9] ),
    .B(_07891_),
    .X(_07981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10938_ (.A(_07900_),
    .X(_07982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10939_ (.A1(_07980_),
    .A2(_07981_),
    .B1(_07982_),
    .X(_04541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _10940_ (.A1(\design_top.uart0.UART_RBAUD[7] ),
    .A2(_07889_),
    .B1_N(_07890_),
    .Y(_07983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10941_ (.A1(_07897_),
    .A2(_07983_),
    .B1(_07982_),
    .Y(_04540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10942_ (.A(_07889_),
    .Y(_07984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10943_ (.A(\design_top.uart0.UART_RBAUD[6] ),
    .B(_07888_),
    .X(_07985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10944_ (.A1(_07984_),
    .A2(_07985_),
    .B1(_07982_),
    .X(_04539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _10945_ (.A1(\design_top.uart0.UART_RBAUD[4] ),
    .A2(_07886_),
    .B1_N(_07887_),
    .Y(_07986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10946_ (.A1(_07897_),
    .A2(_07986_),
    .B1(_07982_),
    .Y(_04538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _10947_ (.A1_N(\design_top.uart0.UART_RBAUD[2] ),
    .A2_N(_07885_),
    .B1(\design_top.uart0.UART_RBAUD[2] ),
    .B2(_07885_),
    .Y(_07987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10948_ (.A(_01370_),
    .B(_07987_),
    .Y(_04537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _10949_ (.A1(\design_top.uart0.UART_RBAUD[1] ),
    .A2(\design_top.uart0.UART_RBAUD[0] ),
    .B1_N(_07885_),
    .Y(_07988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10950_ (.A1(_07897_),
    .A2(_07988_),
    .B1(_07982_),
    .Y(_04536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10951_ (.A(_07723_),
    .B(_00003_),
    .X(_04535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10952_ (.A(_07723_),
    .B(_00002_),
    .X(_04534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10953_ (.A(_07723_),
    .B(_00001_),
    .X(_04533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _10954_ (.A(_07723_),
    .B(_00000_),
    .X(_04532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10955_ (.A(\design_top.core0.RESMODE[2] ),
    .Y(_07989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10956_ (.A(\design_top.core0.RESMODE[0] ),
    .B(\design_top.core0.RESMODE[1] ),
    .Y(_01330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _10957_ (.A(_07989_),
    .B(_01330_),
    .Y(_07990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _10958_ (.A1(\design_top.core0.RESMODE[3] ),
    .A2(_07990_),
    .B1(_07624_),
    .X(_04531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10959_ (.A1(_07989_),
    .A2(_01330_),
    .B1(_07031_),
    .Y(_07991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _10960_ (.A1(_07989_),
    .A2(_01330_),
    .A3(\design_top.core0.RESMODE[3] ),
    .B1(_07991_),
    .X(_04530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10961_ (.A(_07624_),
    .B(_00078_),
    .X(_04529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10962_ (.A(\design_top.core0.RESMODE[0] ),
    .Y(_07992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10963_ (.A(\design_top.core0.RESMODE[2] ),
    .B(\design_top.core0.RESMODE[3] ),
    .X(_07993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10964_ (.A(_07993_),
    .X(_01331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _10965_ (.A(\design_top.core0.RESMODE[0] ),
    .B(\design_top.core0.RESMODE[1] ),
    .C(_01331_),
    .X(_00046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _10966_ (.A1(_07992_),
    .A2(_00046_),
    .B1(_07624_),
    .X(_04528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10967_ (.A(_07031_),
    .X(_07994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10968_ (.A(\design_top.IRES[0] ),
    .B(\design_top.IRES[1] ),
    .X(_07995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _10969_ (.A(\design_top.IRES[2] ),
    .B(_07995_),
    .C(\design_top.IRES[3] ),
    .X(_07996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10970_ (.A(\design_top.IRES[4] ),
    .B(_07996_),
    .X(_07997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10971_ (.A(\design_top.IRES[5] ),
    .B(_07997_),
    .X(_07998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _10972_ (.A(\design_top.IRES[6] ),
    .B(_07998_),
    .Y(_07999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10973_ (.A(_06862_),
    .X(_08000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10974_ (.A1(_07994_),
    .A2(_07999_),
    .B1(_08000_),
    .Y(_04527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _10975_ (.A1(\design_top.IRES[6] ),
    .A2(_07998_),
    .B1(_07999_),
    .Y(_08001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10976_ (.A1(_07994_),
    .A2(_08001_),
    .B1(_08000_),
    .Y(_04526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _10977_ (.A1(\design_top.IRES[5] ),
    .A2(_07997_),
    .B1_N(_07998_),
    .Y(_08002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10978_ (.A1(_07994_),
    .A2(_08002_),
    .B1(_08000_),
    .Y(_04525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _10979_ (.A1(\design_top.IRES[4] ),
    .A2(_07996_),
    .B1_N(_07997_),
    .Y(_08003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10980_ (.A1(_07994_),
    .A2(_08003_),
    .B1(_08000_),
    .Y(_04524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _10981_ (.A1(\design_top.IRES[2] ),
    .A2(_07995_),
    .B1(\design_top.IRES[3] ),
    .X(_08004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2b_2 _10982_ (.A_N(_08004_),
    .B(_07996_),
    .X(_08005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10983_ (.A1(_07994_),
    .A2(_08005_),
    .B1(_08000_),
    .Y(_04523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _10984_ (.A1_N(\design_top.IRES[2] ),
    .A2_N(_07995_),
    .B1(\design_top.IRES[2] ),
    .B2(_07995_),
    .Y(_08006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10985_ (.A1(_06992_),
    .A2(_08006_),
    .B1(_06862_),
    .Y(_04522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _10986_ (.A1(\design_top.IRES[0] ),
    .A2(\design_top.IRES[1] ),
    .B1_N(_07995_),
    .Y(_08007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10987_ (.A1(_06992_),
    .A2(_08007_),
    .B1(_06862_),
    .Y(_04521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _10988_ (.A1(_06992_),
    .A2(\design_top.IRES[0] ),
    .B1(_06862_),
    .Y(_04520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _10989_ (.A(\design_top.DACK[1] ),
    .B(_02944_),
    .C(_01380_),
    .Y(_08008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _10990_ (.A(_06986_),
    .B(_07154_),
    .X(_08009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10991_ (.A(_08009_),
    .Y(_08010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _10992_ (.A1(io_out[12]),
    .A2(_08008_),
    .A3(_08010_),
    .B1(_07623_),
    .X(_08011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _10993_ (.A0(\design_top.uart0.UART_RACK ),
    .A1(\design_top.uart0.UART_RREQ ),
    .S(_08011_),
    .X(_04519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _10994_ (.A(\design_top.uart0.UART_XACK ),
    .Y(_08012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _10995_ (.A(_07658_),
    .B(_06664_),
    .C(_01380_),
    .D(_08009_),
    .X(_08013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _10996_ (.A(_08013_),
    .X(_08014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _10997_ (.A0(_08012_),
    .A1(\design_top.uart0.UART_XREQ ),
    .S(_08014_),
    .X(_04518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _10998_ (.A0(\design_top.DATAO[15] ),
    .A1(\design_top.uart0.UART_XFIFO[7] ),
    .S(_08014_),
    .X(_04517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _10999_ (.A0(\design_top.DATAO[14] ),
    .A1(\design_top.uart0.UART_XFIFO[6] ),
    .S(_08014_),
    .X(_04516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _11000_ (.A0(\design_top.DATAO[13] ),
    .A1(\design_top.uart0.UART_XFIFO[5] ),
    .S(_08014_),
    .X(_04515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _11001_ (.A0(\design_top.DATAO[12] ),
    .A1(\design_top.uart0.UART_XFIFO[4] ),
    .S(_08014_),
    .X(_04514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _11002_ (.A0(\design_top.DATAO[11] ),
    .A1(\design_top.uart0.UART_XFIFO[3] ),
    .S(_08013_),
    .X(_04513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _11003_ (.A0(\design_top.DATAO[10] ),
    .A1(\design_top.uart0.UART_XFIFO[2] ),
    .S(_08013_),
    .X(_04512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _11004_ (.A0(\design_top.DATAO[9] ),
    .A1(\design_top.uart0.UART_XFIFO[1] ),
    .S(_08013_),
    .X(_04511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _11005_ (.A0(\design_top.DATAO[8] ),
    .A1(\design_top.uart0.UART_XFIFO[0] ),
    .S(_08013_),
    .X(_04510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11006_ (.A(_01382_),
    .B(_06843_),
    .X(_08015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11007_ (.A(_08015_),
    .X(_08016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11008_ (.A1(_07150_),
    .A2(_06903_),
    .B1(_06897_),
    .B2(_08016_),
    .X(_08017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11009_ (.A(_08017_),
    .Y(_08018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11010_ (.A(_08018_),
    .X(_08019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11011_ (.A(_08017_),
    .X(_08020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11012_ (.A1(_00180_),
    .A2(_08019_),
    .B1(\design_top.MEM[0][7] ),
    .B2(_08020_),
    .X(_04509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11013_ (.A1(_00179_),
    .A2(_08019_),
    .B1(\design_top.MEM[0][6] ),
    .B2(_08020_),
    .X(_04508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11014_ (.A1(_00178_),
    .A2(_08019_),
    .B1(\design_top.MEM[0][5] ),
    .B2(_08020_),
    .X(_04507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11015_ (.A1(_00177_),
    .A2(_08019_),
    .B1(\design_top.MEM[0][4] ),
    .B2(_08020_),
    .X(_04506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11016_ (.A1(_00176_),
    .A2(_08019_),
    .B1(\design_top.MEM[0][3] ),
    .B2(_08020_),
    .X(_04505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11017_ (.A1(_00175_),
    .A2(_08018_),
    .B1(\design_top.MEM[0][2] ),
    .B2(_08017_),
    .X(_04504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11018_ (.A1(_00174_),
    .A2(_08018_),
    .B1(\design_top.MEM[0][1] ),
    .B2(_08017_),
    .X(_04503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11019_ (.A1(_00173_),
    .A2(_08018_),
    .B1(\design_top.MEM[0][0] ),
    .B2(_08017_),
    .X(_04502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11020_ (.A(_06976_),
    .X(_08021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11021_ (.A(_08015_),
    .X(_08022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11022_ (.A(_08022_),
    .X(_08023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11023_ (.A1(_06869_),
    .A2(_08021_),
    .B1(_06972_),
    .B2(_08023_),
    .X(_08024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11024_ (.A(_08024_),
    .Y(_08025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11025_ (.A(_08025_),
    .X(_08026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11026_ (.A(_08024_),
    .X(_08027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11027_ (.A1(_00188_),
    .A2(_08026_),
    .B1(\design_top.MEM[10][7] ),
    .B2(_08027_),
    .X(_04501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11028_ (.A1(_00187_),
    .A2(_08026_),
    .B1(\design_top.MEM[10][6] ),
    .B2(_08027_),
    .X(_04500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11029_ (.A1(_00186_),
    .A2(_08026_),
    .B1(\design_top.MEM[10][5] ),
    .B2(_08027_),
    .X(_04499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11030_ (.A1(_00185_),
    .A2(_08026_),
    .B1(\design_top.MEM[10][4] ),
    .B2(_08027_),
    .X(_04498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11031_ (.A1(_00184_),
    .A2(_08026_),
    .B1(\design_top.MEM[10][3] ),
    .B2(_08027_),
    .X(_04497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11032_ (.A1(_00183_),
    .A2(_08025_),
    .B1(\design_top.MEM[10][2] ),
    .B2(_08024_),
    .X(_04496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11033_ (.A1(_00182_),
    .A2(_08025_),
    .B1(\design_top.MEM[10][1] ),
    .B2(_08024_),
    .X(_04495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11034_ (.A1(_00181_),
    .A2(_08025_),
    .B1(\design_top.MEM[10][0] ),
    .B2(_08024_),
    .X(_04494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11035_ (.A(\design_top.IRES[7] ),
    .B(_07003_),
    .X(_08028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11036_ (.A(_08028_),
    .X(_08029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11037_ (.A(_08029_),
    .X(_08030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11038_ (.A(_08030_),
    .X(_08031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11039_ (.A(_08028_),
    .Y(_08032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11040_ (.A(_08032_),
    .X(_08033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11041_ (.A1(\design_top.TIMER[31] ),
    .A2(_08031_),
    .B1(_00037_),
    .B2(_08033_),
    .X(_04493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11042_ (.A1(\design_top.TIMER[30] ),
    .A2(_08031_),
    .B1(_00036_),
    .B2(_08033_),
    .X(_04492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11043_ (.A1(\design_top.TIMER[29] ),
    .A2(_08031_),
    .B1(_00034_),
    .B2(_08033_),
    .X(_04491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11044_ (.A1(\design_top.TIMER[28] ),
    .A2(_08031_),
    .B1(_00033_),
    .B2(_08033_),
    .X(_04490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11045_ (.A(_08032_),
    .X(_08034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11046_ (.A(_08034_),
    .X(_08035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11047_ (.A1(\design_top.TIMER[27] ),
    .A2(_08031_),
    .B1(_00032_),
    .B2(_08035_),
    .X(_04489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11048_ (.A(_08030_),
    .X(_08036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11049_ (.A1(\design_top.TIMER[26] ),
    .A2(_08036_),
    .B1(_00031_),
    .B2(_08035_),
    .X(_04488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11050_ (.A1(\design_top.TIMER[25] ),
    .A2(_08036_),
    .B1(_00030_),
    .B2(_08035_),
    .X(_04487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11051_ (.A1(\design_top.TIMER[24] ),
    .A2(_08036_),
    .B1(_00029_),
    .B2(_08035_),
    .X(_04486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11052_ (.A1(\design_top.TIMER[23] ),
    .A2(_08036_),
    .B1(_00028_),
    .B2(_08035_),
    .X(_04485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11053_ (.A(_08034_),
    .X(_08037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11054_ (.A1(\design_top.TIMER[22] ),
    .A2(_08036_),
    .B1(_00027_),
    .B2(_08037_),
    .X(_04484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11055_ (.A(_08029_),
    .X(_08038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11056_ (.A1(\design_top.TIMER[21] ),
    .A2(_08038_),
    .B1(_00026_),
    .B2(_08037_),
    .X(_04483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11057_ (.A1(\design_top.TIMER[20] ),
    .A2(_08038_),
    .B1(_00025_),
    .B2(_08037_),
    .X(_04482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11058_ (.A1(\design_top.TIMER[19] ),
    .A2(_08038_),
    .B1(_00023_),
    .B2(_08037_),
    .X(_04481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11059_ (.A1(\design_top.TIMER[18] ),
    .A2(_08038_),
    .B1(_00022_),
    .B2(_08037_),
    .X(_04480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11060_ (.A(_08032_),
    .X(_08039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11061_ (.A1(\design_top.TIMER[17] ),
    .A2(_08038_),
    .B1(_00021_),
    .B2(_08039_),
    .X(_04479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11062_ (.A(_08029_),
    .X(_08040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11063_ (.A1(\design_top.TIMER[16] ),
    .A2(_08040_),
    .B1(_00020_),
    .B2(_08039_),
    .X(_04478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11064_ (.A1(\design_top.TIMER[15] ),
    .A2(_08040_),
    .B1(_00019_),
    .B2(_08039_),
    .X(_04477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11065_ (.A1(\design_top.TIMER[14] ),
    .A2(_08040_),
    .B1(_00018_),
    .B2(_08039_),
    .X(_04476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11066_ (.A1(\design_top.TIMER[13] ),
    .A2(_08040_),
    .B1(_00017_),
    .B2(_08039_),
    .X(_04475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11067_ (.A(_08032_),
    .X(_08041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11068_ (.A1(\design_top.TIMER[12] ),
    .A2(_08040_),
    .B1(_00016_),
    .B2(_08041_),
    .X(_04474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11069_ (.A(_08029_),
    .X(_08042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11070_ (.A1(\design_top.TIMER[11] ),
    .A2(_08042_),
    .B1(_00015_),
    .B2(_08041_),
    .X(_04473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11071_ (.A1(\design_top.TIMER[10] ),
    .A2(_08042_),
    .B1(_00014_),
    .B2(_08041_),
    .X(_04472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11072_ (.A1(\design_top.TIMER[9] ),
    .A2(_08042_),
    .B1(_00044_),
    .B2(_08041_),
    .X(_04471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11073_ (.A1(\design_top.TIMER[8] ),
    .A2(_08042_),
    .B1(_00043_),
    .B2(_08041_),
    .X(_04470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11074_ (.A(_08032_),
    .X(_08043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11075_ (.A1(\design_top.TIMER[7] ),
    .A2(_08042_),
    .B1(_00042_),
    .B2(_08043_),
    .X(_04469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11076_ (.A(_08029_),
    .X(_08044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11077_ (.A1(\design_top.TIMER[6] ),
    .A2(_08044_),
    .B1(_00041_),
    .B2(_08043_),
    .X(_04468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11078_ (.A1(\design_top.TIMER[5] ),
    .A2(_08044_),
    .B1(_00040_),
    .B2(_08043_),
    .X(_04467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11079_ (.A1(\design_top.TIMER[4] ),
    .A2(_08044_),
    .B1(_00039_),
    .B2(_08043_),
    .X(_04466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11080_ (.A1(\design_top.TIMER[3] ),
    .A2(_08044_),
    .B1(_00038_),
    .B2(_08043_),
    .X(_04465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11081_ (.A1(\design_top.TIMER[2] ),
    .A2(_08044_),
    .B1(_00035_),
    .B2(_08034_),
    .X(_04464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11082_ (.A1(\design_top.TIMER[1] ),
    .A2(_08030_),
    .B1(_00024_),
    .B2(_08034_),
    .X(_04463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11083_ (.A1(\design_top.TIMER[0] ),
    .A2(_08030_),
    .B1(_00013_),
    .B2(_08034_),
    .X(_04462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11084_ (.A(_07047_),
    .X(_08045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11085_ (.A1(_06868_),
    .A2(_08045_),
    .B1(_07044_),
    .B2(_08023_),
    .X(_08046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11086_ (.A(_08046_),
    .Y(_08047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11087_ (.A(_08047_),
    .X(_08048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11088_ (.A(_08046_),
    .X(_08049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11089_ (.A1(_00196_),
    .A2(_08048_),
    .B1(\design_top.MEM[11][7] ),
    .B2(_08049_),
    .X(_04461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11090_ (.A1(_00195_),
    .A2(_08048_),
    .B1(\design_top.MEM[11][6] ),
    .B2(_08049_),
    .X(_04460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11091_ (.A1(_00194_),
    .A2(_08048_),
    .B1(\design_top.MEM[11][5] ),
    .B2(_08049_),
    .X(_04459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11092_ (.A1(_00193_),
    .A2(_08048_),
    .B1(\design_top.MEM[11][4] ),
    .B2(_08049_),
    .X(_04458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11093_ (.A1(_00192_),
    .A2(_08048_),
    .B1(\design_top.MEM[11][3] ),
    .B2(_08049_),
    .X(_04457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11094_ (.A1(_00191_),
    .A2(_08047_),
    .B1(\design_top.MEM[11][2] ),
    .B2(_08046_),
    .X(_04456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11095_ (.A1(_00190_),
    .A2(_08047_),
    .B1(\design_top.MEM[11][1] ),
    .B2(_08046_),
    .X(_04455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11096_ (.A1(_00189_),
    .A2(_08047_),
    .B1(\design_top.MEM[11][0] ),
    .B2(_08046_),
    .X(_04454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11097_ (.A(_07027_),
    .Y(_01375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11098_ (.A(io_out[14]),
    .Y(_08050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11099_ (.A1(_07027_),
    .A2(_08030_),
    .B1(io_out[14]),
    .X(_08051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _11100_ (.A1(_01375_),
    .A2(_08033_),
    .A3(_08050_),
    .B1(_08051_),
    .X(_04453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11101_ (.A1(_06977_),
    .A2(_07067_),
    .B1(_07060_),
    .B2(_08023_),
    .X(_08052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11102_ (.A(_08052_),
    .Y(_08053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11103_ (.A(_08053_),
    .X(_08054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11104_ (.A(_08052_),
    .X(_08055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11105_ (.A1(_00364_),
    .A2(_08054_),
    .B1(\design_top.MEM[30][7] ),
    .B2(_08055_),
    .X(_04452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11106_ (.A1(_00363_),
    .A2(_08054_),
    .B1(\design_top.MEM[30][6] ),
    .B2(_08055_),
    .X(_04451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11107_ (.A1(_00362_),
    .A2(_08054_),
    .B1(\design_top.MEM[30][5] ),
    .B2(_08055_),
    .X(_04450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11108_ (.A1(_00361_),
    .A2(_08054_),
    .B1(\design_top.MEM[30][4] ),
    .B2(_08055_),
    .X(_04449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11109_ (.A1(_00360_),
    .A2(_08054_),
    .B1(\design_top.MEM[30][3] ),
    .B2(_08055_),
    .X(_04448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11110_ (.A1(_00359_),
    .A2(_08053_),
    .B1(\design_top.MEM[30][2] ),
    .B2(_08052_),
    .X(_04447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11111_ (.A1(_00358_),
    .A2(_08053_),
    .B1(\design_top.MEM[30][1] ),
    .B2(_08052_),
    .X(_04446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11112_ (.A1(_00357_),
    .A2(_08053_),
    .B1(\design_top.MEM[30][0] ),
    .B2(_08052_),
    .X(_04445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11113_ (.A1(_07048_),
    .A2(_07066_),
    .B1(_07080_),
    .B2(_08023_),
    .X(_08056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11114_ (.A(_08056_),
    .Y(_08057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11115_ (.A(_08057_),
    .X(_08058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11116_ (.A(_08056_),
    .X(_08059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11117_ (.A1(_00372_),
    .A2(_08058_),
    .B1(\design_top.MEM[31][7] ),
    .B2(_08059_),
    .X(_04444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11118_ (.A1(_00371_),
    .A2(_08058_),
    .B1(\design_top.MEM[31][6] ),
    .B2(_08059_),
    .X(_04443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11119_ (.A1(_00370_),
    .A2(_08058_),
    .B1(\design_top.MEM[31][5] ),
    .B2(_08059_),
    .X(_04442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11120_ (.A1(_00369_),
    .A2(_08058_),
    .B1(\design_top.MEM[31][4] ),
    .B2(_08059_),
    .X(_04441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11121_ (.A1(_00368_),
    .A2(_08058_),
    .B1(\design_top.MEM[31][3] ),
    .B2(_08059_),
    .X(_04440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11122_ (.A1(_00367_),
    .A2(_08057_),
    .B1(\design_top.MEM[31][2] ),
    .B2(_08056_),
    .X(_04439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11123_ (.A1(_00366_),
    .A2(_08057_),
    .B1(\design_top.MEM[31][1] ),
    .B2(_08056_),
    .X(_04438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11124_ (.A1(_00365_),
    .A2(_08057_),
    .B1(\design_top.MEM[31][0] ),
    .B2(_08056_),
    .X(_04437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11125_ (.A1(_06904_),
    .A2(_07047_),
    .B1(_07105_),
    .B2(_08023_),
    .X(_08060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11126_ (.A(_08060_),
    .Y(_08061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11127_ (.A(_08061_),
    .X(_08062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11128_ (.A(_08060_),
    .X(_08063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11129_ (.A1(_00380_),
    .A2(_08062_),
    .B1(\design_top.MEM[3][7] ),
    .B2(_08063_),
    .X(_04436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11130_ (.A1(_00379_),
    .A2(_08062_),
    .B1(\design_top.MEM[3][6] ),
    .B2(_08063_),
    .X(_04435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11131_ (.A1(_00378_),
    .A2(_08062_),
    .B1(\design_top.MEM[3][5] ),
    .B2(_08063_),
    .X(_04434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11132_ (.A1(_00377_),
    .A2(_08062_),
    .B1(\design_top.MEM[3][4] ),
    .B2(_08063_),
    .X(_04433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11133_ (.A1(_00376_),
    .A2(_08062_),
    .B1(\design_top.MEM[3][3] ),
    .B2(_08063_),
    .X(_04432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11134_ (.A1(_00375_),
    .A2(_08061_),
    .B1(\design_top.MEM[3][2] ),
    .B2(_08060_),
    .X(_04431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11135_ (.A1(_00374_),
    .A2(_08061_),
    .B1(\design_top.MEM[3][1] ),
    .B2(_08060_),
    .X(_04430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11136_ (.A1(_00373_),
    .A2(_08061_),
    .B1(\design_top.MEM[3][0] ),
    .B2(_08060_),
    .X(_04429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11137_ (.A(_01600_),
    .Y(_08064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11138_ (.A(_08064_),
    .X(_08065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11139_ (.A(_01599_),
    .Y(_08066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11140_ (.A(_08066_),
    .X(_08067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11141_ (.A(_01602_),
    .Y(_08068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11142_ (.A(_08068_),
    .X(_08069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11143_ (.A(_01601_),
    .Y(_08070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11144_ (.A(_08070_),
    .X(_08071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11145_ (.A(_08065_),
    .B(_08067_),
    .C(_08069_),
    .D(_08071_),
    .X(_08072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11146_ (.A(\design_top.core0.XJALR ),
    .B(\design_top.core0.XJAL ),
    .C(\design_top.core0.XRCC ),
    .D(\design_top.core0.XMCC ),
    .X(_08073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11147_ (.A(\design_top.core0.XLCC ),
    .B(\design_top.core0.XAUIPC ),
    .C(\design_top.core0.XLUI ),
    .D(_08073_),
    .X(_08074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11148_ (.A(_01600_),
    .B(_01599_),
    .C(_01602_),
    .D(_01601_),
    .X(_08075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11149_ (.A(_08075_),
    .Y(_08076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _11150_ (.A1(_00786_),
    .A2(_08074_),
    .B1(_08076_),
    .Y(_08077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _11151_ (.A1(_06662_),
    .A2(_08077_),
    .B1(_07721_),
    .X(_08078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11152_ (.A(_08072_),
    .B(_08078_),
    .X(_08079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11153_ (.A(_08079_),
    .X(_08080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11154_ (.A(_08080_),
    .X(_08081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11155_ (.A(_08079_),
    .Y(_08082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11156_ (.A(_08082_),
    .X(_08083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11157_ (.A(_08083_),
    .X(_08084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11158_ (.A(\design_top.core0.XRES ),
    .B(_08076_),
    .X(_08085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11159_ (.A(_08085_),
    .X(_08086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11160_ (.A(_08086_),
    .X(_08087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11161_ (.A(_00781_),
    .B(_08087_),
    .Y(_08088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11162_ (.A(_08088_),
    .X(_08089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11163_ (.A1(\design_top.core0.REG1[15][31] ),
    .A2(_08081_),
    .B1(_08084_),
    .B2(_08089_),
    .X(_04428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11164_ (.A(_02467_),
    .B(_08087_),
    .Y(_08090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11165_ (.A(_08090_),
    .X(_08091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11166_ (.A1(\design_top.core0.REG1[15][30] ),
    .A2(_08081_),
    .B1(_08084_),
    .B2(_08091_),
    .X(_04427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11167_ (.A(_02446_),
    .B(_08087_),
    .Y(_08092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11168_ (.A(_08092_),
    .X(_08093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11169_ (.A1(\design_top.core0.REG1[15][29] ),
    .A2(_08081_),
    .B1(_08084_),
    .B2(_08093_),
    .X(_04426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11170_ (.A(_02425_),
    .B(_08087_),
    .Y(_08094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11171_ (.A(_08094_),
    .X(_08095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11172_ (.A1(\design_top.core0.REG1[15][28] ),
    .A2(_08081_),
    .B1(_08084_),
    .B2(_08095_),
    .X(_04425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11173_ (.A(_08080_),
    .X(_08096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11174_ (.A(_02403_),
    .B(_08087_),
    .Y(_08097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11175_ (.A(_08097_),
    .X(_08098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11176_ (.A1(\design_top.core0.REG1[15][27] ),
    .A2(_08096_),
    .B1(_08084_),
    .B2(_08098_),
    .X(_04424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11177_ (.A(_08083_),
    .X(_08099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11178_ (.A(_08086_),
    .X(_08100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11179_ (.A(_02382_),
    .B(_08100_),
    .Y(_08101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11180_ (.A(_08101_),
    .X(_08102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11181_ (.A1(\design_top.core0.REG1[15][26] ),
    .A2(_08096_),
    .B1(_08099_),
    .B2(_08102_),
    .X(_04423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11182_ (.A(_02360_),
    .B(_08100_),
    .Y(_08103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11183_ (.A(_08103_),
    .X(_08104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11184_ (.A1(\design_top.core0.REG1[15][25] ),
    .A2(_08096_),
    .B1(_08099_),
    .B2(_08104_),
    .X(_04422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11185_ (.A(_02339_),
    .B(_08100_),
    .Y(_08105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11186_ (.A(_08105_),
    .X(_08106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11187_ (.A1(\design_top.core0.REG1[15][24] ),
    .A2(_08096_),
    .B1(_08099_),
    .B2(_08106_),
    .X(_04421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11188_ (.A(_02317_),
    .B(_08100_),
    .Y(_08107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11189_ (.A(_08107_),
    .X(_08108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11190_ (.A1(\design_top.core0.REG1[15][23] ),
    .A2(_08096_),
    .B1(_08099_),
    .B2(_08108_),
    .X(_04420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11191_ (.A(_08080_),
    .X(_08109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11192_ (.A(_02296_),
    .B(_08100_),
    .Y(_08110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11193_ (.A(_08110_),
    .X(_08111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11194_ (.A1(\design_top.core0.REG1[15][22] ),
    .A2(_08109_),
    .B1(_08099_),
    .B2(_08111_),
    .X(_04419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11195_ (.A(_08083_),
    .X(_08112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11196_ (.A(_08086_),
    .X(_08113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11197_ (.A(_02274_),
    .B(_08113_),
    .Y(_08114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11198_ (.A(_08114_),
    .X(_08115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11199_ (.A1(\design_top.core0.REG1[15][21] ),
    .A2(_08109_),
    .B1(_08112_),
    .B2(_08115_),
    .X(_04418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11200_ (.A(_02253_),
    .B(_08113_),
    .Y(_08116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11201_ (.A(_08116_),
    .X(_08117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11202_ (.A1(\design_top.core0.REG1[15][20] ),
    .A2(_08109_),
    .B1(_08112_),
    .B2(_08117_),
    .X(_04417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11203_ (.A(_02231_),
    .B(_08113_),
    .Y(_08118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11204_ (.A(_08118_),
    .X(_08119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11205_ (.A1(\design_top.core0.REG1[15][19] ),
    .A2(_08109_),
    .B1(_08112_),
    .B2(_08119_),
    .X(_04416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11206_ (.A(_02210_),
    .B(_08113_),
    .Y(_08120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11207_ (.A(_08120_),
    .X(_08121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11208_ (.A1(\design_top.core0.REG1[15][18] ),
    .A2(_08109_),
    .B1(_08112_),
    .B2(_08121_),
    .X(_04415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11209_ (.A(_08079_),
    .X(_08122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11210_ (.A(_02188_),
    .B(_08113_),
    .Y(_08123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11211_ (.A(_08123_),
    .X(_08124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11212_ (.A1(\design_top.core0.REG1[15][17] ),
    .A2(_08122_),
    .B1(_08112_),
    .B2(_08124_),
    .X(_04414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11213_ (.A(_08082_),
    .X(_08125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11214_ (.A(_08086_),
    .X(_08126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11215_ (.A(_02167_),
    .B(_08126_),
    .Y(_08127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11216_ (.A(_08127_),
    .X(_08128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11217_ (.A1(\design_top.core0.REG1[15][16] ),
    .A2(_08122_),
    .B1(_08125_),
    .B2(_08128_),
    .X(_04413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11218_ (.A(_02144_),
    .B(_08126_),
    .Y(_08129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11219_ (.A(_08129_),
    .X(_08130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11220_ (.A1(\design_top.core0.REG1[15][15] ),
    .A2(_08122_),
    .B1(_08125_),
    .B2(_08130_),
    .X(_04412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11221_ (.A(_02122_),
    .B(_08126_),
    .Y(_08131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11222_ (.A(_08131_),
    .X(_08132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11223_ (.A1(\design_top.core0.REG1[15][14] ),
    .A2(_08122_),
    .B1(_08125_),
    .B2(_08132_),
    .X(_04411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11224_ (.A(_00045_),
    .X(_08133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11225_ (.A1(\design_top.core0.REG1[15][13] ),
    .A2(_08083_),
    .B1(_08133_),
    .B2(_08081_),
    .X(_04410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11226_ (.A(_02073_),
    .B(_08126_),
    .Y(_08134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11227_ (.A(_08134_),
    .X(_08135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11228_ (.A1(\design_top.core0.REG1[15][12] ),
    .A2(_08122_),
    .B1(_08125_),
    .B2(_08135_),
    .X(_04409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11229_ (.A(_08079_),
    .X(_08136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11230_ (.A(_02049_),
    .B(_08126_),
    .Y(_08137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11231_ (.A(_08137_),
    .X(_08138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11232_ (.A1(\design_top.core0.REG1[15][11] ),
    .A2(_08136_),
    .B1(_08125_),
    .B2(_08138_),
    .X(_04408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11233_ (.A(_08082_),
    .X(_08139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11234_ (.A(_08085_),
    .X(_08140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11235_ (.A(_02026_),
    .B(_08140_),
    .Y(_08141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11236_ (.A(_08141_),
    .X(_08142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11237_ (.A1(\design_top.core0.REG1[15][10] ),
    .A2(_08136_),
    .B1(_08139_),
    .B2(_08142_),
    .X(_04407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11238_ (.A(_02002_),
    .B(_08140_),
    .Y(_08143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11239_ (.A(_08143_),
    .X(_08144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11240_ (.A1(\design_top.core0.REG1[15][9] ),
    .A2(_08136_),
    .B1(_08139_),
    .B2(_08144_),
    .X(_04406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11241_ (.A(_01979_),
    .B(_08140_),
    .Y(_08145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11242_ (.A(_08145_),
    .X(_08146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11243_ (.A1(\design_top.core0.REG1[15][8] ),
    .A2(_08136_),
    .B1(_08139_),
    .B2(_08146_),
    .X(_04405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11244_ (.A(_01954_),
    .B(_08140_),
    .Y(_08147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11245_ (.A(_08147_),
    .X(_08148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11246_ (.A1(\design_top.core0.REG1[15][7] ),
    .A2(_08136_),
    .B1(_08139_),
    .B2(_08148_),
    .X(_04404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11247_ (.A(_08079_),
    .X(_08149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11248_ (.A(_01911_),
    .B(_08140_),
    .Y(_08150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11249_ (.A(_08150_),
    .X(_08151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11250_ (.A1(\design_top.core0.REG1[15][6] ),
    .A2(_08149_),
    .B1(_08139_),
    .B2(_08151_),
    .X(_04403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11251_ (.A(_08082_),
    .X(_08152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11252_ (.A(_08085_),
    .X(_08153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11253_ (.A(_01866_),
    .B(_08153_),
    .Y(_08154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11254_ (.A(_08154_),
    .X(_08155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11255_ (.A1(\design_top.core0.REG1[15][5] ),
    .A2(_08149_),
    .B1(_08152_),
    .B2(_08155_),
    .X(_04402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11256_ (.A(_01822_),
    .B(_08153_),
    .Y(_08156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11257_ (.A(_08156_),
    .X(_08157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11258_ (.A1(\design_top.core0.REG1[15][4] ),
    .A2(_08149_),
    .B1(_08152_),
    .B2(_08157_),
    .X(_04401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11259_ (.A(_01778_),
    .B(_08153_),
    .Y(_08158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11260_ (.A(_08158_),
    .X(_08159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11261_ (.A1(\design_top.core0.REG1[15][3] ),
    .A2(_08149_),
    .B1(_08152_),
    .B2(_08159_),
    .X(_04400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11262_ (.A(_01727_),
    .B(_08153_),
    .Y(_08160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11263_ (.A(_08160_),
    .X(_08161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11264_ (.A1(\design_top.core0.REG1[15][2] ),
    .A2(_08149_),
    .B1(_08152_),
    .B2(_08161_),
    .X(_04399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11265_ (.A(_01673_),
    .B(_08153_),
    .Y(_08162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11266_ (.A(_08162_),
    .X(_08163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11267_ (.A1(\design_top.core0.REG1[15][1] ),
    .A2(_08080_),
    .B1(_08152_),
    .B2(_08163_),
    .X(_04398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11268_ (.A(_01598_),
    .B(_08086_),
    .Y(_08164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11269_ (.A(_08164_),
    .X(_08165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11270_ (.A1(\design_top.core0.REG1[15][0] ),
    .A2(_08080_),
    .B1(_08083_),
    .B2(_08165_),
    .X(_04397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11271_ (.A(_08078_),
    .X(_08166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11272_ (.A(_01602_),
    .X(_08167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11273_ (.A(_01601_),
    .X(_08168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11274_ (.A(_01600_),
    .X(_08169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11275_ (.A(_08167_),
    .B(_08168_),
    .C(_08169_),
    .D(_08066_),
    .X(_08170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11276_ (.A(_08166_),
    .B(_08170_),
    .X(_08171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11277_ (.A(_08171_),
    .X(_08172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11278_ (.A(_08172_),
    .X(_08173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11279_ (.A(_08088_),
    .X(_08174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11280_ (.A(_08174_),
    .X(_08175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11281_ (.A(_08171_),
    .Y(_08176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11282_ (.A(_08176_),
    .X(_08177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11283_ (.A(_08177_),
    .X(_08178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11284_ (.A1(\design_top.core0.REG1[1][31] ),
    .A2(_08173_),
    .B1(_08175_),
    .B2(_08178_),
    .X(_04396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11285_ (.A(_08090_),
    .X(_08179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11286_ (.A(_08179_),
    .X(_08180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11287_ (.A1(\design_top.core0.REG1[1][30] ),
    .A2(_08173_),
    .B1(_08180_),
    .B2(_08178_),
    .X(_04395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11288_ (.A(_08092_),
    .X(_08181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11289_ (.A(_08181_),
    .X(_08182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11290_ (.A1(\design_top.core0.REG1[1][29] ),
    .A2(_08173_),
    .B1(_08182_),
    .B2(_08178_),
    .X(_04394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11291_ (.A(_08094_),
    .X(_08183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11292_ (.A(_08183_),
    .X(_08184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11293_ (.A1(\design_top.core0.REG1[1][28] ),
    .A2(_08173_),
    .B1(_08184_),
    .B2(_08178_),
    .X(_04393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11294_ (.A(_08172_),
    .X(_08185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11295_ (.A(_08097_),
    .X(_08186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11296_ (.A(_08186_),
    .X(_08187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11297_ (.A1(\design_top.core0.REG1[1][27] ),
    .A2(_08185_),
    .B1(_08187_),
    .B2(_08178_),
    .X(_04392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11298_ (.A(_08101_),
    .X(_08188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11299_ (.A(_08188_),
    .X(_08189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11300_ (.A(_08177_),
    .X(_08190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11301_ (.A1(\design_top.core0.REG1[1][26] ),
    .A2(_08185_),
    .B1(_08189_),
    .B2(_08190_),
    .X(_04391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11302_ (.A(_08103_),
    .X(_08191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11303_ (.A(_08191_),
    .X(_08192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11304_ (.A1(\design_top.core0.REG1[1][25] ),
    .A2(_08185_),
    .B1(_08192_),
    .B2(_08190_),
    .X(_04390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11305_ (.A(_08105_),
    .X(_08193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11306_ (.A(_08193_),
    .X(_08194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11307_ (.A1(\design_top.core0.REG1[1][24] ),
    .A2(_08185_),
    .B1(_08194_),
    .B2(_08190_),
    .X(_04389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11308_ (.A(_08107_),
    .X(_08195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11309_ (.A(_08195_),
    .X(_08196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11310_ (.A1(\design_top.core0.REG1[1][23] ),
    .A2(_08185_),
    .B1(_08196_),
    .B2(_08190_),
    .X(_04388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11311_ (.A(_08172_),
    .X(_08197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11312_ (.A(_08110_),
    .X(_08198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11313_ (.A(_08198_),
    .X(_08199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11314_ (.A1(\design_top.core0.REG1[1][22] ),
    .A2(_08197_),
    .B1(_08199_),
    .B2(_08190_),
    .X(_04387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11315_ (.A(_08114_),
    .X(_08200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11316_ (.A(_08200_),
    .X(_08201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11317_ (.A(_08177_),
    .X(_08202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11318_ (.A1(\design_top.core0.REG1[1][21] ),
    .A2(_08197_),
    .B1(_08201_),
    .B2(_08202_),
    .X(_04386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11319_ (.A(_08116_),
    .X(_08203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11320_ (.A(_08203_),
    .X(_08204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11321_ (.A1(\design_top.core0.REG1[1][20] ),
    .A2(_08197_),
    .B1(_08204_),
    .B2(_08202_),
    .X(_04385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11322_ (.A(_08118_),
    .X(_08205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11323_ (.A(_08205_),
    .X(_08206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11324_ (.A1(\design_top.core0.REG1[1][19] ),
    .A2(_08197_),
    .B1(_08206_),
    .B2(_08202_),
    .X(_04384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11325_ (.A(_08120_),
    .X(_08207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11326_ (.A(_08207_),
    .X(_08208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11327_ (.A1(\design_top.core0.REG1[1][18] ),
    .A2(_08197_),
    .B1(_08208_),
    .B2(_08202_),
    .X(_04383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11328_ (.A(_08171_),
    .X(_08209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11329_ (.A(_08123_),
    .X(_08210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11330_ (.A(_08210_),
    .X(_08211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11331_ (.A1(\design_top.core0.REG1[1][17] ),
    .A2(_08209_),
    .B1(_08211_),
    .B2(_08202_),
    .X(_04382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11332_ (.A(_08127_),
    .X(_08212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11333_ (.A(_08212_),
    .X(_08213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11334_ (.A(_08176_),
    .X(_08214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11335_ (.A1(\design_top.core0.REG1[1][16] ),
    .A2(_08209_),
    .B1(_08213_),
    .B2(_08214_),
    .X(_04381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11336_ (.A(_08129_),
    .X(_08215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11337_ (.A(_08215_),
    .X(_08216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11338_ (.A1(\design_top.core0.REG1[1][15] ),
    .A2(_08209_),
    .B1(_08216_),
    .B2(_08214_),
    .X(_04380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11339_ (.A(_08131_),
    .X(_08217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11340_ (.A(_08217_),
    .X(_08218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11341_ (.A1(\design_top.core0.REG1[1][14] ),
    .A2(_08209_),
    .B1(_08218_),
    .B2(_08214_),
    .X(_04379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11342_ (.A1(\design_top.core0.REG1[1][13] ),
    .A2(_08177_),
    .B1(_08133_),
    .B2(_08173_),
    .X(_04378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11343_ (.A(_08134_),
    .X(_08219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11344_ (.A(_08219_),
    .X(_08220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11345_ (.A1(\design_top.core0.REG1[1][12] ),
    .A2(_08209_),
    .B1(_08220_),
    .B2(_08214_),
    .X(_04377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11346_ (.A(_08171_),
    .X(_08221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11347_ (.A(_08137_),
    .X(_08222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11348_ (.A(_08222_),
    .X(_08223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11349_ (.A1(\design_top.core0.REG1[1][11] ),
    .A2(_08221_),
    .B1(_08223_),
    .B2(_08214_),
    .X(_04376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11350_ (.A(_08141_),
    .X(_08224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11351_ (.A(_08224_),
    .X(_08225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11352_ (.A(_08176_),
    .X(_08226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11353_ (.A1(\design_top.core0.REG1[1][10] ),
    .A2(_08221_),
    .B1(_08225_),
    .B2(_08226_),
    .X(_04375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11354_ (.A(_08143_),
    .X(_08227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11355_ (.A(_08227_),
    .X(_08228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11356_ (.A1(\design_top.core0.REG1[1][9] ),
    .A2(_08221_),
    .B1(_08228_),
    .B2(_08226_),
    .X(_04374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11357_ (.A(_08145_),
    .X(_08229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11358_ (.A(_08229_),
    .X(_08230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11359_ (.A1(\design_top.core0.REG1[1][8] ),
    .A2(_08221_),
    .B1(_08230_),
    .B2(_08226_),
    .X(_04373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11360_ (.A(_08147_),
    .X(_08231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11361_ (.A(_08231_),
    .X(_08232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11362_ (.A1(\design_top.core0.REG1[1][7] ),
    .A2(_08221_),
    .B1(_08232_),
    .B2(_08226_),
    .X(_04372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11363_ (.A(_08171_),
    .X(_08233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11364_ (.A(_08150_),
    .X(_08234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11365_ (.A(_08234_),
    .X(_08235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11366_ (.A1(\design_top.core0.REG1[1][6] ),
    .A2(_08233_),
    .B1(_08235_),
    .B2(_08226_),
    .X(_04371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11367_ (.A(_08154_),
    .X(_08236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11368_ (.A(_08236_),
    .X(_08237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11369_ (.A(_08176_),
    .X(_08238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11370_ (.A1(\design_top.core0.REG1[1][5] ),
    .A2(_08233_),
    .B1(_08237_),
    .B2(_08238_),
    .X(_04370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11371_ (.A(_08156_),
    .X(_08239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11372_ (.A(_08239_),
    .X(_08240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11373_ (.A1(\design_top.core0.REG1[1][4] ),
    .A2(_08233_),
    .B1(_08240_),
    .B2(_08238_),
    .X(_04369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11374_ (.A(_08158_),
    .X(_08241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11375_ (.A(_08241_),
    .X(_08242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11376_ (.A1(\design_top.core0.REG1[1][3] ),
    .A2(_08233_),
    .B1(_08242_),
    .B2(_08238_),
    .X(_04368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11377_ (.A(_08160_),
    .X(_08243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11378_ (.A(_08243_),
    .X(_08244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11379_ (.A1(\design_top.core0.REG1[1][2] ),
    .A2(_08233_),
    .B1(_08244_),
    .B2(_08238_),
    .X(_04367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11380_ (.A(_08162_),
    .X(_08245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11381_ (.A(_08245_),
    .X(_08246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11382_ (.A1(\design_top.core0.REG1[1][1] ),
    .A2(_08172_),
    .B1(_08246_),
    .B2(_08238_),
    .X(_04366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11383_ (.A(_08164_),
    .X(_08247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11384_ (.A(_08247_),
    .X(_08248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11385_ (.A1(\design_top.core0.REG1[1][0] ),
    .A2(_08172_),
    .B1(_08248_),
    .B2(_08177_),
    .X(_04365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11386_ (.A(_01599_),
    .X(_08249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11387_ (.A(_08167_),
    .B(_08168_),
    .C(_08064_),
    .D(_08249_),
    .X(_08250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11388_ (.A(_08166_),
    .B(_08250_),
    .X(_08251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11389_ (.A(_08251_),
    .X(_08252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11390_ (.A(_08252_),
    .X(_08253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11391_ (.A(_08251_),
    .Y(_08254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11392_ (.A(_08254_),
    .X(_08255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11393_ (.A(_08255_),
    .X(_08256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11394_ (.A1(\design_top.core0.REG1[2][31] ),
    .A2(_08253_),
    .B1(_08175_),
    .B2(_08256_),
    .X(_04364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11395_ (.A1(\design_top.core0.REG1[2][30] ),
    .A2(_08253_),
    .B1(_08180_),
    .B2(_08256_),
    .X(_04363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11396_ (.A1(\design_top.core0.REG1[2][29] ),
    .A2(_08253_),
    .B1(_08182_),
    .B2(_08256_),
    .X(_04362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11397_ (.A1(\design_top.core0.REG1[2][28] ),
    .A2(_08253_),
    .B1(_08184_),
    .B2(_08256_),
    .X(_04361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11398_ (.A(_08252_),
    .X(_08257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11399_ (.A1(\design_top.core0.REG1[2][27] ),
    .A2(_08257_),
    .B1(_08187_),
    .B2(_08256_),
    .X(_04360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11400_ (.A(_08255_),
    .X(_08258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11401_ (.A1(\design_top.core0.REG1[2][26] ),
    .A2(_08257_),
    .B1(_08189_),
    .B2(_08258_),
    .X(_04359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11402_ (.A1(\design_top.core0.REG1[2][25] ),
    .A2(_08257_),
    .B1(_08192_),
    .B2(_08258_),
    .X(_04358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11403_ (.A1(\design_top.core0.REG1[2][24] ),
    .A2(_08257_),
    .B1(_08194_),
    .B2(_08258_),
    .X(_04357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11404_ (.A1(\design_top.core0.REG1[2][23] ),
    .A2(_08257_),
    .B1(_08196_),
    .B2(_08258_),
    .X(_04356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11405_ (.A(_08252_),
    .X(_08259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11406_ (.A1(\design_top.core0.REG1[2][22] ),
    .A2(_08259_),
    .B1(_08199_),
    .B2(_08258_),
    .X(_04355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11407_ (.A(_08255_),
    .X(_08260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11408_ (.A1(\design_top.core0.REG1[2][21] ),
    .A2(_08259_),
    .B1(_08201_),
    .B2(_08260_),
    .X(_04354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11409_ (.A1(\design_top.core0.REG1[2][20] ),
    .A2(_08259_),
    .B1(_08204_),
    .B2(_08260_),
    .X(_04353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11410_ (.A1(\design_top.core0.REG1[2][19] ),
    .A2(_08259_),
    .B1(_08206_),
    .B2(_08260_),
    .X(_04352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11411_ (.A1(\design_top.core0.REG1[2][18] ),
    .A2(_08259_),
    .B1(_08208_),
    .B2(_08260_),
    .X(_04351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11412_ (.A(_08251_),
    .X(_08261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11413_ (.A1(\design_top.core0.REG1[2][17] ),
    .A2(_08261_),
    .B1(_08211_),
    .B2(_08260_),
    .X(_04350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11414_ (.A(_08254_),
    .X(_08262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11415_ (.A1(\design_top.core0.REG1[2][16] ),
    .A2(_08261_),
    .B1(_08213_),
    .B2(_08262_),
    .X(_04349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11416_ (.A1(\design_top.core0.REG1[2][15] ),
    .A2(_08261_),
    .B1(_08216_),
    .B2(_08262_),
    .X(_04348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11417_ (.A1(\design_top.core0.REG1[2][14] ),
    .A2(_08261_),
    .B1(_08218_),
    .B2(_08262_),
    .X(_04347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11418_ (.A1(\design_top.core0.REG1[2][13] ),
    .A2(_08255_),
    .B1(_08133_),
    .B2(_08253_),
    .X(_04346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11419_ (.A1(\design_top.core0.REG1[2][12] ),
    .A2(_08261_),
    .B1(_08220_),
    .B2(_08262_),
    .X(_04345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11420_ (.A(_08251_),
    .X(_08263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11421_ (.A1(\design_top.core0.REG1[2][11] ),
    .A2(_08263_),
    .B1(_08223_),
    .B2(_08262_),
    .X(_04344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11422_ (.A(_08254_),
    .X(_08264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11423_ (.A1(\design_top.core0.REG1[2][10] ),
    .A2(_08263_),
    .B1(_08225_),
    .B2(_08264_),
    .X(_04343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11424_ (.A1(\design_top.core0.REG1[2][9] ),
    .A2(_08263_),
    .B1(_08228_),
    .B2(_08264_),
    .X(_04342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11425_ (.A1(\design_top.core0.REG1[2][8] ),
    .A2(_08263_),
    .B1(_08230_),
    .B2(_08264_),
    .X(_04341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11426_ (.A1(\design_top.core0.REG1[2][7] ),
    .A2(_08263_),
    .B1(_08232_),
    .B2(_08264_),
    .X(_04340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11427_ (.A(_08251_),
    .X(_08265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11428_ (.A1(\design_top.core0.REG1[2][6] ),
    .A2(_08265_),
    .B1(_08235_),
    .B2(_08264_),
    .X(_04339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11429_ (.A(_08254_),
    .X(_08266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11430_ (.A1(\design_top.core0.REG1[2][5] ),
    .A2(_08265_),
    .B1(_08237_),
    .B2(_08266_),
    .X(_04338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11431_ (.A1(\design_top.core0.REG1[2][4] ),
    .A2(_08265_),
    .B1(_08240_),
    .B2(_08266_),
    .X(_04337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11432_ (.A1(\design_top.core0.REG1[2][3] ),
    .A2(_08265_),
    .B1(_08242_),
    .B2(_08266_),
    .X(_04336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11433_ (.A1(\design_top.core0.REG1[2][2] ),
    .A2(_08265_),
    .B1(_08244_),
    .B2(_08266_),
    .X(_04335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11434_ (.A1(\design_top.core0.REG1[2][1] ),
    .A2(_08252_),
    .B1(_08246_),
    .B2(_08266_),
    .X(_04334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11435_ (.A1(\design_top.core0.REG1[2][0] ),
    .A2(_08252_),
    .B1(_08248_),
    .B2(_08255_),
    .X(_04333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11436_ (.A(_08065_),
    .B(_08067_),
    .C(_08167_),
    .D(_08168_),
    .X(_08267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11437_ (.A(_08166_),
    .B(_08267_),
    .X(_08268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11438_ (.A(_08268_),
    .X(_08269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11439_ (.A(_08269_),
    .X(_08270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11440_ (.A(_08268_),
    .Y(_08271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11441_ (.A(_08271_),
    .X(_08272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11442_ (.A(_08272_),
    .X(_08273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11443_ (.A1(\design_top.core0.REG1[3][31] ),
    .A2(_08270_),
    .B1(_08175_),
    .B2(_08273_),
    .X(_04332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11444_ (.A1(\design_top.core0.REG1[3][30] ),
    .A2(_08270_),
    .B1(_08180_),
    .B2(_08273_),
    .X(_04331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11445_ (.A1(\design_top.core0.REG1[3][29] ),
    .A2(_08270_),
    .B1(_08182_),
    .B2(_08273_),
    .X(_04330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11446_ (.A1(\design_top.core0.REG1[3][28] ),
    .A2(_08270_),
    .B1(_08184_),
    .B2(_08273_),
    .X(_04329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11447_ (.A(_08269_),
    .X(_08274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11448_ (.A1(\design_top.core0.REG1[3][27] ),
    .A2(_08274_),
    .B1(_08187_),
    .B2(_08273_),
    .X(_04328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11449_ (.A(_08272_),
    .X(_08275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11450_ (.A1(\design_top.core0.REG1[3][26] ),
    .A2(_08274_),
    .B1(_08189_),
    .B2(_08275_),
    .X(_04327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11451_ (.A1(\design_top.core0.REG1[3][25] ),
    .A2(_08274_),
    .B1(_08192_),
    .B2(_08275_),
    .X(_04326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11452_ (.A1(\design_top.core0.REG1[3][24] ),
    .A2(_08274_),
    .B1(_08194_),
    .B2(_08275_),
    .X(_04325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11453_ (.A1(\design_top.core0.REG1[3][23] ),
    .A2(_08274_),
    .B1(_08196_),
    .B2(_08275_),
    .X(_04324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11454_ (.A(_08269_),
    .X(_08276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11455_ (.A1(\design_top.core0.REG1[3][22] ),
    .A2(_08276_),
    .B1(_08199_),
    .B2(_08275_),
    .X(_04323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11456_ (.A(_08272_),
    .X(_08277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11457_ (.A1(\design_top.core0.REG1[3][21] ),
    .A2(_08276_),
    .B1(_08201_),
    .B2(_08277_),
    .X(_04322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11458_ (.A1(\design_top.core0.REG1[3][20] ),
    .A2(_08276_),
    .B1(_08204_),
    .B2(_08277_),
    .X(_04321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11459_ (.A1(\design_top.core0.REG1[3][19] ),
    .A2(_08276_),
    .B1(_08206_),
    .B2(_08277_),
    .X(_04320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11460_ (.A1(\design_top.core0.REG1[3][18] ),
    .A2(_08276_),
    .B1(_08208_),
    .B2(_08277_),
    .X(_04319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11461_ (.A(_08268_),
    .X(_08278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11462_ (.A1(\design_top.core0.REG1[3][17] ),
    .A2(_08278_),
    .B1(_08211_),
    .B2(_08277_),
    .X(_04318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11463_ (.A(_08271_),
    .X(_08279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11464_ (.A1(\design_top.core0.REG1[3][16] ),
    .A2(_08278_),
    .B1(_08213_),
    .B2(_08279_),
    .X(_04317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11465_ (.A1(\design_top.core0.REG1[3][15] ),
    .A2(_08278_),
    .B1(_08216_),
    .B2(_08279_),
    .X(_04316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11466_ (.A1(\design_top.core0.REG1[3][14] ),
    .A2(_08278_),
    .B1(_08218_),
    .B2(_08279_),
    .X(_04315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11467_ (.A1(\design_top.core0.REG1[3][13] ),
    .A2(_08272_),
    .B1(_08133_),
    .B2(_08270_),
    .X(_04314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11468_ (.A1(\design_top.core0.REG1[3][12] ),
    .A2(_08278_),
    .B1(_08220_),
    .B2(_08279_),
    .X(_04313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11469_ (.A(_08268_),
    .X(_08280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11470_ (.A1(\design_top.core0.REG1[3][11] ),
    .A2(_08280_),
    .B1(_08223_),
    .B2(_08279_),
    .X(_04312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11471_ (.A(_08271_),
    .X(_08281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11472_ (.A1(\design_top.core0.REG1[3][10] ),
    .A2(_08280_),
    .B1(_08225_),
    .B2(_08281_),
    .X(_04311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11473_ (.A1(\design_top.core0.REG1[3][9] ),
    .A2(_08280_),
    .B1(_08228_),
    .B2(_08281_),
    .X(_04310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11474_ (.A1(\design_top.core0.REG1[3][8] ),
    .A2(_08280_),
    .B1(_08230_),
    .B2(_08281_),
    .X(_04309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11475_ (.A1(\design_top.core0.REG1[3][7] ),
    .A2(_08280_),
    .B1(_08232_),
    .B2(_08281_),
    .X(_04308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11476_ (.A(_08268_),
    .X(_08282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11477_ (.A1(\design_top.core0.REG1[3][6] ),
    .A2(_08282_),
    .B1(_08235_),
    .B2(_08281_),
    .X(_04307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11478_ (.A(_08271_),
    .X(_08283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11479_ (.A1(\design_top.core0.REG1[3][5] ),
    .A2(_08282_),
    .B1(_08237_),
    .B2(_08283_),
    .X(_04306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11480_ (.A1(\design_top.core0.REG1[3][4] ),
    .A2(_08282_),
    .B1(_08240_),
    .B2(_08283_),
    .X(_04305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11481_ (.A1(\design_top.core0.REG1[3][3] ),
    .A2(_08282_),
    .B1(_08242_),
    .B2(_08283_),
    .X(_04304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11482_ (.A1(\design_top.core0.REG1[3][2] ),
    .A2(_08282_),
    .B1(_08244_),
    .B2(_08283_),
    .X(_04303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11483_ (.A1(\design_top.core0.REG1[3][1] ),
    .A2(_08269_),
    .B1(_08246_),
    .B2(_08283_),
    .X(_04302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11484_ (.A1(\design_top.core0.REG1[3][0] ),
    .A2(_08269_),
    .B1(_08248_),
    .B2(_08272_),
    .X(_04301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11485_ (.A(_08169_),
    .B(_08249_),
    .C(_08167_),
    .D(_08071_),
    .X(_08284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11486_ (.A(_08166_),
    .B(_08284_),
    .X(_08285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11487_ (.A(_08285_),
    .X(_08286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11488_ (.A(_08286_),
    .X(_08287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11489_ (.A(_08285_),
    .Y(_08288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11490_ (.A(_08288_),
    .X(_08289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11491_ (.A(_08289_),
    .X(_08290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11492_ (.A1(\design_top.core0.REG1[4][31] ),
    .A2(_08287_),
    .B1(_08175_),
    .B2(_08290_),
    .X(_04300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11493_ (.A1(\design_top.core0.REG1[4][30] ),
    .A2(_08287_),
    .B1(_08180_),
    .B2(_08290_),
    .X(_04299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11494_ (.A1(\design_top.core0.REG1[4][29] ),
    .A2(_08287_),
    .B1(_08182_),
    .B2(_08290_),
    .X(_04298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11495_ (.A1(\design_top.core0.REG1[4][28] ),
    .A2(_08287_),
    .B1(_08184_),
    .B2(_08290_),
    .X(_04297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11496_ (.A(_08286_),
    .X(_08291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11497_ (.A1(\design_top.core0.REG1[4][27] ),
    .A2(_08291_),
    .B1(_08187_),
    .B2(_08290_),
    .X(_04296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11498_ (.A(_08289_),
    .X(_08292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11499_ (.A1(\design_top.core0.REG1[4][26] ),
    .A2(_08291_),
    .B1(_08189_),
    .B2(_08292_),
    .X(_04295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11500_ (.A1(\design_top.core0.REG1[4][25] ),
    .A2(_08291_),
    .B1(_08192_),
    .B2(_08292_),
    .X(_04294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11501_ (.A1(\design_top.core0.REG1[4][24] ),
    .A2(_08291_),
    .B1(_08194_),
    .B2(_08292_),
    .X(_04293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11502_ (.A1(\design_top.core0.REG1[4][23] ),
    .A2(_08291_),
    .B1(_08196_),
    .B2(_08292_),
    .X(_04292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11503_ (.A(_08286_),
    .X(_08293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11504_ (.A1(\design_top.core0.REG1[4][22] ),
    .A2(_08293_),
    .B1(_08199_),
    .B2(_08292_),
    .X(_04291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11505_ (.A(_08289_),
    .X(_08294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11506_ (.A1(\design_top.core0.REG1[4][21] ),
    .A2(_08293_),
    .B1(_08201_),
    .B2(_08294_),
    .X(_04290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11507_ (.A1(\design_top.core0.REG1[4][20] ),
    .A2(_08293_),
    .B1(_08204_),
    .B2(_08294_),
    .X(_04289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11508_ (.A1(\design_top.core0.REG1[4][19] ),
    .A2(_08293_),
    .B1(_08206_),
    .B2(_08294_),
    .X(_04288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11509_ (.A1(\design_top.core0.REG1[4][18] ),
    .A2(_08293_),
    .B1(_08208_),
    .B2(_08294_),
    .X(_04287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11510_ (.A(_08285_),
    .X(_08295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11511_ (.A1(\design_top.core0.REG1[4][17] ),
    .A2(_08295_),
    .B1(_08211_),
    .B2(_08294_),
    .X(_04286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11512_ (.A(_08288_),
    .X(_08296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11513_ (.A1(\design_top.core0.REG1[4][16] ),
    .A2(_08295_),
    .B1(_08213_),
    .B2(_08296_),
    .X(_04285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11514_ (.A1(\design_top.core0.REG1[4][15] ),
    .A2(_08295_),
    .B1(_08216_),
    .B2(_08296_),
    .X(_04284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11515_ (.A1(\design_top.core0.REG1[4][14] ),
    .A2(_08295_),
    .B1(_08218_),
    .B2(_08296_),
    .X(_04283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11516_ (.A(_00045_),
    .X(_08297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11517_ (.A1(\design_top.core0.REG1[4][13] ),
    .A2(_08289_),
    .B1(_08297_),
    .B2(_08287_),
    .X(_04282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11518_ (.A1(\design_top.core0.REG1[4][12] ),
    .A2(_08295_),
    .B1(_08220_),
    .B2(_08296_),
    .X(_04281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11519_ (.A(_08285_),
    .X(_08298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11520_ (.A1(\design_top.core0.REG1[4][11] ),
    .A2(_08298_),
    .B1(_08223_),
    .B2(_08296_),
    .X(_04280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11521_ (.A(_08288_),
    .X(_08299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11522_ (.A1(\design_top.core0.REG1[4][10] ),
    .A2(_08298_),
    .B1(_08225_),
    .B2(_08299_),
    .X(_04279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11523_ (.A1(\design_top.core0.REG1[4][9] ),
    .A2(_08298_),
    .B1(_08228_),
    .B2(_08299_),
    .X(_04278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11524_ (.A1(\design_top.core0.REG1[4][8] ),
    .A2(_08298_),
    .B1(_08230_),
    .B2(_08299_),
    .X(_04277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11525_ (.A1(\design_top.core0.REG1[4][7] ),
    .A2(_08298_),
    .B1(_08232_),
    .B2(_08299_),
    .X(_04276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11526_ (.A(_08285_),
    .X(_08300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11527_ (.A1(\design_top.core0.REG1[4][6] ),
    .A2(_08300_),
    .B1(_08235_),
    .B2(_08299_),
    .X(_04275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11528_ (.A(_08288_),
    .X(_08301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11529_ (.A1(\design_top.core0.REG1[4][5] ),
    .A2(_08300_),
    .B1(_08237_),
    .B2(_08301_),
    .X(_04274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11530_ (.A1(\design_top.core0.REG1[4][4] ),
    .A2(_08300_),
    .B1(_08240_),
    .B2(_08301_),
    .X(_04273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11531_ (.A1(\design_top.core0.REG1[4][3] ),
    .A2(_08300_),
    .B1(_08242_),
    .B2(_08301_),
    .X(_04272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11532_ (.A1(\design_top.core0.REG1[4][2] ),
    .A2(_08300_),
    .B1(_08244_),
    .B2(_08301_),
    .X(_04271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11533_ (.A1(\design_top.core0.REG1[4][1] ),
    .A2(_08286_),
    .B1(_08246_),
    .B2(_08301_),
    .X(_04270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11534_ (.A1(\design_top.core0.REG1[4][0] ),
    .A2(_08286_),
    .B1(_08248_),
    .B2(_08289_),
    .X(_04269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11535_ (.A(_08078_),
    .X(_08302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11536_ (.A(_08169_),
    .B(_08067_),
    .C(_08167_),
    .D(_08070_),
    .X(_08303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11537_ (.A(_08302_),
    .B(_08303_),
    .X(_08304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11538_ (.A(_08304_),
    .X(_08305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11539_ (.A(_08305_),
    .X(_08306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11540_ (.A(_08304_),
    .Y(_08307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11541_ (.A(_08307_),
    .X(_08308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11542_ (.A(_08308_),
    .X(_08309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11543_ (.A1(\design_top.core0.REG1[5][31] ),
    .A2(_08306_),
    .B1(_08175_),
    .B2(_08309_),
    .X(_04268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11544_ (.A1(\design_top.core0.REG1[5][30] ),
    .A2(_08306_),
    .B1(_08180_),
    .B2(_08309_),
    .X(_04267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11545_ (.A1(\design_top.core0.REG1[5][29] ),
    .A2(_08306_),
    .B1(_08182_),
    .B2(_08309_),
    .X(_04266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11546_ (.A1(\design_top.core0.REG1[5][28] ),
    .A2(_08306_),
    .B1(_08184_),
    .B2(_08309_),
    .X(_04265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11547_ (.A(_08305_),
    .X(_08310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11548_ (.A1(\design_top.core0.REG1[5][27] ),
    .A2(_08310_),
    .B1(_08187_),
    .B2(_08309_),
    .X(_04264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11549_ (.A(_08308_),
    .X(_08311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11550_ (.A1(\design_top.core0.REG1[5][26] ),
    .A2(_08310_),
    .B1(_08189_),
    .B2(_08311_),
    .X(_04263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11551_ (.A1(\design_top.core0.REG1[5][25] ),
    .A2(_08310_),
    .B1(_08192_),
    .B2(_08311_),
    .X(_04262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11552_ (.A1(\design_top.core0.REG1[5][24] ),
    .A2(_08310_),
    .B1(_08194_),
    .B2(_08311_),
    .X(_04261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11553_ (.A1(\design_top.core0.REG1[5][23] ),
    .A2(_08310_),
    .B1(_08196_),
    .B2(_08311_),
    .X(_04260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11554_ (.A(_08305_),
    .X(_08312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11555_ (.A1(\design_top.core0.REG1[5][22] ),
    .A2(_08312_),
    .B1(_08199_),
    .B2(_08311_),
    .X(_04259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11556_ (.A(_08308_),
    .X(_08313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11557_ (.A1(\design_top.core0.REG1[5][21] ),
    .A2(_08312_),
    .B1(_08201_),
    .B2(_08313_),
    .X(_04258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11558_ (.A1(\design_top.core0.REG1[5][20] ),
    .A2(_08312_),
    .B1(_08204_),
    .B2(_08313_),
    .X(_04257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11559_ (.A1(\design_top.core0.REG1[5][19] ),
    .A2(_08312_),
    .B1(_08206_),
    .B2(_08313_),
    .X(_04256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11560_ (.A1(\design_top.core0.REG1[5][18] ),
    .A2(_08312_),
    .B1(_08208_),
    .B2(_08313_),
    .X(_04255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11561_ (.A(_08304_),
    .X(_08314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11562_ (.A1(\design_top.core0.REG1[5][17] ),
    .A2(_08314_),
    .B1(_08211_),
    .B2(_08313_),
    .X(_04254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11563_ (.A(_08307_),
    .X(_08315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11564_ (.A1(\design_top.core0.REG1[5][16] ),
    .A2(_08314_),
    .B1(_08213_),
    .B2(_08315_),
    .X(_04253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11565_ (.A1(\design_top.core0.REG1[5][15] ),
    .A2(_08314_),
    .B1(_08216_),
    .B2(_08315_),
    .X(_04252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11566_ (.A1(\design_top.core0.REG1[5][14] ),
    .A2(_08314_),
    .B1(_08218_),
    .B2(_08315_),
    .X(_04251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11567_ (.A1(\design_top.core0.REG1[5][13] ),
    .A2(_08308_),
    .B1(_08297_),
    .B2(_08306_),
    .X(_04250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11568_ (.A1(\design_top.core0.REG1[5][12] ),
    .A2(_08314_),
    .B1(_08220_),
    .B2(_08315_),
    .X(_04249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11569_ (.A(_08304_),
    .X(_08316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11570_ (.A1(\design_top.core0.REG1[5][11] ),
    .A2(_08316_),
    .B1(_08223_),
    .B2(_08315_),
    .X(_04248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11571_ (.A(_08307_),
    .X(_08317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11572_ (.A1(\design_top.core0.REG1[5][10] ),
    .A2(_08316_),
    .B1(_08225_),
    .B2(_08317_),
    .X(_04247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11573_ (.A1(\design_top.core0.REG1[5][9] ),
    .A2(_08316_),
    .B1(_08228_),
    .B2(_08317_),
    .X(_04246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11574_ (.A1(\design_top.core0.REG1[5][8] ),
    .A2(_08316_),
    .B1(_08230_),
    .B2(_08317_),
    .X(_04245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11575_ (.A1(\design_top.core0.REG1[5][7] ),
    .A2(_08316_),
    .B1(_08232_),
    .B2(_08317_),
    .X(_04244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11576_ (.A(_08304_),
    .X(_08318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11577_ (.A1(\design_top.core0.REG1[5][6] ),
    .A2(_08318_),
    .B1(_08235_),
    .B2(_08317_),
    .X(_04243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11578_ (.A(_08307_),
    .X(_08319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11579_ (.A1(\design_top.core0.REG1[5][5] ),
    .A2(_08318_),
    .B1(_08237_),
    .B2(_08319_),
    .X(_04242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11580_ (.A1(\design_top.core0.REG1[5][4] ),
    .A2(_08318_),
    .B1(_08240_),
    .B2(_08319_),
    .X(_04241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11581_ (.A1(\design_top.core0.REG1[5][3] ),
    .A2(_08318_),
    .B1(_08242_),
    .B2(_08319_),
    .X(_04240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11582_ (.A1(\design_top.core0.REG1[5][2] ),
    .A2(_08318_),
    .B1(_08244_),
    .B2(_08319_),
    .X(_04239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11583_ (.A1(\design_top.core0.REG1[5][1] ),
    .A2(_08305_),
    .B1(_08246_),
    .B2(_08319_),
    .X(_04238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11584_ (.A1(\design_top.core0.REG1[5][0] ),
    .A2(_08305_),
    .B1(_08248_),
    .B2(_08308_),
    .X(_04237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11585_ (.A(_08065_),
    .B(_08249_),
    .C(_01602_),
    .D(_08070_),
    .X(_08320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11586_ (.A(_08302_),
    .B(_08320_),
    .X(_08321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11587_ (.A(_08321_),
    .X(_08322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11588_ (.A(_08322_),
    .X(_08323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11589_ (.A(_08174_),
    .X(_08324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11590_ (.A(_08321_),
    .Y(_08325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11591_ (.A(_08325_),
    .X(_08326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11592_ (.A(_08326_),
    .X(_08327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11593_ (.A1(\design_top.core0.REG1[6][31] ),
    .A2(_08323_),
    .B1(_08324_),
    .B2(_08327_),
    .X(_04236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11594_ (.A(_08179_),
    .X(_08328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11595_ (.A1(\design_top.core0.REG1[6][30] ),
    .A2(_08323_),
    .B1(_08328_),
    .B2(_08327_),
    .X(_04235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11596_ (.A(_08181_),
    .X(_08329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11597_ (.A1(\design_top.core0.REG1[6][29] ),
    .A2(_08323_),
    .B1(_08329_),
    .B2(_08327_),
    .X(_04234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11598_ (.A(_08183_),
    .X(_08330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11599_ (.A1(\design_top.core0.REG1[6][28] ),
    .A2(_08323_),
    .B1(_08330_),
    .B2(_08327_),
    .X(_04233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11600_ (.A(_08322_),
    .X(_08331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11601_ (.A(_08186_),
    .X(_08332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11602_ (.A1(\design_top.core0.REG1[6][27] ),
    .A2(_08331_),
    .B1(_08332_),
    .B2(_08327_),
    .X(_04232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11603_ (.A(_08188_),
    .X(_08333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11604_ (.A(_08326_),
    .X(_08334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11605_ (.A1(\design_top.core0.REG1[6][26] ),
    .A2(_08331_),
    .B1(_08333_),
    .B2(_08334_),
    .X(_04231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11606_ (.A(_08191_),
    .X(_08335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11607_ (.A1(\design_top.core0.REG1[6][25] ),
    .A2(_08331_),
    .B1(_08335_),
    .B2(_08334_),
    .X(_04230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11608_ (.A(_08193_),
    .X(_08336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11609_ (.A1(\design_top.core0.REG1[6][24] ),
    .A2(_08331_),
    .B1(_08336_),
    .B2(_08334_),
    .X(_04229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11610_ (.A(_08195_),
    .X(_08337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11611_ (.A1(\design_top.core0.REG1[6][23] ),
    .A2(_08331_),
    .B1(_08337_),
    .B2(_08334_),
    .X(_04228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11612_ (.A(_08322_),
    .X(_08338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11613_ (.A(_08198_),
    .X(_08339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11614_ (.A1(\design_top.core0.REG1[6][22] ),
    .A2(_08338_),
    .B1(_08339_),
    .B2(_08334_),
    .X(_04227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11615_ (.A(_08200_),
    .X(_08340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11616_ (.A(_08326_),
    .X(_08341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11617_ (.A1(\design_top.core0.REG1[6][21] ),
    .A2(_08338_),
    .B1(_08340_),
    .B2(_08341_),
    .X(_04226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11618_ (.A(_08203_),
    .X(_08342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11619_ (.A1(\design_top.core0.REG1[6][20] ),
    .A2(_08338_),
    .B1(_08342_),
    .B2(_08341_),
    .X(_04225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11620_ (.A(_08205_),
    .X(_08343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11621_ (.A1(\design_top.core0.REG1[6][19] ),
    .A2(_08338_),
    .B1(_08343_),
    .B2(_08341_),
    .X(_04224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11622_ (.A(_08207_),
    .X(_08344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11623_ (.A1(\design_top.core0.REG1[6][18] ),
    .A2(_08338_),
    .B1(_08344_),
    .B2(_08341_),
    .X(_04223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11624_ (.A(_08321_),
    .X(_08345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11625_ (.A(_08210_),
    .X(_08346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11626_ (.A1(\design_top.core0.REG1[6][17] ),
    .A2(_08345_),
    .B1(_08346_),
    .B2(_08341_),
    .X(_04222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11627_ (.A(_08212_),
    .X(_08347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11628_ (.A(_08325_),
    .X(_08348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11629_ (.A1(\design_top.core0.REG1[6][16] ),
    .A2(_08345_),
    .B1(_08347_),
    .B2(_08348_),
    .X(_04221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11630_ (.A(_08215_),
    .X(_08349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11631_ (.A1(\design_top.core0.REG1[6][15] ),
    .A2(_08345_),
    .B1(_08349_),
    .B2(_08348_),
    .X(_04220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11632_ (.A(_08217_),
    .X(_08350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11633_ (.A1(\design_top.core0.REG1[6][14] ),
    .A2(_08345_),
    .B1(_08350_),
    .B2(_08348_),
    .X(_04219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11634_ (.A1(\design_top.core0.REG1[6][13] ),
    .A2(_08326_),
    .B1(_08297_),
    .B2(_08323_),
    .X(_04218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11635_ (.A(_08219_),
    .X(_08351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11636_ (.A1(\design_top.core0.REG1[6][12] ),
    .A2(_08345_),
    .B1(_08351_),
    .B2(_08348_),
    .X(_04217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11637_ (.A(_08321_),
    .X(_08352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11638_ (.A(_08222_),
    .X(_08353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11639_ (.A1(\design_top.core0.REG1[6][11] ),
    .A2(_08352_),
    .B1(_08353_),
    .B2(_08348_),
    .X(_04216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11640_ (.A(_08224_),
    .X(_08354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11641_ (.A(_08325_),
    .X(_08355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11642_ (.A1(\design_top.core0.REG1[6][10] ),
    .A2(_08352_),
    .B1(_08354_),
    .B2(_08355_),
    .X(_04215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11643_ (.A(_08227_),
    .X(_08356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11644_ (.A1(\design_top.core0.REG1[6][9] ),
    .A2(_08352_),
    .B1(_08356_),
    .B2(_08355_),
    .X(_04214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11645_ (.A(_08229_),
    .X(_08357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11646_ (.A1(\design_top.core0.REG1[6][8] ),
    .A2(_08352_),
    .B1(_08357_),
    .B2(_08355_),
    .X(_04213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11647_ (.A(_08231_),
    .X(_08358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11648_ (.A1(\design_top.core0.REG1[6][7] ),
    .A2(_08352_),
    .B1(_08358_),
    .B2(_08355_),
    .X(_04212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11649_ (.A(_08321_),
    .X(_08359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11650_ (.A(_08234_),
    .X(_08360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11651_ (.A1(\design_top.core0.REG1[6][6] ),
    .A2(_08359_),
    .B1(_08360_),
    .B2(_08355_),
    .X(_04211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11652_ (.A(_08236_),
    .X(_08361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11653_ (.A(_08325_),
    .X(_08362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11654_ (.A1(\design_top.core0.REG1[6][5] ),
    .A2(_08359_),
    .B1(_08361_),
    .B2(_08362_),
    .X(_04210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11655_ (.A(_08239_),
    .X(_08363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11656_ (.A1(\design_top.core0.REG1[6][4] ),
    .A2(_08359_),
    .B1(_08363_),
    .B2(_08362_),
    .X(_04209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11657_ (.A(_08241_),
    .X(_08364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11658_ (.A1(\design_top.core0.REG1[6][3] ),
    .A2(_08359_),
    .B1(_08364_),
    .B2(_08362_),
    .X(_04208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11659_ (.A(_08243_),
    .X(_08365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11660_ (.A1(\design_top.core0.REG1[6][2] ),
    .A2(_08359_),
    .B1(_08365_),
    .B2(_08362_),
    .X(_04207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11661_ (.A(_08245_),
    .X(_08366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11662_ (.A1(\design_top.core0.REG1[6][1] ),
    .A2(_08322_),
    .B1(_08366_),
    .B2(_08362_),
    .X(_04206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11663_ (.A(_08247_),
    .X(_08367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11664_ (.A1(\design_top.core0.REG1[6][0] ),
    .A2(_08322_),
    .B1(_08367_),
    .B2(_08326_),
    .X(_04205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11665_ (.A(_08065_),
    .B(_08067_),
    .C(_01602_),
    .D(_08070_),
    .X(_08368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11666_ (.A(_08302_),
    .B(_08368_),
    .X(_08369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11667_ (.A(_08369_),
    .X(_08370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11668_ (.A(_08370_),
    .X(_08371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11669_ (.A(_08369_),
    .Y(_08372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11670_ (.A(_08372_),
    .X(_08373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11671_ (.A(_08373_),
    .X(_08374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11672_ (.A1(\design_top.core0.REG1[7][31] ),
    .A2(_08371_),
    .B1(_08324_),
    .B2(_08374_),
    .X(_04204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11673_ (.A1(\design_top.core0.REG1[7][30] ),
    .A2(_08371_),
    .B1(_08328_),
    .B2(_08374_),
    .X(_04203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11674_ (.A1(\design_top.core0.REG1[7][29] ),
    .A2(_08371_),
    .B1(_08329_),
    .B2(_08374_),
    .X(_04202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11675_ (.A1(\design_top.core0.REG1[7][28] ),
    .A2(_08371_),
    .B1(_08330_),
    .B2(_08374_),
    .X(_04201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11676_ (.A(_08370_),
    .X(_08375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11677_ (.A1(\design_top.core0.REG1[7][27] ),
    .A2(_08375_),
    .B1(_08332_),
    .B2(_08374_),
    .X(_04200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11678_ (.A(_08373_),
    .X(_08376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11679_ (.A1(\design_top.core0.REG1[7][26] ),
    .A2(_08375_),
    .B1(_08333_),
    .B2(_08376_),
    .X(_04199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11680_ (.A1(\design_top.core0.REG1[7][25] ),
    .A2(_08375_),
    .B1(_08335_),
    .B2(_08376_),
    .X(_04198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11681_ (.A1(\design_top.core0.REG1[7][24] ),
    .A2(_08375_),
    .B1(_08336_),
    .B2(_08376_),
    .X(_04197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11682_ (.A1(\design_top.core0.REG1[7][23] ),
    .A2(_08375_),
    .B1(_08337_),
    .B2(_08376_),
    .X(_04196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11683_ (.A(_08370_),
    .X(_08377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11684_ (.A1(\design_top.core0.REG1[7][22] ),
    .A2(_08377_),
    .B1(_08339_),
    .B2(_08376_),
    .X(_04195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11685_ (.A(_08373_),
    .X(_08378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11686_ (.A1(\design_top.core0.REG1[7][21] ),
    .A2(_08377_),
    .B1(_08340_),
    .B2(_08378_),
    .X(_04194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11687_ (.A1(\design_top.core0.REG1[7][20] ),
    .A2(_08377_),
    .B1(_08342_),
    .B2(_08378_),
    .X(_04193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11688_ (.A1(\design_top.core0.REG1[7][19] ),
    .A2(_08377_),
    .B1(_08343_),
    .B2(_08378_),
    .X(_04192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11689_ (.A1(\design_top.core0.REG1[7][18] ),
    .A2(_08377_),
    .B1(_08344_),
    .B2(_08378_),
    .X(_04191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11690_ (.A(_08369_),
    .X(_08379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11691_ (.A1(\design_top.core0.REG1[7][17] ),
    .A2(_08379_),
    .B1(_08346_),
    .B2(_08378_),
    .X(_04190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11692_ (.A(_08372_),
    .X(_08380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11693_ (.A1(\design_top.core0.REG1[7][16] ),
    .A2(_08379_),
    .B1(_08347_),
    .B2(_08380_),
    .X(_04189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11694_ (.A1(\design_top.core0.REG1[7][15] ),
    .A2(_08379_),
    .B1(_08349_),
    .B2(_08380_),
    .X(_04188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11695_ (.A1(\design_top.core0.REG1[7][14] ),
    .A2(_08379_),
    .B1(_08350_),
    .B2(_08380_),
    .X(_04187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11696_ (.A1(\design_top.core0.REG1[7][13] ),
    .A2(_08373_),
    .B1(_08297_),
    .B2(_08371_),
    .X(_04186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11697_ (.A1(\design_top.core0.REG1[7][12] ),
    .A2(_08379_),
    .B1(_08351_),
    .B2(_08380_),
    .X(_04185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11698_ (.A(_08369_),
    .X(_08381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11699_ (.A1(\design_top.core0.REG1[7][11] ),
    .A2(_08381_),
    .B1(_08353_),
    .B2(_08380_),
    .X(_04184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11700_ (.A(_08372_),
    .X(_08382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11701_ (.A1(\design_top.core0.REG1[7][10] ),
    .A2(_08381_),
    .B1(_08354_),
    .B2(_08382_),
    .X(_04183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11702_ (.A1(\design_top.core0.REG1[7][9] ),
    .A2(_08381_),
    .B1(_08356_),
    .B2(_08382_),
    .X(_04182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11703_ (.A1(\design_top.core0.REG1[7][8] ),
    .A2(_08381_),
    .B1(_08357_),
    .B2(_08382_),
    .X(_04181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11704_ (.A1(\design_top.core0.REG1[7][7] ),
    .A2(_08381_),
    .B1(_08358_),
    .B2(_08382_),
    .X(_04180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11705_ (.A(_08369_),
    .X(_08383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11706_ (.A1(\design_top.core0.REG1[7][6] ),
    .A2(_08383_),
    .B1(_08360_),
    .B2(_08382_),
    .X(_04179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11707_ (.A(_08372_),
    .X(_08384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11708_ (.A1(\design_top.core0.REG1[7][5] ),
    .A2(_08383_),
    .B1(_08361_),
    .B2(_08384_),
    .X(_04178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11709_ (.A1(\design_top.core0.REG1[7][4] ),
    .A2(_08383_),
    .B1(_08363_),
    .B2(_08384_),
    .X(_04177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11710_ (.A1(\design_top.core0.REG1[7][3] ),
    .A2(_08383_),
    .B1(_08364_),
    .B2(_08384_),
    .X(_04176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11711_ (.A1(\design_top.core0.REG1[7][2] ),
    .A2(_08383_),
    .B1(_08365_),
    .B2(_08384_),
    .X(_04175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11712_ (.A1(\design_top.core0.REG1[7][1] ),
    .A2(_08370_),
    .B1(_08366_),
    .B2(_08384_),
    .X(_04174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11713_ (.A1(\design_top.core0.REG1[7][0] ),
    .A2(_08370_),
    .B1(_08367_),
    .B2(_08373_),
    .X(_04173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11714_ (.A(_08022_),
    .X(_08385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11715_ (.A1(_07150_),
    .A2(_07132_),
    .B1(_07128_),
    .B2(_08385_),
    .X(_08386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11716_ (.A(_08386_),
    .Y(_08387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11717_ (.A(_08387_),
    .X(_08388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11718_ (.A(_08386_),
    .X(_08389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11719_ (.A1(_00388_),
    .A2(_08388_),
    .B1(\design_top.MEM[4][7] ),
    .B2(_08389_),
    .X(_04172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11720_ (.A1(_00387_),
    .A2(_08388_),
    .B1(\design_top.MEM[4][6] ),
    .B2(_08389_),
    .X(_04171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11721_ (.A1(_00386_),
    .A2(_08388_),
    .B1(\design_top.MEM[4][5] ),
    .B2(_08389_),
    .X(_04170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11722_ (.A1(_00385_),
    .A2(_08388_),
    .B1(\design_top.MEM[4][4] ),
    .B2(_08389_),
    .X(_04169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11723_ (.A1(_00384_),
    .A2(_08388_),
    .B1(\design_top.MEM[4][3] ),
    .B2(_08389_),
    .X(_04168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11724_ (.A1(_00383_),
    .A2(_08387_),
    .B1(\design_top.MEM[4][2] ),
    .B2(_08386_),
    .X(_04167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11725_ (.A1(_00382_),
    .A2(_08387_),
    .B1(\design_top.MEM[4][1] ),
    .B2(_08386_),
    .X(_04166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11726_ (.A1(_00381_),
    .A2(_08387_),
    .B1(\design_top.MEM[4][0] ),
    .B2(_08386_),
    .X(_04165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11727_ (.A(_08169_),
    .B(_08249_),
    .C(_08069_),
    .D(_08168_),
    .X(_08390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11728_ (.A(_08302_),
    .B(_08390_),
    .X(_08391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11729_ (.A(_08391_),
    .X(_08392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11730_ (.A(_08392_),
    .X(_08393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11731_ (.A(_08391_),
    .Y(_08394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11732_ (.A(_08394_),
    .X(_08395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11733_ (.A(_08395_),
    .X(_08396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11734_ (.A1(\design_top.core0.REG1[8][31] ),
    .A2(_08393_),
    .B1(_08324_),
    .B2(_08396_),
    .X(_04164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11735_ (.A1(\design_top.core0.REG1[8][30] ),
    .A2(_08393_),
    .B1(_08328_),
    .B2(_08396_),
    .X(_04163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11736_ (.A1(\design_top.core0.REG1[8][29] ),
    .A2(_08393_),
    .B1(_08329_),
    .B2(_08396_),
    .X(_04162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11737_ (.A1(\design_top.core0.REG1[8][28] ),
    .A2(_08393_),
    .B1(_08330_),
    .B2(_08396_),
    .X(_04161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11738_ (.A(_08392_),
    .X(_08397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11739_ (.A1(\design_top.core0.REG1[8][27] ),
    .A2(_08397_),
    .B1(_08332_),
    .B2(_08396_),
    .X(_04160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11740_ (.A(_08395_),
    .X(_08398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11741_ (.A1(\design_top.core0.REG1[8][26] ),
    .A2(_08397_),
    .B1(_08333_),
    .B2(_08398_),
    .X(_04159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11742_ (.A1(\design_top.core0.REG1[8][25] ),
    .A2(_08397_),
    .B1(_08335_),
    .B2(_08398_),
    .X(_04158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11743_ (.A1(\design_top.core0.REG1[8][24] ),
    .A2(_08397_),
    .B1(_08336_),
    .B2(_08398_),
    .X(_04157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11744_ (.A1(\design_top.core0.REG1[8][23] ),
    .A2(_08397_),
    .B1(_08337_),
    .B2(_08398_),
    .X(_04156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11745_ (.A(_08392_),
    .X(_08399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11746_ (.A1(\design_top.core0.REG1[8][22] ),
    .A2(_08399_),
    .B1(_08339_),
    .B2(_08398_),
    .X(_04155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11747_ (.A(_08395_),
    .X(_08400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11748_ (.A1(\design_top.core0.REG1[8][21] ),
    .A2(_08399_),
    .B1(_08340_),
    .B2(_08400_),
    .X(_04154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11749_ (.A1(\design_top.core0.REG1[8][20] ),
    .A2(_08399_),
    .B1(_08342_),
    .B2(_08400_),
    .X(_04153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11750_ (.A1(\design_top.core0.REG1[8][19] ),
    .A2(_08399_),
    .B1(_08343_),
    .B2(_08400_),
    .X(_04152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11751_ (.A1(\design_top.core0.REG1[8][18] ),
    .A2(_08399_),
    .B1(_08344_),
    .B2(_08400_),
    .X(_04151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11752_ (.A(_08391_),
    .X(_08401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11753_ (.A1(\design_top.core0.REG1[8][17] ),
    .A2(_08401_),
    .B1(_08346_),
    .B2(_08400_),
    .X(_04150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11754_ (.A(_08394_),
    .X(_08402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11755_ (.A1(\design_top.core0.REG1[8][16] ),
    .A2(_08401_),
    .B1(_08347_),
    .B2(_08402_),
    .X(_04149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11756_ (.A1(\design_top.core0.REG1[8][15] ),
    .A2(_08401_),
    .B1(_08349_),
    .B2(_08402_),
    .X(_04148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11757_ (.A1(\design_top.core0.REG1[8][14] ),
    .A2(_08401_),
    .B1(_08350_),
    .B2(_08402_),
    .X(_04147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11758_ (.A1(\design_top.core0.REG1[8][13] ),
    .A2(_08395_),
    .B1(_08297_),
    .B2(_08393_),
    .X(_04146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11759_ (.A1(\design_top.core0.REG1[8][12] ),
    .A2(_08401_),
    .B1(_08351_),
    .B2(_08402_),
    .X(_04145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11760_ (.A(_08391_),
    .X(_08403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11761_ (.A1(\design_top.core0.REG1[8][11] ),
    .A2(_08403_),
    .B1(_08353_),
    .B2(_08402_),
    .X(_04144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11762_ (.A(_08394_),
    .X(_08404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11763_ (.A1(\design_top.core0.REG1[8][10] ),
    .A2(_08403_),
    .B1(_08354_),
    .B2(_08404_),
    .X(_04143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11764_ (.A1(\design_top.core0.REG1[8][9] ),
    .A2(_08403_),
    .B1(_08356_),
    .B2(_08404_),
    .X(_04142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11765_ (.A1(\design_top.core0.REG1[8][8] ),
    .A2(_08403_),
    .B1(_08357_),
    .B2(_08404_),
    .X(_04141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11766_ (.A1(\design_top.core0.REG1[8][7] ),
    .A2(_08403_),
    .B1(_08358_),
    .B2(_08404_),
    .X(_04140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11767_ (.A(_08391_),
    .X(_08405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11768_ (.A1(\design_top.core0.REG1[8][6] ),
    .A2(_08405_),
    .B1(_08360_),
    .B2(_08404_),
    .X(_04139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11769_ (.A(_08394_),
    .X(_08406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11770_ (.A1(\design_top.core0.REG1[8][5] ),
    .A2(_08405_),
    .B1(_08361_),
    .B2(_08406_),
    .X(_04138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11771_ (.A1(\design_top.core0.REG1[8][4] ),
    .A2(_08405_),
    .B1(_08363_),
    .B2(_08406_),
    .X(_04137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11772_ (.A1(\design_top.core0.REG1[8][3] ),
    .A2(_08405_),
    .B1(_08364_),
    .B2(_08406_),
    .X(_04136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11773_ (.A1(\design_top.core0.REG1[8][2] ),
    .A2(_08405_),
    .B1(_08365_),
    .B2(_08406_),
    .X(_04135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11774_ (.A1(\design_top.core0.REG1[8][1] ),
    .A2(_08392_),
    .B1(_08366_),
    .B2(_08406_),
    .X(_04134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11775_ (.A1(\design_top.core0.REG1[8][0] ),
    .A2(_08392_),
    .B1(_08367_),
    .B2(_08395_),
    .X(_04133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11776_ (.A(\design_top.core0.REG1[0][31] ),
    .Y(_00823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11777_ (.A(_08075_),
    .X(_08407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11778_ (.A(_08407_),
    .B(_08166_),
    .X(_08408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11779_ (.A(_08408_),
    .Y(_08409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11780_ (.A(_00823_),
    .B(_08409_),
    .Y(_04132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11781_ (.A(_08408_),
    .X(_08410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11782_ (.A(_08410_),
    .X(_08411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11783_ (.A(\design_top.core0.REG1[0][30] ),
    .B(_08411_),
    .X(_04131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11784_ (.A(\design_top.core0.REG1[0][29] ),
    .B(_08411_),
    .X(_04130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11785_ (.A(\design_top.core0.REG1[0][28] ),
    .B(_08411_),
    .X(_04129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11786_ (.A(\design_top.core0.REG1[0][27] ),
    .B(_08411_),
    .X(_04128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11787_ (.A(_08410_),
    .X(_08412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11788_ (.A(\design_top.core0.REG1[0][26] ),
    .B(_08412_),
    .X(_04127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11789_ (.A(\design_top.core0.REG1[0][25] ),
    .B(_08412_),
    .X(_04126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11790_ (.A(\design_top.core0.REG1[0][24] ),
    .B(_08412_),
    .X(_04125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11791_ (.A(\design_top.core0.REG1[0][23] ),
    .B(_08412_),
    .X(_04124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11792_ (.A(\design_top.core0.REG1[0][22] ),
    .B(_08412_),
    .X(_04123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11793_ (.A(_08410_),
    .X(_08413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11794_ (.A(\design_top.core0.REG1[0][21] ),
    .B(_08413_),
    .X(_04122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11795_ (.A(\design_top.core0.REG1[0][20] ),
    .B(_08413_),
    .X(_04121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11796_ (.A(\design_top.core0.REG1[0][19] ),
    .B(_08413_),
    .X(_04120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11797_ (.A(\design_top.core0.REG1[0][18] ),
    .B(_08413_),
    .X(_04119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11798_ (.A(\design_top.core0.REG1[0][17] ),
    .Y(_01028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _11799_ (.A(_01028_),
    .B(_08409_),
    .Y(_04118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11800_ (.A(\design_top.core0.REG1[0][16] ),
    .B(_08413_),
    .X(_04117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11801_ (.A(_08410_),
    .X(_08414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11802_ (.A(\design_top.core0.REG1[0][15] ),
    .B(_08414_),
    .X(_04116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11803_ (.A(\design_top.core0.REG1[0][14] ),
    .B(_08414_),
    .X(_04115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11804_ (.A(_00045_),
    .X(_08415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11805_ (.A1(\design_top.core0.REG1[0][13] ),
    .A2(_08409_),
    .B1(_08415_),
    .B2(_08411_),
    .X(_04114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11806_ (.A(\design_top.core0.REG1[0][12] ),
    .B(_08414_),
    .X(_04113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11807_ (.A(\design_top.core0.REG1[0][11] ),
    .B(_08414_),
    .X(_04112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11808_ (.A(\design_top.core0.REG1[0][10] ),
    .B(_08414_),
    .X(_04111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11809_ (.A(_08410_),
    .X(_08416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11810_ (.A(\design_top.core0.REG1[0][9] ),
    .B(_08416_),
    .X(_04110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11811_ (.A(\design_top.core0.REG1[0][8] ),
    .B(_08416_),
    .X(_04109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11812_ (.A(\design_top.core0.REG1[0][7] ),
    .B(_08416_),
    .X(_04108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11813_ (.A(\design_top.core0.REG1[0][6] ),
    .B(_08416_),
    .X(_04107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11814_ (.A(\design_top.core0.REG1[0][5] ),
    .B(_08416_),
    .X(_04106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11815_ (.A(_08408_),
    .X(_08417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11816_ (.A(\design_top.core0.REG1[0][4] ),
    .B(_08417_),
    .X(_04105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11817_ (.A(\design_top.core0.REG1[0][3] ),
    .B(_08417_),
    .X(_04104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11818_ (.A(\design_top.core0.REG1[0][2] ),
    .B(_08417_),
    .X(_04103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11819_ (.A(\design_top.core0.REG1[0][1] ),
    .B(_08417_),
    .X(_04102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _11820_ (.A(\design_top.core0.REG1[0][0] ),
    .B(_08417_),
    .X(_04101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11821_ (.A(_08065_),
    .B(_08249_),
    .C(_08068_),
    .D(_08168_),
    .X(_08418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11822_ (.A(_08302_),
    .B(_08418_),
    .X(_08419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11823_ (.A(_08419_),
    .X(_08420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11824_ (.A(_08420_),
    .X(_08421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11825_ (.A(_08419_),
    .Y(_08422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11826_ (.A(_08422_),
    .X(_08423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11827_ (.A(_08423_),
    .X(_08424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11828_ (.A1(\design_top.core0.REG1[10][31] ),
    .A2(_08421_),
    .B1(_08324_),
    .B2(_08424_),
    .X(_04100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11829_ (.A1(\design_top.core0.REG1[10][30] ),
    .A2(_08421_),
    .B1(_08328_),
    .B2(_08424_),
    .X(_04099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11830_ (.A1(\design_top.core0.REG1[10][29] ),
    .A2(_08421_),
    .B1(_08329_),
    .B2(_08424_),
    .X(_04098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11831_ (.A1(\design_top.core0.REG1[10][28] ),
    .A2(_08421_),
    .B1(_08330_),
    .B2(_08424_),
    .X(_04097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11832_ (.A(_08420_),
    .X(_08425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11833_ (.A1(\design_top.core0.REG1[10][27] ),
    .A2(_08425_),
    .B1(_08332_),
    .B2(_08424_),
    .X(_04096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11834_ (.A(_08423_),
    .X(_08426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11835_ (.A1(\design_top.core0.REG1[10][26] ),
    .A2(_08425_),
    .B1(_08333_),
    .B2(_08426_),
    .X(_04095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11836_ (.A1(\design_top.core0.REG1[10][25] ),
    .A2(_08425_),
    .B1(_08335_),
    .B2(_08426_),
    .X(_04094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11837_ (.A1(\design_top.core0.REG1[10][24] ),
    .A2(_08425_),
    .B1(_08336_),
    .B2(_08426_),
    .X(_04093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11838_ (.A1(\design_top.core0.REG1[10][23] ),
    .A2(_08425_),
    .B1(_08337_),
    .B2(_08426_),
    .X(_04092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11839_ (.A(_08420_),
    .X(_08427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11840_ (.A1(\design_top.core0.REG1[10][22] ),
    .A2(_08427_),
    .B1(_08339_),
    .B2(_08426_),
    .X(_04091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11841_ (.A(_08423_),
    .X(_08428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11842_ (.A1(\design_top.core0.REG1[10][21] ),
    .A2(_08427_),
    .B1(_08340_),
    .B2(_08428_),
    .X(_04090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11843_ (.A1(\design_top.core0.REG1[10][20] ),
    .A2(_08427_),
    .B1(_08342_),
    .B2(_08428_),
    .X(_04089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11844_ (.A1(\design_top.core0.REG1[10][19] ),
    .A2(_08427_),
    .B1(_08343_),
    .B2(_08428_),
    .X(_04088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11845_ (.A1(\design_top.core0.REG1[10][18] ),
    .A2(_08427_),
    .B1(_08344_),
    .B2(_08428_),
    .X(_04087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11846_ (.A(_08419_),
    .X(_08429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11847_ (.A1(\design_top.core0.REG1[10][17] ),
    .A2(_08429_),
    .B1(_08346_),
    .B2(_08428_),
    .X(_04086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11848_ (.A(_08422_),
    .X(_08430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11849_ (.A1(\design_top.core0.REG1[10][16] ),
    .A2(_08429_),
    .B1(_08347_),
    .B2(_08430_),
    .X(_04085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11850_ (.A1(\design_top.core0.REG1[10][15] ),
    .A2(_08429_),
    .B1(_08349_),
    .B2(_08430_),
    .X(_04084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11851_ (.A1(\design_top.core0.REG1[10][14] ),
    .A2(_08429_),
    .B1(_08350_),
    .B2(_08430_),
    .X(_04083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11852_ (.A1(\design_top.core0.REG1[10][13] ),
    .A2(_08423_),
    .B1(_08415_),
    .B2(_08421_),
    .X(_04082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11853_ (.A1(\design_top.core0.REG1[10][12] ),
    .A2(_08429_),
    .B1(_08351_),
    .B2(_08430_),
    .X(_04081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11854_ (.A(_08419_),
    .X(_08431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11855_ (.A1(\design_top.core0.REG1[10][11] ),
    .A2(_08431_),
    .B1(_08353_),
    .B2(_08430_),
    .X(_04080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11856_ (.A(_08422_),
    .X(_08432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11857_ (.A1(\design_top.core0.REG1[10][10] ),
    .A2(_08431_),
    .B1(_08354_),
    .B2(_08432_),
    .X(_04079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11858_ (.A1(\design_top.core0.REG1[10][9] ),
    .A2(_08431_),
    .B1(_08356_),
    .B2(_08432_),
    .X(_04078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11859_ (.A1(\design_top.core0.REG1[10][8] ),
    .A2(_08431_),
    .B1(_08357_),
    .B2(_08432_),
    .X(_04077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11860_ (.A1(\design_top.core0.REG1[10][7] ),
    .A2(_08431_),
    .B1(_08358_),
    .B2(_08432_),
    .X(_04076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11861_ (.A(_08419_),
    .X(_08433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11862_ (.A1(\design_top.core0.REG1[10][6] ),
    .A2(_08433_),
    .B1(_08360_),
    .B2(_08432_),
    .X(_04075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11863_ (.A(_08422_),
    .X(_08434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11864_ (.A1(\design_top.core0.REG1[10][5] ),
    .A2(_08433_),
    .B1(_08361_),
    .B2(_08434_),
    .X(_04074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11865_ (.A1(\design_top.core0.REG1[10][4] ),
    .A2(_08433_),
    .B1(_08363_),
    .B2(_08434_),
    .X(_04073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11866_ (.A1(\design_top.core0.REG1[10][3] ),
    .A2(_08433_),
    .B1(_08364_),
    .B2(_08434_),
    .X(_04072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11867_ (.A1(\design_top.core0.REG1[10][2] ),
    .A2(_08433_),
    .B1(_08365_),
    .B2(_08434_),
    .X(_04071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11868_ (.A1(\design_top.core0.REG1[10][1] ),
    .A2(_08420_),
    .B1(_08366_),
    .B2(_08434_),
    .X(_04070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11869_ (.A1(\design_top.core0.REG1[10][0] ),
    .A2(_08420_),
    .B1(_08367_),
    .B2(_08423_),
    .X(_04069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11870_ (.A(_08078_),
    .X(_08435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11871_ (.A(_08064_),
    .B(_08067_),
    .C(_08068_),
    .D(_01601_),
    .X(_08436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11872_ (.A(_08435_),
    .B(_08436_),
    .X(_08437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11873_ (.A(_08437_),
    .X(_08438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11874_ (.A(_08438_),
    .X(_08439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11875_ (.A(_08437_),
    .Y(_08440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11876_ (.A(_08440_),
    .X(_08441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11877_ (.A(_08441_),
    .X(_08442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11878_ (.A1(\design_top.core0.REG1[11][31] ),
    .A2(_08439_),
    .B1(_08324_),
    .B2(_08442_),
    .X(_04068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11879_ (.A1(\design_top.core0.REG1[11][30] ),
    .A2(_08439_),
    .B1(_08328_),
    .B2(_08442_),
    .X(_04067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11880_ (.A1(\design_top.core0.REG1[11][29] ),
    .A2(_08439_),
    .B1(_08329_),
    .B2(_08442_),
    .X(_04066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11881_ (.A1(\design_top.core0.REG1[11][28] ),
    .A2(_08439_),
    .B1(_08330_),
    .B2(_08442_),
    .X(_04065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11882_ (.A(_08438_),
    .X(_08443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11883_ (.A1(\design_top.core0.REG1[11][27] ),
    .A2(_08443_),
    .B1(_08332_),
    .B2(_08442_),
    .X(_04064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11884_ (.A(_08441_),
    .X(_08444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11885_ (.A1(\design_top.core0.REG1[11][26] ),
    .A2(_08443_),
    .B1(_08333_),
    .B2(_08444_),
    .X(_04063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11886_ (.A1(\design_top.core0.REG1[11][25] ),
    .A2(_08443_),
    .B1(_08335_),
    .B2(_08444_),
    .X(_04062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11887_ (.A1(\design_top.core0.REG1[11][24] ),
    .A2(_08443_),
    .B1(_08336_),
    .B2(_08444_),
    .X(_04061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11888_ (.A1(\design_top.core0.REG1[11][23] ),
    .A2(_08443_),
    .B1(_08337_),
    .B2(_08444_),
    .X(_04060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11889_ (.A(_08438_),
    .X(_08445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11890_ (.A1(\design_top.core0.REG1[11][22] ),
    .A2(_08445_),
    .B1(_08339_),
    .B2(_08444_),
    .X(_04059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11891_ (.A(_08441_),
    .X(_08446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11892_ (.A1(\design_top.core0.REG1[11][21] ),
    .A2(_08445_),
    .B1(_08340_),
    .B2(_08446_),
    .X(_04058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11893_ (.A1(\design_top.core0.REG1[11][20] ),
    .A2(_08445_),
    .B1(_08342_),
    .B2(_08446_),
    .X(_04057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11894_ (.A1(\design_top.core0.REG1[11][19] ),
    .A2(_08445_),
    .B1(_08343_),
    .B2(_08446_),
    .X(_04056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11895_ (.A1(\design_top.core0.REG1[11][18] ),
    .A2(_08445_),
    .B1(_08344_),
    .B2(_08446_),
    .X(_04055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11896_ (.A(_08437_),
    .X(_08447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11897_ (.A1(\design_top.core0.REG1[11][17] ),
    .A2(_08447_),
    .B1(_08346_),
    .B2(_08446_),
    .X(_04054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11898_ (.A(_08440_),
    .X(_08448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11899_ (.A1(\design_top.core0.REG1[11][16] ),
    .A2(_08447_),
    .B1(_08347_),
    .B2(_08448_),
    .X(_04053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11900_ (.A1(\design_top.core0.REG1[11][15] ),
    .A2(_08447_),
    .B1(_08349_),
    .B2(_08448_),
    .X(_04052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11901_ (.A1(\design_top.core0.REG1[11][14] ),
    .A2(_08447_),
    .B1(_08350_),
    .B2(_08448_),
    .X(_04051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11902_ (.A1(\design_top.core0.REG1[11][13] ),
    .A2(_08441_),
    .B1(_08415_),
    .B2(_08439_),
    .X(_04050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11903_ (.A1(\design_top.core0.REG1[11][12] ),
    .A2(_08447_),
    .B1(_08351_),
    .B2(_08448_),
    .X(_04049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11904_ (.A(_08437_),
    .X(_08449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11905_ (.A1(\design_top.core0.REG1[11][11] ),
    .A2(_08449_),
    .B1(_08353_),
    .B2(_08448_),
    .X(_04048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11906_ (.A(_08440_),
    .X(_08450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11907_ (.A1(\design_top.core0.REG1[11][10] ),
    .A2(_08449_),
    .B1(_08354_),
    .B2(_08450_),
    .X(_04047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11908_ (.A1(\design_top.core0.REG1[11][9] ),
    .A2(_08449_),
    .B1(_08356_),
    .B2(_08450_),
    .X(_04046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11909_ (.A1(\design_top.core0.REG1[11][8] ),
    .A2(_08449_),
    .B1(_08357_),
    .B2(_08450_),
    .X(_04045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11910_ (.A1(\design_top.core0.REG1[11][7] ),
    .A2(_08449_),
    .B1(_08358_),
    .B2(_08450_),
    .X(_04044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11911_ (.A(_08437_),
    .X(_08451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11912_ (.A1(\design_top.core0.REG1[11][6] ),
    .A2(_08451_),
    .B1(_08360_),
    .B2(_08450_),
    .X(_04043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11913_ (.A(_08440_),
    .X(_08452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11914_ (.A1(\design_top.core0.REG1[11][5] ),
    .A2(_08451_),
    .B1(_08361_),
    .B2(_08452_),
    .X(_04042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11915_ (.A1(\design_top.core0.REG1[11][4] ),
    .A2(_08451_),
    .B1(_08363_),
    .B2(_08452_),
    .X(_04041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11916_ (.A1(\design_top.core0.REG1[11][3] ),
    .A2(_08451_),
    .B1(_08364_),
    .B2(_08452_),
    .X(_04040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11917_ (.A1(\design_top.core0.REG1[11][2] ),
    .A2(_08451_),
    .B1(_08365_),
    .B2(_08452_),
    .X(_04039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11918_ (.A1(\design_top.core0.REG1[11][1] ),
    .A2(_08438_),
    .B1(_08366_),
    .B2(_08452_),
    .X(_04038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11919_ (.A1(\design_top.core0.REG1[11][0] ),
    .A2(_08438_),
    .B1(_08367_),
    .B2(_08441_),
    .X(_04037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _11920_ (.A(_08069_),
    .B(_08071_),
    .C(_01600_),
    .D(_01599_),
    .X(_08453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _11921_ (.A(_08435_),
    .B(_08453_),
    .X(_08454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11922_ (.A(_08454_),
    .X(_08455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11923_ (.A(_08455_),
    .X(_08456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11924_ (.A(_08174_),
    .X(_08457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _11925_ (.A(_08454_),
    .Y(_08458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11926_ (.A(_08458_),
    .X(_08459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11927_ (.A(_08459_),
    .X(_08460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11928_ (.A1(\design_top.core0.REG1[12][31] ),
    .A2(_08456_),
    .B1(_08457_),
    .B2(_08460_),
    .X(_04036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11929_ (.A(_08179_),
    .X(_08461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11930_ (.A1(\design_top.core0.REG1[12][30] ),
    .A2(_08456_),
    .B1(_08461_),
    .B2(_08460_),
    .X(_04035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11931_ (.A(_08181_),
    .X(_08462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11932_ (.A1(\design_top.core0.REG1[12][29] ),
    .A2(_08456_),
    .B1(_08462_),
    .B2(_08460_),
    .X(_04034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11933_ (.A(_08183_),
    .X(_08463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11934_ (.A1(\design_top.core0.REG1[12][28] ),
    .A2(_08456_),
    .B1(_08463_),
    .B2(_08460_),
    .X(_04033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11935_ (.A(_08455_),
    .X(_08464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11936_ (.A(_08186_),
    .X(_08465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11937_ (.A1(\design_top.core0.REG1[12][27] ),
    .A2(_08464_),
    .B1(_08465_),
    .B2(_08460_),
    .X(_04032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11938_ (.A(_08188_),
    .X(_08466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11939_ (.A(_08459_),
    .X(_08467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11940_ (.A1(\design_top.core0.REG1[12][26] ),
    .A2(_08464_),
    .B1(_08466_),
    .B2(_08467_),
    .X(_04031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11941_ (.A(_08191_),
    .X(_08468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11942_ (.A1(\design_top.core0.REG1[12][25] ),
    .A2(_08464_),
    .B1(_08468_),
    .B2(_08467_),
    .X(_04030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11943_ (.A(_08193_),
    .X(_08469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11944_ (.A1(\design_top.core0.REG1[12][24] ),
    .A2(_08464_),
    .B1(_08469_),
    .B2(_08467_),
    .X(_04029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11945_ (.A(_08195_),
    .X(_08470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11946_ (.A1(\design_top.core0.REG1[12][23] ),
    .A2(_08464_),
    .B1(_08470_),
    .B2(_08467_),
    .X(_04028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11947_ (.A(_08455_),
    .X(_08471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11948_ (.A(_08198_),
    .X(_08472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11949_ (.A1(\design_top.core0.REG1[12][22] ),
    .A2(_08471_),
    .B1(_08472_),
    .B2(_08467_),
    .X(_04027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11950_ (.A(_08200_),
    .X(_08473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11951_ (.A(_08459_),
    .X(_08474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11952_ (.A1(\design_top.core0.REG1[12][21] ),
    .A2(_08471_),
    .B1(_08473_),
    .B2(_08474_),
    .X(_04026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11953_ (.A(_08203_),
    .X(_08475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11954_ (.A1(\design_top.core0.REG1[12][20] ),
    .A2(_08471_),
    .B1(_08475_),
    .B2(_08474_),
    .X(_04025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11955_ (.A(_08205_),
    .X(_08476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11956_ (.A1(\design_top.core0.REG1[12][19] ),
    .A2(_08471_),
    .B1(_08476_),
    .B2(_08474_),
    .X(_04024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11957_ (.A(_08207_),
    .X(_08477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11958_ (.A1(\design_top.core0.REG1[12][18] ),
    .A2(_08471_),
    .B1(_08477_),
    .B2(_08474_),
    .X(_04023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11959_ (.A(_08454_),
    .X(_08478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11960_ (.A(_08210_),
    .X(_08479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11961_ (.A1(\design_top.core0.REG1[12][17] ),
    .A2(_08478_),
    .B1(_08479_),
    .B2(_08474_),
    .X(_04022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11962_ (.A(_08212_),
    .X(_08480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11963_ (.A(_08458_),
    .X(_08481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11964_ (.A1(\design_top.core0.REG1[12][16] ),
    .A2(_08478_),
    .B1(_08480_),
    .B2(_08481_),
    .X(_04021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11965_ (.A(_08215_),
    .X(_08482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11966_ (.A1(\design_top.core0.REG1[12][15] ),
    .A2(_08478_),
    .B1(_08482_),
    .B2(_08481_),
    .X(_04020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11967_ (.A(_08217_),
    .X(_08483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11968_ (.A1(\design_top.core0.REG1[12][14] ),
    .A2(_08478_),
    .B1(_08483_),
    .B2(_08481_),
    .X(_04019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _11969_ (.A1(\design_top.core0.REG1[12][13] ),
    .A2(_08459_),
    .B1(_08415_),
    .B2(_08456_),
    .X(_04018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11970_ (.A(_08219_),
    .X(_08484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11971_ (.A1(\design_top.core0.REG1[12][12] ),
    .A2(_08478_),
    .B1(_08484_),
    .B2(_08481_),
    .X(_04017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11972_ (.A(_08454_),
    .X(_08485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11973_ (.A(_08222_),
    .X(_08486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11974_ (.A1(\design_top.core0.REG1[12][11] ),
    .A2(_08485_),
    .B1(_08486_),
    .B2(_08481_),
    .X(_04016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11975_ (.A(_08224_),
    .X(_08487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11976_ (.A(_08458_),
    .X(_08488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11977_ (.A1(\design_top.core0.REG1[12][10] ),
    .A2(_08485_),
    .B1(_08487_),
    .B2(_08488_),
    .X(_04015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11978_ (.A(_08227_),
    .X(_08489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11979_ (.A1(\design_top.core0.REG1[12][9] ),
    .A2(_08485_),
    .B1(_08489_),
    .B2(_08488_),
    .X(_04014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11980_ (.A(_08229_),
    .X(_08490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11981_ (.A1(\design_top.core0.REG1[12][8] ),
    .A2(_08485_),
    .B1(_08490_),
    .B2(_08488_),
    .X(_04013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11982_ (.A(_08231_),
    .X(_08491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11983_ (.A1(\design_top.core0.REG1[12][7] ),
    .A2(_08485_),
    .B1(_08491_),
    .B2(_08488_),
    .X(_04012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11984_ (.A(_08454_),
    .X(_08492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11985_ (.A(_08234_),
    .X(_08493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11986_ (.A1(\design_top.core0.REG1[12][6] ),
    .A2(_08492_),
    .B1(_08493_),
    .B2(_08488_),
    .X(_04011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11987_ (.A(_08236_),
    .X(_08494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11988_ (.A(_08458_),
    .X(_08495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11989_ (.A1(\design_top.core0.REG1[12][5] ),
    .A2(_08492_),
    .B1(_08494_),
    .B2(_08495_),
    .X(_04010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11990_ (.A(_08239_),
    .X(_08496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11991_ (.A1(\design_top.core0.REG1[12][4] ),
    .A2(_08492_),
    .B1(_08496_),
    .B2(_08495_),
    .X(_04009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11992_ (.A(_08241_),
    .X(_08497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11993_ (.A1(\design_top.core0.REG1[12][3] ),
    .A2(_08492_),
    .B1(_08497_),
    .B2(_08495_),
    .X(_04008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11994_ (.A(_08243_),
    .X(_08498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11995_ (.A1(\design_top.core0.REG1[12][2] ),
    .A2(_08492_),
    .B1(_08498_),
    .B2(_08495_),
    .X(_04007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11996_ (.A(_08245_),
    .X(_08499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11997_ (.A1(\design_top.core0.REG1[12][1] ),
    .A2(_08455_),
    .B1(_08499_),
    .B2(_08495_),
    .X(_04006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _11998_ (.A(_08247_),
    .X(_08500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _11999_ (.A1(\design_top.core0.REG1[12][0] ),
    .A2(_08455_),
    .B1(_08500_),
    .B2(_08459_),
    .X(_04005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _12000_ (.A(_08069_),
    .B(_08071_),
    .C(_01600_),
    .D(_08066_),
    .X(_08501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12001_ (.A(_08435_),
    .B(_08501_),
    .X(_08502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12002_ (.A(_08502_),
    .X(_08503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12003_ (.A(_08503_),
    .X(_08504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12004_ (.A(_08502_),
    .Y(_08505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12005_ (.A(_08505_),
    .X(_08506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12006_ (.A(_08506_),
    .X(_08507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12007_ (.A1(\design_top.core0.REG1[13][31] ),
    .A2(_08504_),
    .B1(_08457_),
    .B2(_08507_),
    .X(_04004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12008_ (.A1(\design_top.core0.REG1[13][30] ),
    .A2(_08504_),
    .B1(_08461_),
    .B2(_08507_),
    .X(_04003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12009_ (.A1(\design_top.core0.REG1[13][29] ),
    .A2(_08504_),
    .B1(_08462_),
    .B2(_08507_),
    .X(_04002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12010_ (.A1(\design_top.core0.REG1[13][28] ),
    .A2(_08504_),
    .B1(_08463_),
    .B2(_08507_),
    .X(_04001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12011_ (.A(_08503_),
    .X(_08508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12012_ (.A1(\design_top.core0.REG1[13][27] ),
    .A2(_08508_),
    .B1(_08465_),
    .B2(_08507_),
    .X(_04000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12013_ (.A(_08506_),
    .X(_08509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12014_ (.A1(\design_top.core0.REG1[13][26] ),
    .A2(_08508_),
    .B1(_08466_),
    .B2(_08509_),
    .X(_03999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12015_ (.A1(\design_top.core0.REG1[13][25] ),
    .A2(_08508_),
    .B1(_08468_),
    .B2(_08509_),
    .X(_03998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12016_ (.A1(\design_top.core0.REG1[13][24] ),
    .A2(_08508_),
    .B1(_08469_),
    .B2(_08509_),
    .X(_03997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12017_ (.A1(\design_top.core0.REG1[13][23] ),
    .A2(_08508_),
    .B1(_08470_),
    .B2(_08509_),
    .X(_03996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12018_ (.A(_08503_),
    .X(_08510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12019_ (.A1(\design_top.core0.REG1[13][22] ),
    .A2(_08510_),
    .B1(_08472_),
    .B2(_08509_),
    .X(_03995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12020_ (.A(_08506_),
    .X(_08511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12021_ (.A1(\design_top.core0.REG1[13][21] ),
    .A2(_08510_),
    .B1(_08473_),
    .B2(_08511_),
    .X(_03994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12022_ (.A1(\design_top.core0.REG1[13][20] ),
    .A2(_08510_),
    .B1(_08475_),
    .B2(_08511_),
    .X(_03993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12023_ (.A1(\design_top.core0.REG1[13][19] ),
    .A2(_08510_),
    .B1(_08476_),
    .B2(_08511_),
    .X(_03992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12024_ (.A1(\design_top.core0.REG1[13][18] ),
    .A2(_08510_),
    .B1(_08477_),
    .B2(_08511_),
    .X(_03991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12025_ (.A(_08502_),
    .X(_08512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12026_ (.A1(\design_top.core0.REG1[13][17] ),
    .A2(_08512_),
    .B1(_08479_),
    .B2(_08511_),
    .X(_03990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12027_ (.A(_08505_),
    .X(_08513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12028_ (.A1(\design_top.core0.REG1[13][16] ),
    .A2(_08512_),
    .B1(_08480_),
    .B2(_08513_),
    .X(_03989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12029_ (.A1(\design_top.core0.REG1[13][15] ),
    .A2(_08512_),
    .B1(_08482_),
    .B2(_08513_),
    .X(_03988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12030_ (.A1(\design_top.core0.REG1[13][14] ),
    .A2(_08512_),
    .B1(_08483_),
    .B2(_08513_),
    .X(_03987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12031_ (.A1(\design_top.core0.REG1[13][13] ),
    .A2(_08506_),
    .B1(_08415_),
    .B2(_08504_),
    .X(_03986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12032_ (.A1(\design_top.core0.REG1[13][12] ),
    .A2(_08512_),
    .B1(_08484_),
    .B2(_08513_),
    .X(_03985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12033_ (.A(_08502_),
    .X(_08514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12034_ (.A1(\design_top.core0.REG1[13][11] ),
    .A2(_08514_),
    .B1(_08486_),
    .B2(_08513_),
    .X(_03984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12035_ (.A(_08505_),
    .X(_08515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12036_ (.A1(\design_top.core0.REG1[13][10] ),
    .A2(_08514_),
    .B1(_08487_),
    .B2(_08515_),
    .X(_03983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12037_ (.A1(\design_top.core0.REG1[13][9] ),
    .A2(_08514_),
    .B1(_08489_),
    .B2(_08515_),
    .X(_03982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12038_ (.A1(\design_top.core0.REG1[13][8] ),
    .A2(_08514_),
    .B1(_08490_),
    .B2(_08515_),
    .X(_03981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12039_ (.A1(\design_top.core0.REG1[13][7] ),
    .A2(_08514_),
    .B1(_08491_),
    .B2(_08515_),
    .X(_03980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12040_ (.A(_08502_),
    .X(_08516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12041_ (.A1(\design_top.core0.REG1[13][6] ),
    .A2(_08516_),
    .B1(_08493_),
    .B2(_08515_),
    .X(_03979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12042_ (.A(_08505_),
    .X(_08517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12043_ (.A1(\design_top.core0.REG1[13][5] ),
    .A2(_08516_),
    .B1(_08494_),
    .B2(_08517_),
    .X(_03978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12044_ (.A1(\design_top.core0.REG1[13][4] ),
    .A2(_08516_),
    .B1(_08496_),
    .B2(_08517_),
    .X(_03977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12045_ (.A1(\design_top.core0.REG1[13][3] ),
    .A2(_08516_),
    .B1(_08497_),
    .B2(_08517_),
    .X(_03976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12046_ (.A1(\design_top.core0.REG1[13][2] ),
    .A2(_08516_),
    .B1(_08498_),
    .B2(_08517_),
    .X(_03975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12047_ (.A1(\design_top.core0.REG1[13][1] ),
    .A2(_08503_),
    .B1(_08499_),
    .B2(_08517_),
    .X(_03974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12048_ (.A1(\design_top.core0.REG1[13][0] ),
    .A2(_08503_),
    .B1(_08500_),
    .B2(_08506_),
    .X(_03973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _12049_ (.A(_08069_),
    .B(_08071_),
    .C(_08064_),
    .D(_01599_),
    .X(_08518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12050_ (.A(_08435_),
    .B(_08518_),
    .X(_08519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12051_ (.A(_08519_),
    .X(_08520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12052_ (.A(_08520_),
    .X(_08521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12053_ (.A(_08519_),
    .Y(_08522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12054_ (.A(_08522_),
    .X(_08523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12055_ (.A(_08523_),
    .X(_08524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12056_ (.A1(\design_top.core0.REG1[14][31] ),
    .A2(_08521_),
    .B1(_08457_),
    .B2(_08524_),
    .X(_03972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12057_ (.A1(\design_top.core0.REG1[14][30] ),
    .A2(_08521_),
    .B1(_08461_),
    .B2(_08524_),
    .X(_03971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12058_ (.A1(\design_top.core0.REG1[14][29] ),
    .A2(_08521_),
    .B1(_08462_),
    .B2(_08524_),
    .X(_03970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12059_ (.A1(\design_top.core0.REG1[14][28] ),
    .A2(_08521_),
    .B1(_08463_),
    .B2(_08524_),
    .X(_03969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12060_ (.A(_08520_),
    .X(_08525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12061_ (.A1(\design_top.core0.REG1[14][27] ),
    .A2(_08525_),
    .B1(_08465_),
    .B2(_08524_),
    .X(_03968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12062_ (.A(_08523_),
    .X(_08526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12063_ (.A1(\design_top.core0.REG1[14][26] ),
    .A2(_08525_),
    .B1(_08466_),
    .B2(_08526_),
    .X(_03967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12064_ (.A1(\design_top.core0.REG1[14][25] ),
    .A2(_08525_),
    .B1(_08468_),
    .B2(_08526_),
    .X(_03966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12065_ (.A1(\design_top.core0.REG1[14][24] ),
    .A2(_08525_),
    .B1(_08469_),
    .B2(_08526_),
    .X(_03965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12066_ (.A1(\design_top.core0.REG1[14][23] ),
    .A2(_08525_),
    .B1(_08470_),
    .B2(_08526_),
    .X(_03964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12067_ (.A(_08520_),
    .X(_08527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12068_ (.A1(\design_top.core0.REG1[14][22] ),
    .A2(_08527_),
    .B1(_08472_),
    .B2(_08526_),
    .X(_03963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12069_ (.A(_08523_),
    .X(_08528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12070_ (.A1(\design_top.core0.REG1[14][21] ),
    .A2(_08527_),
    .B1(_08473_),
    .B2(_08528_),
    .X(_03962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12071_ (.A1(\design_top.core0.REG1[14][20] ),
    .A2(_08527_),
    .B1(_08475_),
    .B2(_08528_),
    .X(_03961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12072_ (.A1(\design_top.core0.REG1[14][19] ),
    .A2(_08527_),
    .B1(_08476_),
    .B2(_08528_),
    .X(_03960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12073_ (.A1(\design_top.core0.REG1[14][18] ),
    .A2(_08527_),
    .B1(_08477_),
    .B2(_08528_),
    .X(_03959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12074_ (.A(_08519_),
    .X(_08529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12075_ (.A1(\design_top.core0.REG1[14][17] ),
    .A2(_08529_),
    .B1(_08479_),
    .B2(_08528_),
    .X(_03958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12076_ (.A(_08522_),
    .X(_08530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12077_ (.A1(\design_top.core0.REG1[14][16] ),
    .A2(_08529_),
    .B1(_08480_),
    .B2(_08530_),
    .X(_03957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12078_ (.A1(\design_top.core0.REG1[14][15] ),
    .A2(_08529_),
    .B1(_08482_),
    .B2(_08530_),
    .X(_03956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12079_ (.A1(\design_top.core0.REG1[14][14] ),
    .A2(_08529_),
    .B1(_08483_),
    .B2(_08530_),
    .X(_03955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12080_ (.A(_00045_),
    .X(_08531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12081_ (.A1(\design_top.core0.REG1[14][13] ),
    .A2(_08523_),
    .B1(_08531_),
    .B2(_08521_),
    .X(_03954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12082_ (.A1(\design_top.core0.REG1[14][12] ),
    .A2(_08529_),
    .B1(_08484_),
    .B2(_08530_),
    .X(_03953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12083_ (.A(_08519_),
    .X(_08532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12084_ (.A1(\design_top.core0.REG1[14][11] ),
    .A2(_08532_),
    .B1(_08486_),
    .B2(_08530_),
    .X(_03952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12085_ (.A(_08522_),
    .X(_08533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12086_ (.A1(\design_top.core0.REG1[14][10] ),
    .A2(_08532_),
    .B1(_08487_),
    .B2(_08533_),
    .X(_03951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12087_ (.A1(\design_top.core0.REG1[14][9] ),
    .A2(_08532_),
    .B1(_08489_),
    .B2(_08533_),
    .X(_03950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12088_ (.A1(\design_top.core0.REG1[14][8] ),
    .A2(_08532_),
    .B1(_08490_),
    .B2(_08533_),
    .X(_03949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12089_ (.A1(\design_top.core0.REG1[14][7] ),
    .A2(_08532_),
    .B1(_08491_),
    .B2(_08533_),
    .X(_03948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12090_ (.A(_08519_),
    .X(_08534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12091_ (.A1(\design_top.core0.REG1[14][6] ),
    .A2(_08534_),
    .B1(_08493_),
    .B2(_08533_),
    .X(_03947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12092_ (.A(_08522_),
    .X(_08535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12093_ (.A1(\design_top.core0.REG1[14][5] ),
    .A2(_08534_),
    .B1(_08494_),
    .B2(_08535_),
    .X(_03946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12094_ (.A1(\design_top.core0.REG1[14][4] ),
    .A2(_08534_),
    .B1(_08496_),
    .B2(_08535_),
    .X(_03945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12095_ (.A1(\design_top.core0.REG1[14][3] ),
    .A2(_08534_),
    .B1(_08497_),
    .B2(_08535_),
    .X(_03944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12096_ (.A1(\design_top.core0.REG1[14][2] ),
    .A2(_08534_),
    .B1(_08498_),
    .B2(_08535_),
    .X(_03943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12097_ (.A1(\design_top.core0.REG1[14][1] ),
    .A2(_08520_),
    .B1(_08499_),
    .B2(_08535_),
    .X(_03942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12098_ (.A1(\design_top.core0.REG1[14][0] ),
    .A2(_08520_),
    .B1(_08500_),
    .B2(_08523_),
    .X(_03941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12099_ (.A1(_07189_),
    .A2(_07131_),
    .B1(_07155_),
    .B2(_08385_),
    .X(_08536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12100_ (.A(_08536_),
    .Y(_08537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12101_ (.A(_08537_),
    .X(_08538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12102_ (.A(_08536_),
    .X(_08539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12103_ (.A1(_00396_),
    .A2(_08538_),
    .B1(\design_top.MEM[5][7] ),
    .B2(_08539_),
    .X(_03940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12104_ (.A1(_00395_),
    .A2(_08538_),
    .B1(\design_top.MEM[5][6] ),
    .B2(_08539_),
    .X(_03939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12105_ (.A1(_00394_),
    .A2(_08538_),
    .B1(\design_top.MEM[5][5] ),
    .B2(_08539_),
    .X(_03938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12106_ (.A1(_00393_),
    .A2(_08538_),
    .B1(\design_top.MEM[5][4] ),
    .B2(_08539_),
    .X(_03937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12107_ (.A1(_00392_),
    .A2(_08538_),
    .B1(\design_top.MEM[5][3] ),
    .B2(_08539_),
    .X(_03936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12108_ (.A1(_00391_),
    .A2(_08537_),
    .B1(\design_top.MEM[5][2] ),
    .B2(_08536_),
    .X(_03935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12109_ (.A1(_00390_),
    .A2(_08537_),
    .B1(\design_top.MEM[5][1] ),
    .B2(_08536_),
    .X(_03934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12110_ (.A1(_00389_),
    .A2(_08537_),
    .B1(\design_top.MEM[5][0] ),
    .B2(_08536_),
    .X(_03933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12111_ (.A1(_06977_),
    .A2(_07131_),
    .B1(_07169_),
    .B2(_08385_),
    .X(_08540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12112_ (.A(_08540_),
    .Y(_08541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12113_ (.A(_08541_),
    .X(_08542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12114_ (.A(_08540_),
    .X(_08543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12115_ (.A1(_00404_),
    .A2(_08542_),
    .B1(\design_top.MEM[6][7] ),
    .B2(_08543_),
    .X(_03932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12116_ (.A1(_00403_),
    .A2(_08542_),
    .B1(\design_top.MEM[6][6] ),
    .B2(_08543_),
    .X(_03931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12117_ (.A1(_00402_),
    .A2(_08542_),
    .B1(\design_top.MEM[6][5] ),
    .B2(_08543_),
    .X(_03930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12118_ (.A1(_00401_),
    .A2(_08542_),
    .B1(\design_top.MEM[6][4] ),
    .B2(_08543_),
    .X(_03929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12119_ (.A1(_00400_),
    .A2(_08542_),
    .B1(\design_top.MEM[6][3] ),
    .B2(_08543_),
    .X(_03928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12120_ (.A1(_00399_),
    .A2(_08541_),
    .B1(\design_top.MEM[6][2] ),
    .B2(_08540_),
    .X(_03927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12121_ (.A1(_00398_),
    .A2(_08541_),
    .B1(\design_top.MEM[6][1] ),
    .B2(_08540_),
    .X(_03926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12122_ (.A1(_00397_),
    .A2(_08541_),
    .B1(\design_top.MEM[6][0] ),
    .B2(_08540_),
    .X(_03925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _12123_ (.A(_08169_),
    .B(_08066_),
    .C(_08068_),
    .D(_01601_),
    .X(_08544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _12124_ (.A(_08435_),
    .B(_08544_),
    .X(_08545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12125_ (.A(_08545_),
    .X(_08546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12126_ (.A(_08546_),
    .X(_08547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12127_ (.A(_08545_),
    .Y(_08548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12128_ (.A(_08548_),
    .X(_08549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12129_ (.A(_08549_),
    .X(_08550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12130_ (.A1(\design_top.core0.REG1[9][31] ),
    .A2(_08547_),
    .B1(_08457_),
    .B2(_08550_),
    .X(_03924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12131_ (.A1(\design_top.core0.REG1[9][30] ),
    .A2(_08547_),
    .B1(_08461_),
    .B2(_08550_),
    .X(_03923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12132_ (.A1(\design_top.core0.REG1[9][29] ),
    .A2(_08547_),
    .B1(_08462_),
    .B2(_08550_),
    .X(_03922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12133_ (.A1(\design_top.core0.REG1[9][28] ),
    .A2(_08547_),
    .B1(_08463_),
    .B2(_08550_),
    .X(_03921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12134_ (.A(_08546_),
    .X(_08551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12135_ (.A1(\design_top.core0.REG1[9][27] ),
    .A2(_08551_),
    .B1(_08465_),
    .B2(_08550_),
    .X(_03920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12136_ (.A(_08549_),
    .X(_08552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12137_ (.A1(\design_top.core0.REG1[9][26] ),
    .A2(_08551_),
    .B1(_08466_),
    .B2(_08552_),
    .X(_03919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12138_ (.A1(\design_top.core0.REG1[9][25] ),
    .A2(_08551_),
    .B1(_08468_),
    .B2(_08552_),
    .X(_03918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12139_ (.A1(\design_top.core0.REG1[9][24] ),
    .A2(_08551_),
    .B1(_08469_),
    .B2(_08552_),
    .X(_03917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12140_ (.A1(\design_top.core0.REG1[9][23] ),
    .A2(_08551_),
    .B1(_08470_),
    .B2(_08552_),
    .X(_03916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12141_ (.A(_08546_),
    .X(_08553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12142_ (.A1(\design_top.core0.REG1[9][22] ),
    .A2(_08553_),
    .B1(_08472_),
    .B2(_08552_),
    .X(_03915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12143_ (.A(_08549_),
    .X(_08554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12144_ (.A1(\design_top.core0.REG1[9][21] ),
    .A2(_08553_),
    .B1(_08473_),
    .B2(_08554_),
    .X(_03914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12145_ (.A1(\design_top.core0.REG1[9][20] ),
    .A2(_08553_),
    .B1(_08475_),
    .B2(_08554_),
    .X(_03913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12146_ (.A1(\design_top.core0.REG1[9][19] ),
    .A2(_08553_),
    .B1(_08476_),
    .B2(_08554_),
    .X(_03912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12147_ (.A1(\design_top.core0.REG1[9][18] ),
    .A2(_08553_),
    .B1(_08477_),
    .B2(_08554_),
    .X(_03911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12148_ (.A(_08545_),
    .X(_08555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12149_ (.A1(\design_top.core0.REG1[9][17] ),
    .A2(_08555_),
    .B1(_08479_),
    .B2(_08554_),
    .X(_03910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12150_ (.A(_08548_),
    .X(_08556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12151_ (.A1(\design_top.core0.REG1[9][16] ),
    .A2(_08555_),
    .B1(_08480_),
    .B2(_08556_),
    .X(_03909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12152_ (.A1(\design_top.core0.REG1[9][15] ),
    .A2(_08555_),
    .B1(_08482_),
    .B2(_08556_),
    .X(_03908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12153_ (.A1(\design_top.core0.REG1[9][14] ),
    .A2(_08555_),
    .B1(_08483_),
    .B2(_08556_),
    .X(_03907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12154_ (.A1(\design_top.core0.REG1[9][13] ),
    .A2(_08549_),
    .B1(_08531_),
    .B2(_08547_),
    .X(_03906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12155_ (.A1(\design_top.core0.REG1[9][12] ),
    .A2(_08555_),
    .B1(_08484_),
    .B2(_08556_),
    .X(_03905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12156_ (.A(_08545_),
    .X(_08557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12157_ (.A1(\design_top.core0.REG1[9][11] ),
    .A2(_08557_),
    .B1(_08486_),
    .B2(_08556_),
    .X(_03904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12158_ (.A(_08548_),
    .X(_08558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12159_ (.A1(\design_top.core0.REG1[9][10] ),
    .A2(_08557_),
    .B1(_08487_),
    .B2(_08558_),
    .X(_03903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12160_ (.A1(\design_top.core0.REG1[9][9] ),
    .A2(_08557_),
    .B1(_08489_),
    .B2(_08558_),
    .X(_03902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12161_ (.A1(\design_top.core0.REG1[9][8] ),
    .A2(_08557_),
    .B1(_08490_),
    .B2(_08558_),
    .X(_03901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12162_ (.A1(\design_top.core0.REG1[9][7] ),
    .A2(_08557_),
    .B1(_08491_),
    .B2(_08558_),
    .X(_03900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12163_ (.A(_08545_),
    .X(_08559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12164_ (.A1(\design_top.core0.REG1[9][6] ),
    .A2(_08559_),
    .B1(_08493_),
    .B2(_08558_),
    .X(_03899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12165_ (.A(_08548_),
    .X(_08560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12166_ (.A1(\design_top.core0.REG1[9][5] ),
    .A2(_08559_),
    .B1(_08494_),
    .B2(_08560_),
    .X(_03898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12167_ (.A1(\design_top.core0.REG1[9][4] ),
    .A2(_08559_),
    .B1(_08496_),
    .B2(_08560_),
    .X(_03897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12168_ (.A1(\design_top.core0.REG1[9][3] ),
    .A2(_08559_),
    .B1(_08497_),
    .B2(_08560_),
    .X(_03896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12169_ (.A1(\design_top.core0.REG1[9][2] ),
    .A2(_08559_),
    .B1(_08498_),
    .B2(_08560_),
    .X(_03895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12170_ (.A1(\design_top.core0.REG1[9][1] ),
    .A2(_08546_),
    .B1(_08499_),
    .B2(_08560_),
    .X(_03894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12171_ (.A1(\design_top.core0.REG1[9][0] ),
    .A2(_08546_),
    .B1(_08500_),
    .B2(_08549_),
    .X(_03893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12172_ (.A1(_08021_),
    .A2(_07183_),
    .B1(_07194_),
    .B2(_08385_),
    .X(_05495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12173_ (.A(_05495_),
    .Y(_05496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12174_ (.A(_05496_),
    .X(_05497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12175_ (.A(_05495_),
    .X(_05498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12176_ (.A1(_00220_),
    .A2(_05497_),
    .B1(\design_top.MEM[14][7] ),
    .B2(_05498_),
    .X(_03892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12177_ (.A1(_00219_),
    .A2(_05497_),
    .B1(\design_top.MEM[14][6] ),
    .B2(_05498_),
    .X(_03891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12178_ (.A1(_00218_),
    .A2(_05497_),
    .B1(\design_top.MEM[14][5] ),
    .B2(_05498_),
    .X(_03890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12179_ (.A1(_00217_),
    .A2(_05497_),
    .B1(\design_top.MEM[14][4] ),
    .B2(_05498_),
    .X(_03889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12180_ (.A1(_00216_),
    .A2(_05497_),
    .B1(\design_top.MEM[14][3] ),
    .B2(_05498_),
    .X(_03888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12181_ (.A1(_00215_),
    .A2(_05496_),
    .B1(\design_top.MEM[14][2] ),
    .B2(_05495_),
    .X(_03887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12182_ (.A1(_00214_),
    .A2(_05496_),
    .B1(\design_top.MEM[14][1] ),
    .B2(_05495_),
    .X(_03886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12183_ (.A1(_00213_),
    .A2(_05496_),
    .B1(\design_top.MEM[14][0] ),
    .B2(_05495_),
    .X(_03885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12184_ (.A1(_07048_),
    .A2(_07182_),
    .B1(_07218_),
    .B2(_08385_),
    .X(_05499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12185_ (.A(_05499_),
    .Y(_05500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12186_ (.A(_05500_),
    .X(_05501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12187_ (.A(_05499_),
    .X(_05502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12188_ (.A1(_00228_),
    .A2(_05501_),
    .B1(\design_top.MEM[15][7] ),
    .B2(_05502_),
    .X(_03884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12189_ (.A1(_00227_),
    .A2(_05501_),
    .B1(\design_top.MEM[15][6] ),
    .B2(_05502_),
    .X(_03883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12190_ (.A1(_00226_),
    .A2(_05501_),
    .B1(\design_top.MEM[15][5] ),
    .B2(_05502_),
    .X(_03882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12191_ (.A1(_00225_),
    .A2(_05501_),
    .B1(\design_top.MEM[15][4] ),
    .B2(_05502_),
    .X(_03881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12192_ (.A1(_00224_),
    .A2(_05501_),
    .B1(\design_top.MEM[15][3] ),
    .B2(_05502_),
    .X(_03880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12193_ (.A1(_00223_),
    .A2(_05500_),
    .B1(\design_top.MEM[15][2] ),
    .B2(_05499_),
    .X(_03879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12194_ (.A1(_00222_),
    .A2(_05500_),
    .B1(\design_top.MEM[15][1] ),
    .B2(_05499_),
    .X(_03878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12195_ (.A1(_00221_),
    .A2(_05500_),
    .B1(\design_top.MEM[15][0] ),
    .B2(_05499_),
    .X(_03877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12196_ (.A(_06900_),
    .X(_05503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12197_ (.A(_08022_),
    .X(_05504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12198_ (.A1(_05503_),
    .A2(_07255_),
    .B1(_07251_),
    .B2(_05504_),
    .X(_05505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12199_ (.A(_05505_),
    .Y(_05506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12200_ (.A(_05506_),
    .X(_05507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12201_ (.A(_05505_),
    .X(_05508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12202_ (.A1(_00236_),
    .A2(_05507_),
    .B1(\design_top.MEM[16][7] ),
    .B2(_05508_),
    .X(_03876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12203_ (.A1(_00235_),
    .A2(_05507_),
    .B1(\design_top.MEM[16][6] ),
    .B2(_05508_),
    .X(_03875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12204_ (.A1(_00234_),
    .A2(_05507_),
    .B1(\design_top.MEM[16][5] ),
    .B2(_05508_),
    .X(_03874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12205_ (.A1(_00233_),
    .A2(_05507_),
    .B1(\design_top.MEM[16][4] ),
    .B2(_05508_),
    .X(_03873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12206_ (.A1(_00232_),
    .A2(_05507_),
    .B1(\design_top.MEM[16][3] ),
    .B2(_05508_),
    .X(_03872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12207_ (.A1(_00231_),
    .A2(_05506_),
    .B1(\design_top.MEM[16][2] ),
    .B2(_05505_),
    .X(_03871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12208_ (.A1(_00230_),
    .A2(_05506_),
    .B1(\design_top.MEM[16][1] ),
    .B2(_05505_),
    .X(_03870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12209_ (.A1(_00229_),
    .A2(_05506_),
    .B1(\design_top.MEM[16][0] ),
    .B2(_05505_),
    .X(_03869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12210_ (.A1(_07189_),
    .A2(_07254_),
    .B1(_07267_),
    .B2(_05504_),
    .X(_05509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12211_ (.A(_05509_),
    .Y(_05510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12212_ (.A(_05510_),
    .X(_05511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12213_ (.A(_05509_),
    .X(_05512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12214_ (.A1(_00244_),
    .A2(_05511_),
    .B1(\design_top.MEM[17][7] ),
    .B2(_05512_),
    .X(_03868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12215_ (.A1(_00243_),
    .A2(_05511_),
    .B1(\design_top.MEM[17][6] ),
    .B2(_05512_),
    .X(_03867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12216_ (.A1(_00242_),
    .A2(_05511_),
    .B1(\design_top.MEM[17][5] ),
    .B2(_05512_),
    .X(_03866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12217_ (.A1(_00241_),
    .A2(_05511_),
    .B1(\design_top.MEM[17][4] ),
    .B2(_05512_),
    .X(_03865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12218_ (.A1(_00240_),
    .A2(_05511_),
    .B1(\design_top.MEM[17][3] ),
    .B2(_05512_),
    .X(_03864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12219_ (.A1(_00239_),
    .A2(_05510_),
    .B1(\design_top.MEM[17][2] ),
    .B2(_05509_),
    .X(_03863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12220_ (.A1(_00238_),
    .A2(_05510_),
    .B1(\design_top.MEM[17][1] ),
    .B2(_05509_),
    .X(_03862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12221_ (.A1(_00237_),
    .A2(_05510_),
    .B1(\design_top.MEM[17][0] ),
    .B2(_05509_),
    .X(_03861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12222_ (.A1(_08021_),
    .A2(_07254_),
    .B1(_07281_),
    .B2(_05504_),
    .X(_05513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12223_ (.A(_05513_),
    .Y(_05514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12224_ (.A(_05514_),
    .X(_05515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12225_ (.A(_05513_),
    .X(_05516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12226_ (.A1(_00252_),
    .A2(_05515_),
    .B1(\design_top.MEM[18][7] ),
    .B2(_05516_),
    .X(_03860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12227_ (.A1(_00251_),
    .A2(_05515_),
    .B1(\design_top.MEM[18][6] ),
    .B2(_05516_),
    .X(_03859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12228_ (.A1(_00250_),
    .A2(_05515_),
    .B1(\design_top.MEM[18][5] ),
    .B2(_05516_),
    .X(_03858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12229_ (.A1(_00249_),
    .A2(_05515_),
    .B1(\design_top.MEM[18][4] ),
    .B2(_05516_),
    .X(_03857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12230_ (.A1(_00248_),
    .A2(_05515_),
    .B1(\design_top.MEM[18][3] ),
    .B2(_05516_),
    .X(_03856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12231_ (.A1(_00247_),
    .A2(_05514_),
    .B1(\design_top.MEM[18][2] ),
    .B2(_05513_),
    .X(_03855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12232_ (.A1(_00246_),
    .A2(_05514_),
    .B1(\design_top.MEM[18][1] ),
    .B2(_05513_),
    .X(_03854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12233_ (.A1(_00245_),
    .A2(_05514_),
    .B1(\design_top.MEM[18][0] ),
    .B2(_05513_),
    .X(_03853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12234_ (.A1(_08045_),
    .A2(_07254_),
    .B1(_07296_),
    .B2(_05504_),
    .X(_05517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12235_ (.A(_05517_),
    .Y(_05518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12236_ (.A(_05518_),
    .X(_05519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12237_ (.A(_05517_),
    .X(_05520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12238_ (.A1(_00260_),
    .A2(_05519_),
    .B1(\design_top.MEM[19][7] ),
    .B2(_05520_),
    .X(_03852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12239_ (.A1(_00259_),
    .A2(_05519_),
    .B1(\design_top.MEM[19][6] ),
    .B2(_05520_),
    .X(_03851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12240_ (.A1(_00258_),
    .A2(_05519_),
    .B1(\design_top.MEM[19][5] ),
    .B2(_05520_),
    .X(_03850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12241_ (.A1(_00257_),
    .A2(_05519_),
    .B1(\design_top.MEM[19][4] ),
    .B2(_05520_),
    .X(_03849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12242_ (.A1(_00256_),
    .A2(_05519_),
    .B1(\design_top.MEM[19][3] ),
    .B2(_05520_),
    .X(_03848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12243_ (.A1(_00255_),
    .A2(_05518_),
    .B1(\design_top.MEM[19][2] ),
    .B2(_05517_),
    .X(_03847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12244_ (.A1(_00254_),
    .A2(_05518_),
    .B1(\design_top.MEM[19][1] ),
    .B2(_05517_),
    .X(_03846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12245_ (.A1(_00253_),
    .A2(_05518_),
    .B1(\design_top.MEM[19][0] ),
    .B2(_05517_),
    .X(_03845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12246_ (.A(_06864_),
    .X(_05521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12247_ (.A1(_05521_),
    .A2(_06903_),
    .B1(_07319_),
    .B2(_05504_),
    .X(_05522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12248_ (.A(_05522_),
    .Y(_05523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12249_ (.A(_05523_),
    .X(_05524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12250_ (.A(_05522_),
    .X(_05525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12251_ (.A1(_00268_),
    .A2(_05524_),
    .B1(\design_top.MEM[1][7] ),
    .B2(_05525_),
    .X(_03844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12252_ (.A1(_00267_),
    .A2(_05524_),
    .B1(\design_top.MEM[1][6] ),
    .B2(_05525_),
    .X(_03843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12253_ (.A1(_00266_),
    .A2(_05524_),
    .B1(\design_top.MEM[1][5] ),
    .B2(_05525_),
    .X(_03842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12254_ (.A1(_00265_),
    .A2(_05524_),
    .B1(\design_top.MEM[1][4] ),
    .B2(_05525_),
    .X(_03841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12255_ (.A1(_00264_),
    .A2(_05524_),
    .B1(\design_top.MEM[1][3] ),
    .B2(_05525_),
    .X(_03840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12256_ (.A1(_00263_),
    .A2(_05523_),
    .B1(\design_top.MEM[1][2] ),
    .B2(_05522_),
    .X(_03839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12257_ (.A1(_00262_),
    .A2(_05523_),
    .B1(\design_top.MEM[1][1] ),
    .B2(_05522_),
    .X(_03838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12258_ (.A1(_00261_),
    .A2(_05523_),
    .B1(\design_top.MEM[1][0] ),
    .B2(_05522_),
    .X(_03837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12259_ (.A(_08072_),
    .X(_05526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12260_ (.A(_05526_),
    .X(_05527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12261_ (.A(_05527_),
    .X(_05528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12262_ (.A(_05526_),
    .Y(_05529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12263_ (.A(_05529_),
    .X(_05530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12264_ (.A(_05530_),
    .X(_05531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12265_ (.A1(_05528_),
    .A2(_08089_),
    .B1(\design_top.core0.REG2[15][31] ),
    .B2(_05531_),
    .X(_03836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12266_ (.A1(_05528_),
    .A2(_08091_),
    .B1(\design_top.core0.REG2[15][30] ),
    .B2(_05531_),
    .X(_03835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12267_ (.A1(_05528_),
    .A2(_08093_),
    .B1(\design_top.core0.REG2[15][29] ),
    .B2(_05531_),
    .X(_03834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12268_ (.A1(_05528_),
    .A2(_08095_),
    .B1(\design_top.core0.REG2[15][28] ),
    .B2(_05531_),
    .X(_03833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12269_ (.A1(_05528_),
    .A2(_08098_),
    .B1(\design_top.core0.REG2[15][27] ),
    .B2(_05531_),
    .X(_03832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12270_ (.A(_05527_),
    .X(_05532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12271_ (.A(_05530_),
    .X(_05533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12272_ (.A1(_05532_),
    .A2(_08102_),
    .B1(\design_top.core0.REG2[15][26] ),
    .B2(_05533_),
    .X(_03831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12273_ (.A1(_05532_),
    .A2(_08104_),
    .B1(\design_top.core0.REG2[15][25] ),
    .B2(_05533_),
    .X(_03830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12274_ (.A1(_05532_),
    .A2(_08106_),
    .B1(\design_top.core0.REG2[15][24] ),
    .B2(_05533_),
    .X(_03829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12275_ (.A1(_05532_),
    .A2(_08108_),
    .B1(\design_top.core0.REG2[15][23] ),
    .B2(_05533_),
    .X(_03828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12276_ (.A1(_05532_),
    .A2(_08111_),
    .B1(\design_top.core0.REG2[15][22] ),
    .B2(_05533_),
    .X(_03827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12277_ (.A(_05527_),
    .X(_05534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12278_ (.A(_05530_),
    .X(_05535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12279_ (.A1(_05534_),
    .A2(_08115_),
    .B1(\design_top.core0.REG2[15][21] ),
    .B2(_05535_),
    .X(_03826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12280_ (.A1(_05534_),
    .A2(_08117_),
    .B1(\design_top.core0.REG2[15][20] ),
    .B2(_05535_),
    .X(_03825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12281_ (.A1(_05534_),
    .A2(_08119_),
    .B1(\design_top.core0.REG2[15][19] ),
    .B2(_05535_),
    .X(_03824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12282_ (.A1(_05534_),
    .A2(_08121_),
    .B1(\design_top.core0.REG2[15][18] ),
    .B2(_05535_),
    .X(_03823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12283_ (.A1(_05534_),
    .A2(_08124_),
    .B1(\design_top.core0.REG2[15][17] ),
    .B2(_05535_),
    .X(_03822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12284_ (.A(_05526_),
    .X(_05536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12285_ (.A(_05529_),
    .X(_05537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12286_ (.A1(_05536_),
    .A2(_08128_),
    .B1(\design_top.core0.REG2[15][16] ),
    .B2(_05537_),
    .X(_03821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12287_ (.A1(_05536_),
    .A2(_08130_),
    .B1(\design_top.core0.REG2[15][15] ),
    .B2(_05537_),
    .X(_03820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12288_ (.A1(_05536_),
    .A2(_08132_),
    .B1(\design_top.core0.REG2[15][14] ),
    .B2(_05537_),
    .X(_03819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12289_ (.A(_08531_),
    .X(_05538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12290_ (.A1(\design_top.core0.REG2[15][13] ),
    .A2(_05527_),
    .B1(_05538_),
    .B2(_05530_),
    .X(_03818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12291_ (.A1(_05536_),
    .A2(_08135_),
    .B1(\design_top.core0.REG2[15][12] ),
    .B2(_05537_),
    .X(_03817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12292_ (.A1(_05536_),
    .A2(_08138_),
    .B1(\design_top.core0.REG2[15][11] ),
    .B2(_05537_),
    .X(_03816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12293_ (.A(_05526_),
    .X(_05539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12294_ (.A(_05529_),
    .X(_05540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12295_ (.A1(_05539_),
    .A2(_08142_),
    .B1(\design_top.core0.REG2[15][10] ),
    .B2(_05540_),
    .X(_03815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12296_ (.A1(_05539_),
    .A2(_08144_),
    .B1(\design_top.core0.REG2[15][9] ),
    .B2(_05540_),
    .X(_03814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12297_ (.A1(_05539_),
    .A2(_08146_),
    .B1(\design_top.core0.REG2[15][8] ),
    .B2(_05540_),
    .X(_03813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12298_ (.A1(_05539_),
    .A2(_08148_),
    .B1(\design_top.core0.REG2[15][7] ),
    .B2(_05540_),
    .X(_03812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12299_ (.A1(_05539_),
    .A2(_08151_),
    .B1(\design_top.core0.REG2[15][6] ),
    .B2(_05540_),
    .X(_03811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12300_ (.A(_05526_),
    .X(_05541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12301_ (.A(_05529_),
    .X(_05542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12302_ (.A1(_05541_),
    .A2(_08155_),
    .B1(\design_top.core0.REG2[15][5] ),
    .B2(_05542_),
    .X(_03810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12303_ (.A1(_05541_),
    .A2(_08157_),
    .B1(\design_top.core0.REG2[15][4] ),
    .B2(_05542_),
    .X(_03809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12304_ (.A1(_05541_),
    .A2(_08159_),
    .B1(\design_top.core0.REG2[15][3] ),
    .B2(_05542_),
    .X(_03808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12305_ (.A1(_05541_),
    .A2(_08161_),
    .B1(\design_top.core0.REG2[15][2] ),
    .B2(_05542_),
    .X(_03807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12306_ (.A1(_05541_),
    .A2(_08163_),
    .B1(\design_top.core0.REG2[15][1] ),
    .B2(_05542_),
    .X(_03806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12307_ (.A1(_05527_),
    .A2(_08165_),
    .B1(\design_top.core0.REG2[15][0] ),
    .B2(_05530_),
    .X(_03805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12308_ (.A(_08170_),
    .X(_05543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12309_ (.A(_05543_),
    .X(_05544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12310_ (.A(_05544_),
    .X(_05545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12311_ (.A(_05543_),
    .Y(_05546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12312_ (.A(_05546_),
    .X(_05547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12313_ (.A(_05547_),
    .X(_05548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12314_ (.A1(_08457_),
    .A2(_05545_),
    .B1(\design_top.core0.REG2[1][31] ),
    .B2(_05548_),
    .X(_03804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12315_ (.A1(_08461_),
    .A2(_05545_),
    .B1(\design_top.core0.REG2[1][30] ),
    .B2(_05548_),
    .X(_03803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12316_ (.A1(_08462_),
    .A2(_05545_),
    .B1(\design_top.core0.REG2[1][29] ),
    .B2(_05548_),
    .X(_03802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12317_ (.A1(_08463_),
    .A2(_05545_),
    .B1(\design_top.core0.REG2[1][28] ),
    .B2(_05548_),
    .X(_03801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12318_ (.A1(_08465_),
    .A2(_05545_),
    .B1(\design_top.core0.REG2[1][27] ),
    .B2(_05548_),
    .X(_03800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12319_ (.A(_05544_),
    .X(_05549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12320_ (.A(_05547_),
    .X(_05550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12321_ (.A1(_08466_),
    .A2(_05549_),
    .B1(\design_top.core0.REG2[1][26] ),
    .B2(_05550_),
    .X(_03799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12322_ (.A1(_08468_),
    .A2(_05549_),
    .B1(\design_top.core0.REG2[1][25] ),
    .B2(_05550_),
    .X(_03798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12323_ (.A1(_08469_),
    .A2(_05549_),
    .B1(\design_top.core0.REG2[1][24] ),
    .B2(_05550_),
    .X(_03797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12324_ (.A1(_08470_),
    .A2(_05549_),
    .B1(\design_top.core0.REG2[1][23] ),
    .B2(_05550_),
    .X(_03796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12325_ (.A1(_08472_),
    .A2(_05549_),
    .B1(\design_top.core0.REG2[1][22] ),
    .B2(_05550_),
    .X(_03795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12326_ (.A(_05544_),
    .X(_05551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12327_ (.A(_05547_),
    .X(_05552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12328_ (.A1(_08473_),
    .A2(_05551_),
    .B1(\design_top.core0.REG2[1][21] ),
    .B2(_05552_),
    .X(_03794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12329_ (.A1(_08475_),
    .A2(_05551_),
    .B1(\design_top.core0.REG2[1][20] ),
    .B2(_05552_),
    .X(_03793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12330_ (.A1(_08476_),
    .A2(_05551_),
    .B1(\design_top.core0.REG2[1][19] ),
    .B2(_05552_),
    .X(_03792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12331_ (.A1(_08477_),
    .A2(_05551_),
    .B1(\design_top.core0.REG2[1][18] ),
    .B2(_05552_),
    .X(_03791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12332_ (.A1(_08479_),
    .A2(_05551_),
    .B1(\design_top.core0.REG2[1][17] ),
    .B2(_05552_),
    .X(_03790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12333_ (.A(_05543_),
    .X(_05553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12334_ (.A(_05546_),
    .X(_05554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12335_ (.A1(_08480_),
    .A2(_05553_),
    .B1(\design_top.core0.REG2[1][16] ),
    .B2(_05554_),
    .X(_03789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12336_ (.A1(_08482_),
    .A2(_05553_),
    .B1(\design_top.core0.REG2[1][15] ),
    .B2(_05554_),
    .X(_03788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12337_ (.A1(_08483_),
    .A2(_05553_),
    .B1(\design_top.core0.REG2[1][14] ),
    .B2(_05554_),
    .X(_03787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12338_ (.A1(\design_top.core0.REG2[1][13] ),
    .A2(_05544_),
    .B1(_05538_),
    .B2(_05547_),
    .X(_03786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12339_ (.A1(_08484_),
    .A2(_05553_),
    .B1(\design_top.core0.REG2[1][12] ),
    .B2(_05554_),
    .X(_03785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12340_ (.A1(_08486_),
    .A2(_05553_),
    .B1(\design_top.core0.REG2[1][11] ),
    .B2(_05554_),
    .X(_03784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12341_ (.A(_05543_),
    .X(_05555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12342_ (.A(_05546_),
    .X(_05556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12343_ (.A1(_08487_),
    .A2(_05555_),
    .B1(\design_top.core0.REG2[1][10] ),
    .B2(_05556_),
    .X(_03783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12344_ (.A1(_08489_),
    .A2(_05555_),
    .B1(\design_top.core0.REG2[1][9] ),
    .B2(_05556_),
    .X(_03782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12345_ (.A1(_08490_),
    .A2(_05555_),
    .B1(\design_top.core0.REG2[1][8] ),
    .B2(_05556_),
    .X(_03781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12346_ (.A1(_08491_),
    .A2(_05555_),
    .B1(\design_top.core0.REG2[1][7] ),
    .B2(_05556_),
    .X(_03780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12347_ (.A1(_08493_),
    .A2(_05555_),
    .B1(\design_top.core0.REG2[1][6] ),
    .B2(_05556_),
    .X(_03779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12348_ (.A(_05543_),
    .X(_05557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12349_ (.A(_05546_),
    .X(_05558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12350_ (.A1(_08494_),
    .A2(_05557_),
    .B1(\design_top.core0.REG2[1][5] ),
    .B2(_05558_),
    .X(_03778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12351_ (.A1(_08496_),
    .A2(_05557_),
    .B1(\design_top.core0.REG2[1][4] ),
    .B2(_05558_),
    .X(_03777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12352_ (.A1(_08497_),
    .A2(_05557_),
    .B1(\design_top.core0.REG2[1][3] ),
    .B2(_05558_),
    .X(_03776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12353_ (.A1(_08498_),
    .A2(_05557_),
    .B1(\design_top.core0.REG2[1][2] ),
    .B2(_05558_),
    .X(_03775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12354_ (.A1(_08499_),
    .A2(_05557_),
    .B1(\design_top.core0.REG2[1][1] ),
    .B2(_05558_),
    .X(_03774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12355_ (.A1(_08500_),
    .A2(_05544_),
    .B1(\design_top.core0.REG2[1][0] ),
    .B2(_05547_),
    .X(_03773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12356_ (.A(_08174_),
    .X(_05559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12357_ (.A(_08250_),
    .X(_05560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12358_ (.A(_05560_),
    .X(_05561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12359_ (.A(_05561_),
    .X(_05562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12360_ (.A(_05560_),
    .Y(_05563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12361_ (.A(_05563_),
    .X(_05564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12362_ (.A(_05564_),
    .X(_05565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12363_ (.A1(_05559_),
    .A2(_05562_),
    .B1(\design_top.core0.REG2[2][31] ),
    .B2(_05565_),
    .X(_03772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12364_ (.A(_08179_),
    .X(_05566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12365_ (.A1(_05566_),
    .A2(_05562_),
    .B1(\design_top.core0.REG2[2][30] ),
    .B2(_05565_),
    .X(_03771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12366_ (.A(_08181_),
    .X(_05567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12367_ (.A1(_05567_),
    .A2(_05562_),
    .B1(\design_top.core0.REG2[2][29] ),
    .B2(_05565_),
    .X(_03770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12368_ (.A(_08183_),
    .X(_05568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12369_ (.A1(_05568_),
    .A2(_05562_),
    .B1(\design_top.core0.REG2[2][28] ),
    .B2(_05565_),
    .X(_03769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12370_ (.A(_08186_),
    .X(_05569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12371_ (.A1(_05569_),
    .A2(_05562_),
    .B1(\design_top.core0.REG2[2][27] ),
    .B2(_05565_),
    .X(_03768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12372_ (.A(_08188_),
    .X(_05570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12373_ (.A(_05561_),
    .X(_05571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12374_ (.A(_05564_),
    .X(_05572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12375_ (.A1(_05570_),
    .A2(_05571_),
    .B1(\design_top.core0.REG2[2][26] ),
    .B2(_05572_),
    .X(_03767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12376_ (.A(_08191_),
    .X(_05573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12377_ (.A1(_05573_),
    .A2(_05571_),
    .B1(\design_top.core0.REG2[2][25] ),
    .B2(_05572_),
    .X(_03766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12378_ (.A(_08193_),
    .X(_05574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12379_ (.A1(_05574_),
    .A2(_05571_),
    .B1(\design_top.core0.REG2[2][24] ),
    .B2(_05572_),
    .X(_03765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12380_ (.A(_08195_),
    .X(_05575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12381_ (.A1(_05575_),
    .A2(_05571_),
    .B1(\design_top.core0.REG2[2][23] ),
    .B2(_05572_),
    .X(_03764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12382_ (.A(_08198_),
    .X(_05576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12383_ (.A1(_05576_),
    .A2(_05571_),
    .B1(\design_top.core0.REG2[2][22] ),
    .B2(_05572_),
    .X(_03763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12384_ (.A(_08200_),
    .X(_05577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12385_ (.A(_05561_),
    .X(_05578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12386_ (.A(_05564_),
    .X(_05579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12387_ (.A1(_05577_),
    .A2(_05578_),
    .B1(\design_top.core0.REG2[2][21] ),
    .B2(_05579_),
    .X(_03762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12388_ (.A(_08203_),
    .X(_05580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12389_ (.A1(_05580_),
    .A2(_05578_),
    .B1(\design_top.core0.REG2[2][20] ),
    .B2(_05579_),
    .X(_03761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12390_ (.A(_08205_),
    .X(_05581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12391_ (.A1(_05581_),
    .A2(_05578_),
    .B1(\design_top.core0.REG2[2][19] ),
    .B2(_05579_),
    .X(_03760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12392_ (.A(_08207_),
    .X(_05582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12393_ (.A1(_05582_),
    .A2(_05578_),
    .B1(\design_top.core0.REG2[2][18] ),
    .B2(_05579_),
    .X(_03759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12394_ (.A(_08210_),
    .X(_05583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12395_ (.A1(_05583_),
    .A2(_05578_),
    .B1(\design_top.core0.REG2[2][17] ),
    .B2(_05579_),
    .X(_03758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12396_ (.A(_08212_),
    .X(_05584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12397_ (.A(_05560_),
    .X(_05585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12398_ (.A(_05563_),
    .X(_05586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12399_ (.A1(_05584_),
    .A2(_05585_),
    .B1(\design_top.core0.REG2[2][16] ),
    .B2(_05586_),
    .X(_03757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12400_ (.A(_08215_),
    .X(_05587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12401_ (.A1(_05587_),
    .A2(_05585_),
    .B1(\design_top.core0.REG2[2][15] ),
    .B2(_05586_),
    .X(_03756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12402_ (.A(_08217_),
    .X(_05588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12403_ (.A1(_05588_),
    .A2(_05585_),
    .B1(\design_top.core0.REG2[2][14] ),
    .B2(_05586_),
    .X(_03755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12404_ (.A1(\design_top.core0.REG2[2][13] ),
    .A2(_05561_),
    .B1(_05538_),
    .B2(_05564_),
    .X(_03754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12405_ (.A(_08219_),
    .X(_05589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12406_ (.A1(_05589_),
    .A2(_05585_),
    .B1(\design_top.core0.REG2[2][12] ),
    .B2(_05586_),
    .X(_03753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12407_ (.A(_08222_),
    .X(_05590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12408_ (.A1(_05590_),
    .A2(_05585_),
    .B1(\design_top.core0.REG2[2][11] ),
    .B2(_05586_),
    .X(_03752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12409_ (.A(_08224_),
    .X(_05591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12410_ (.A(_05560_),
    .X(_05592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12411_ (.A(_05563_),
    .X(_05593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12412_ (.A1(_05591_),
    .A2(_05592_),
    .B1(\design_top.core0.REG2[2][10] ),
    .B2(_05593_),
    .X(_03751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12413_ (.A(_08227_),
    .X(_05594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12414_ (.A1(_05594_),
    .A2(_05592_),
    .B1(\design_top.core0.REG2[2][9] ),
    .B2(_05593_),
    .X(_03750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12415_ (.A(_08229_),
    .X(_05595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12416_ (.A1(_05595_),
    .A2(_05592_),
    .B1(\design_top.core0.REG2[2][8] ),
    .B2(_05593_),
    .X(_03749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12417_ (.A(_08231_),
    .X(_05596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12418_ (.A1(_05596_),
    .A2(_05592_),
    .B1(\design_top.core0.REG2[2][7] ),
    .B2(_05593_),
    .X(_03748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12419_ (.A(_08234_),
    .X(_05597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12420_ (.A1(_05597_),
    .A2(_05592_),
    .B1(\design_top.core0.REG2[2][6] ),
    .B2(_05593_),
    .X(_03747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12421_ (.A(_08236_),
    .X(_05598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12422_ (.A(_05560_),
    .X(_05599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12423_ (.A(_05563_),
    .X(_05600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12424_ (.A1(_05598_),
    .A2(_05599_),
    .B1(\design_top.core0.REG2[2][5] ),
    .B2(_05600_),
    .X(_03746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12425_ (.A(_08239_),
    .X(_05601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12426_ (.A1(_05601_),
    .A2(_05599_),
    .B1(\design_top.core0.REG2[2][4] ),
    .B2(_05600_),
    .X(_03745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12427_ (.A(_08241_),
    .X(_05602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12428_ (.A1(_05602_),
    .A2(_05599_),
    .B1(\design_top.core0.REG2[2][3] ),
    .B2(_05600_),
    .X(_03744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12429_ (.A(_08243_),
    .X(_05603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12430_ (.A1(_05603_),
    .A2(_05599_),
    .B1(\design_top.core0.REG2[2][2] ),
    .B2(_05600_),
    .X(_03743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12431_ (.A(_08245_),
    .X(_05604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12432_ (.A1(_05604_),
    .A2(_05599_),
    .B1(\design_top.core0.REG2[2][1] ),
    .B2(_05600_),
    .X(_03742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12433_ (.A(_08247_),
    .X(_05605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12434_ (.A1(_05605_),
    .A2(_05561_),
    .B1(\design_top.core0.REG2[2][0] ),
    .B2(_05564_),
    .X(_03741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12435_ (.A(_08267_),
    .X(_05606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12436_ (.A(_05606_),
    .X(_05607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12437_ (.A(_05607_),
    .X(_05608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12438_ (.A(_05606_),
    .Y(_05609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12439_ (.A(_05609_),
    .X(_05610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12440_ (.A(_05610_),
    .X(_05611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12441_ (.A1(_05559_),
    .A2(_05608_),
    .B1(\design_top.core0.REG2[3][31] ),
    .B2(_05611_),
    .X(_03740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12442_ (.A1(_05566_),
    .A2(_05608_),
    .B1(\design_top.core0.REG2[3][30] ),
    .B2(_05611_),
    .X(_03739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12443_ (.A1(_05567_),
    .A2(_05608_),
    .B1(\design_top.core0.REG2[3][29] ),
    .B2(_05611_),
    .X(_03738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12444_ (.A1(_05568_),
    .A2(_05608_),
    .B1(\design_top.core0.REG2[3][28] ),
    .B2(_05611_),
    .X(_03737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12445_ (.A1(_05569_),
    .A2(_05608_),
    .B1(\design_top.core0.REG2[3][27] ),
    .B2(_05611_),
    .X(_03736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12446_ (.A(_05607_),
    .X(_05612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12447_ (.A(_05610_),
    .X(_05613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12448_ (.A1(_05570_),
    .A2(_05612_),
    .B1(\design_top.core0.REG2[3][26] ),
    .B2(_05613_),
    .X(_03735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12449_ (.A1(_05573_),
    .A2(_05612_),
    .B1(\design_top.core0.REG2[3][25] ),
    .B2(_05613_),
    .X(_03734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12450_ (.A1(_05574_),
    .A2(_05612_),
    .B1(\design_top.core0.REG2[3][24] ),
    .B2(_05613_),
    .X(_03733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12451_ (.A1(_05575_),
    .A2(_05612_),
    .B1(\design_top.core0.REG2[3][23] ),
    .B2(_05613_),
    .X(_03732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12452_ (.A1(_05576_),
    .A2(_05612_),
    .B1(\design_top.core0.REG2[3][22] ),
    .B2(_05613_),
    .X(_03731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12453_ (.A(_05607_),
    .X(_05614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12454_ (.A(_05610_),
    .X(_05615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12455_ (.A1(_05577_),
    .A2(_05614_),
    .B1(\design_top.core0.REG2[3][21] ),
    .B2(_05615_),
    .X(_03730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12456_ (.A1(_05580_),
    .A2(_05614_),
    .B1(\design_top.core0.REG2[3][20] ),
    .B2(_05615_),
    .X(_03729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12457_ (.A1(_05581_),
    .A2(_05614_),
    .B1(\design_top.core0.REG2[3][19] ),
    .B2(_05615_),
    .X(_03728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12458_ (.A1(_05582_),
    .A2(_05614_),
    .B1(\design_top.core0.REG2[3][18] ),
    .B2(_05615_),
    .X(_03727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12459_ (.A1(_05583_),
    .A2(_05614_),
    .B1(\design_top.core0.REG2[3][17] ),
    .B2(_05615_),
    .X(_03726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12460_ (.A(_05606_),
    .X(_05616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12461_ (.A(_05609_),
    .X(_05617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12462_ (.A1(_05584_),
    .A2(_05616_),
    .B1(\design_top.core0.REG2[3][16] ),
    .B2(_05617_),
    .X(_03725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12463_ (.A1(_05587_),
    .A2(_05616_),
    .B1(\design_top.core0.REG2[3][15] ),
    .B2(_05617_),
    .X(_03724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12464_ (.A1(_05588_),
    .A2(_05616_),
    .B1(\design_top.core0.REG2[3][14] ),
    .B2(_05617_),
    .X(_03723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12465_ (.A1(\design_top.core0.REG2[3][13] ),
    .A2(_05607_),
    .B1(_05538_),
    .B2(_05610_),
    .X(_03722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12466_ (.A1(_05589_),
    .A2(_05616_),
    .B1(\design_top.core0.REG2[3][12] ),
    .B2(_05617_),
    .X(_03721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12467_ (.A1(_05590_),
    .A2(_05616_),
    .B1(\design_top.core0.REG2[3][11] ),
    .B2(_05617_),
    .X(_03720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12468_ (.A(_05606_),
    .X(_05618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12469_ (.A(_05609_),
    .X(_05619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12470_ (.A1(_05591_),
    .A2(_05618_),
    .B1(\design_top.core0.REG2[3][10] ),
    .B2(_05619_),
    .X(_03719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12471_ (.A1(_05594_),
    .A2(_05618_),
    .B1(\design_top.core0.REG2[3][9] ),
    .B2(_05619_),
    .X(_03718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12472_ (.A1(_05595_),
    .A2(_05618_),
    .B1(\design_top.core0.REG2[3][8] ),
    .B2(_05619_),
    .X(_03717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12473_ (.A1(_05596_),
    .A2(_05618_),
    .B1(\design_top.core0.REG2[3][7] ),
    .B2(_05619_),
    .X(_03716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12474_ (.A1(_05597_),
    .A2(_05618_),
    .B1(\design_top.core0.REG2[3][6] ),
    .B2(_05619_),
    .X(_03715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12475_ (.A(_05606_),
    .X(_05620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12476_ (.A(_05609_),
    .X(_05621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12477_ (.A1(_05598_),
    .A2(_05620_),
    .B1(\design_top.core0.REG2[3][5] ),
    .B2(_05621_),
    .X(_03714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12478_ (.A1(_05601_),
    .A2(_05620_),
    .B1(\design_top.core0.REG2[3][4] ),
    .B2(_05621_),
    .X(_03713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12479_ (.A1(_05602_),
    .A2(_05620_),
    .B1(\design_top.core0.REG2[3][3] ),
    .B2(_05621_),
    .X(_03712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12480_ (.A1(_05603_),
    .A2(_05620_),
    .B1(\design_top.core0.REG2[3][2] ),
    .B2(_05621_),
    .X(_03711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12481_ (.A1(_05604_),
    .A2(_05620_),
    .B1(\design_top.core0.REG2[3][1] ),
    .B2(_05621_),
    .X(_03710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12482_ (.A1(_05605_),
    .A2(_05607_),
    .B1(\design_top.core0.REG2[3][0] ),
    .B2(_05610_),
    .X(_03709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12483_ (.A(_08284_),
    .X(_05622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12484_ (.A(_05622_),
    .X(_05623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12485_ (.A(_05623_),
    .X(_05624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12486_ (.A(_05622_),
    .Y(_05625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12487_ (.A(_05625_),
    .X(_05626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12488_ (.A(_05626_),
    .X(_05627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12489_ (.A1(_05559_),
    .A2(_05624_),
    .B1(\design_top.core0.REG2[4][31] ),
    .B2(_05627_),
    .X(_03708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12490_ (.A1(_05566_),
    .A2(_05624_),
    .B1(\design_top.core0.REG2[4][30] ),
    .B2(_05627_),
    .X(_03707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12491_ (.A1(_05567_),
    .A2(_05624_),
    .B1(\design_top.core0.REG2[4][29] ),
    .B2(_05627_),
    .X(_03706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12492_ (.A1(_05568_),
    .A2(_05624_),
    .B1(\design_top.core0.REG2[4][28] ),
    .B2(_05627_),
    .X(_03705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12493_ (.A1(_05569_),
    .A2(_05624_),
    .B1(\design_top.core0.REG2[4][27] ),
    .B2(_05627_),
    .X(_03704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12494_ (.A(_05623_),
    .X(_05628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12495_ (.A(_05626_),
    .X(_05629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12496_ (.A1(_05570_),
    .A2(_05628_),
    .B1(\design_top.core0.REG2[4][26] ),
    .B2(_05629_),
    .X(_03703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12497_ (.A1(_05573_),
    .A2(_05628_),
    .B1(\design_top.core0.REG2[4][25] ),
    .B2(_05629_),
    .X(_03702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12498_ (.A1(_05574_),
    .A2(_05628_),
    .B1(\design_top.core0.REG2[4][24] ),
    .B2(_05629_),
    .X(_03701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12499_ (.A1(_05575_),
    .A2(_05628_),
    .B1(\design_top.core0.REG2[4][23] ),
    .B2(_05629_),
    .X(_03700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12500_ (.A1(_05576_),
    .A2(_05628_),
    .B1(\design_top.core0.REG2[4][22] ),
    .B2(_05629_),
    .X(_03699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12501_ (.A(_05623_),
    .X(_05630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12502_ (.A(_05626_),
    .X(_05631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12503_ (.A1(_05577_),
    .A2(_05630_),
    .B1(\design_top.core0.REG2[4][21] ),
    .B2(_05631_),
    .X(_03698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12504_ (.A1(_05580_),
    .A2(_05630_),
    .B1(\design_top.core0.REG2[4][20] ),
    .B2(_05631_),
    .X(_03697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12505_ (.A1(_05581_),
    .A2(_05630_),
    .B1(\design_top.core0.REG2[4][19] ),
    .B2(_05631_),
    .X(_03696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12506_ (.A1(_05582_),
    .A2(_05630_),
    .B1(\design_top.core0.REG2[4][18] ),
    .B2(_05631_),
    .X(_03695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12507_ (.A1(_05583_),
    .A2(_05630_),
    .B1(\design_top.core0.REG2[4][17] ),
    .B2(_05631_),
    .X(_03694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12508_ (.A(_05622_),
    .X(_05632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12509_ (.A(_05625_),
    .X(_05633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12510_ (.A1(_05584_),
    .A2(_05632_),
    .B1(\design_top.core0.REG2[4][16] ),
    .B2(_05633_),
    .X(_03693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12511_ (.A1(_05587_),
    .A2(_05632_),
    .B1(\design_top.core0.REG2[4][15] ),
    .B2(_05633_),
    .X(_03692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12512_ (.A1(_05588_),
    .A2(_05632_),
    .B1(\design_top.core0.REG2[4][14] ),
    .B2(_05633_),
    .X(_03691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12513_ (.A1(\design_top.core0.REG2[4][13] ),
    .A2(_05623_),
    .B1(_05538_),
    .B2(_05626_),
    .X(_03690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12514_ (.A1(_05589_),
    .A2(_05632_),
    .B1(\design_top.core0.REG2[4][12] ),
    .B2(_05633_),
    .X(_03689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12515_ (.A1(_05590_),
    .A2(_05632_),
    .B1(\design_top.core0.REG2[4][11] ),
    .B2(_05633_),
    .X(_03688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12516_ (.A(_05622_),
    .X(_05634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12517_ (.A(_05625_),
    .X(_05635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12518_ (.A1(_05591_),
    .A2(_05634_),
    .B1(\design_top.core0.REG2[4][10] ),
    .B2(_05635_),
    .X(_03687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12519_ (.A1(_05594_),
    .A2(_05634_),
    .B1(\design_top.core0.REG2[4][9] ),
    .B2(_05635_),
    .X(_03686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12520_ (.A1(_05595_),
    .A2(_05634_),
    .B1(\design_top.core0.REG2[4][8] ),
    .B2(_05635_),
    .X(_03685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12521_ (.A1(_05596_),
    .A2(_05634_),
    .B1(\design_top.core0.REG2[4][7] ),
    .B2(_05635_),
    .X(_03684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12522_ (.A1(_05597_),
    .A2(_05634_),
    .B1(\design_top.core0.REG2[4][6] ),
    .B2(_05635_),
    .X(_03683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12523_ (.A(_05622_),
    .X(_05636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12524_ (.A(_05625_),
    .X(_05637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12525_ (.A1(_05598_),
    .A2(_05636_),
    .B1(\design_top.core0.REG2[4][5] ),
    .B2(_05637_),
    .X(_03682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12526_ (.A1(_05601_),
    .A2(_05636_),
    .B1(\design_top.core0.REG2[4][4] ),
    .B2(_05637_),
    .X(_03681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12527_ (.A1(_05602_),
    .A2(_05636_),
    .B1(\design_top.core0.REG2[4][3] ),
    .B2(_05637_),
    .X(_03680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12528_ (.A1(_05603_),
    .A2(_05636_),
    .B1(\design_top.core0.REG2[4][2] ),
    .B2(_05637_),
    .X(_03679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12529_ (.A1(_05604_),
    .A2(_05636_),
    .B1(\design_top.core0.REG2[4][1] ),
    .B2(_05637_),
    .X(_03678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12530_ (.A1(_05605_),
    .A2(_05623_),
    .B1(\design_top.core0.REG2[4][0] ),
    .B2(_05626_),
    .X(_03677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12531_ (.A(_08022_),
    .X(_05638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12532_ (.A1(_08045_),
    .A2(_07131_),
    .B1(_07353_),
    .B2(_05638_),
    .X(_05639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12533_ (.A(_05639_),
    .Y(_05640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12534_ (.A(_05640_),
    .X(_05641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12535_ (.A(_05639_),
    .X(_05642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12536_ (.A1(_00412_),
    .A2(_05641_),
    .B1(\design_top.MEM[7][7] ),
    .B2(_05642_),
    .X(_03676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12537_ (.A1(_00411_),
    .A2(_05641_),
    .B1(\design_top.MEM[7][6] ),
    .B2(_05642_),
    .X(_03675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12538_ (.A1(_00410_),
    .A2(_05641_),
    .B1(\design_top.MEM[7][5] ),
    .B2(_05642_),
    .X(_03674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12539_ (.A1(_00409_),
    .A2(_05641_),
    .B1(\design_top.MEM[7][4] ),
    .B2(_05642_),
    .X(_03673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12540_ (.A1(_00408_),
    .A2(_05641_),
    .B1(\design_top.MEM[7][3] ),
    .B2(_05642_),
    .X(_03672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12541_ (.A1(_00407_),
    .A2(_05640_),
    .B1(\design_top.MEM[7][2] ),
    .B2(_05639_),
    .X(_03671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12542_ (.A1(_00406_),
    .A2(_05640_),
    .B1(\design_top.MEM[7][1] ),
    .B2(_05639_),
    .X(_03670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12543_ (.A1(_00405_),
    .A2(_05640_),
    .B1(\design_top.MEM[7][0] ),
    .B2(_05639_),
    .X(_03669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12544_ (.A(_08303_),
    .X(_05643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12545_ (.A(_05643_),
    .X(_05644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12546_ (.A(_05644_),
    .X(_05645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12547_ (.A(_05643_),
    .Y(_05646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12548_ (.A(_05646_),
    .X(_05647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12549_ (.A(_05647_),
    .X(_05648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12550_ (.A1(_05559_),
    .A2(_05645_),
    .B1(\design_top.core0.REG2[5][31] ),
    .B2(_05648_),
    .X(_03668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12551_ (.A1(_05566_),
    .A2(_05645_),
    .B1(\design_top.core0.REG2[5][30] ),
    .B2(_05648_),
    .X(_03667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12552_ (.A1(_05567_),
    .A2(_05645_),
    .B1(\design_top.core0.REG2[5][29] ),
    .B2(_05648_),
    .X(_03666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12553_ (.A1(_05568_),
    .A2(_05645_),
    .B1(\design_top.core0.REG2[5][28] ),
    .B2(_05648_),
    .X(_03665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12554_ (.A1(_05569_),
    .A2(_05645_),
    .B1(\design_top.core0.REG2[5][27] ),
    .B2(_05648_),
    .X(_03664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12555_ (.A(_05644_),
    .X(_05649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12556_ (.A(_05647_),
    .X(_05650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12557_ (.A1(_05570_),
    .A2(_05649_),
    .B1(\design_top.core0.REG2[5][26] ),
    .B2(_05650_),
    .X(_03663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12558_ (.A1(_05573_),
    .A2(_05649_),
    .B1(\design_top.core0.REG2[5][25] ),
    .B2(_05650_),
    .X(_03662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12559_ (.A1(_05574_),
    .A2(_05649_),
    .B1(\design_top.core0.REG2[5][24] ),
    .B2(_05650_),
    .X(_03661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12560_ (.A1(_05575_),
    .A2(_05649_),
    .B1(\design_top.core0.REG2[5][23] ),
    .B2(_05650_),
    .X(_03660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12561_ (.A1(_05576_),
    .A2(_05649_),
    .B1(\design_top.core0.REG2[5][22] ),
    .B2(_05650_),
    .X(_03659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12562_ (.A(_05644_),
    .X(_05651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12563_ (.A(_05647_),
    .X(_05652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12564_ (.A1(_05577_),
    .A2(_05651_),
    .B1(\design_top.core0.REG2[5][21] ),
    .B2(_05652_),
    .X(_03658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12565_ (.A1(_05580_),
    .A2(_05651_),
    .B1(\design_top.core0.REG2[5][20] ),
    .B2(_05652_),
    .X(_03657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12566_ (.A1(_05581_),
    .A2(_05651_),
    .B1(\design_top.core0.REG2[5][19] ),
    .B2(_05652_),
    .X(_03656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12567_ (.A1(_05582_),
    .A2(_05651_),
    .B1(\design_top.core0.REG2[5][18] ),
    .B2(_05652_),
    .X(_03655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12568_ (.A1(_05583_),
    .A2(_05651_),
    .B1(\design_top.core0.REG2[5][17] ),
    .B2(_05652_),
    .X(_03654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12569_ (.A(_05643_),
    .X(_05653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12570_ (.A(_05646_),
    .X(_05654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12571_ (.A1(_05584_),
    .A2(_05653_),
    .B1(\design_top.core0.REG2[5][16] ),
    .B2(_05654_),
    .X(_03653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12572_ (.A1(_05587_),
    .A2(_05653_),
    .B1(\design_top.core0.REG2[5][15] ),
    .B2(_05654_),
    .X(_03652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12573_ (.A1(_05588_),
    .A2(_05653_),
    .B1(\design_top.core0.REG2[5][14] ),
    .B2(_05654_),
    .X(_03651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12574_ (.A(_08531_),
    .X(_05655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12575_ (.A1(\design_top.core0.REG2[5][13] ),
    .A2(_05644_),
    .B1(_05655_),
    .B2(_05647_),
    .X(_03650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12576_ (.A1(_05589_),
    .A2(_05653_),
    .B1(\design_top.core0.REG2[5][12] ),
    .B2(_05654_),
    .X(_03649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12577_ (.A1(_05590_),
    .A2(_05653_),
    .B1(\design_top.core0.REG2[5][11] ),
    .B2(_05654_),
    .X(_03648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12578_ (.A(_05643_),
    .X(_05656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12579_ (.A(_05646_),
    .X(_05657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12580_ (.A1(_05591_),
    .A2(_05656_),
    .B1(\design_top.core0.REG2[5][10] ),
    .B2(_05657_),
    .X(_03647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12581_ (.A1(_05594_),
    .A2(_05656_),
    .B1(\design_top.core0.REG2[5][9] ),
    .B2(_05657_),
    .X(_03646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12582_ (.A1(_05595_),
    .A2(_05656_),
    .B1(\design_top.core0.REG2[5][8] ),
    .B2(_05657_),
    .X(_03645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12583_ (.A1(_05596_),
    .A2(_05656_),
    .B1(\design_top.core0.REG2[5][7] ),
    .B2(_05657_),
    .X(_03644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12584_ (.A1(_05597_),
    .A2(_05656_),
    .B1(\design_top.core0.REG2[5][6] ),
    .B2(_05657_),
    .X(_03643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12585_ (.A(_05643_),
    .X(_05658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12586_ (.A(_05646_),
    .X(_05659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12587_ (.A1(_05598_),
    .A2(_05658_),
    .B1(\design_top.core0.REG2[5][5] ),
    .B2(_05659_),
    .X(_03642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12588_ (.A1(_05601_),
    .A2(_05658_),
    .B1(\design_top.core0.REG2[5][4] ),
    .B2(_05659_),
    .X(_03641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12589_ (.A1(_05602_),
    .A2(_05658_),
    .B1(\design_top.core0.REG2[5][3] ),
    .B2(_05659_),
    .X(_03640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12590_ (.A1(_05603_),
    .A2(_05658_),
    .B1(\design_top.core0.REG2[5][2] ),
    .B2(_05659_),
    .X(_03639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12591_ (.A1(_05604_),
    .A2(_05658_),
    .B1(\design_top.core0.REG2[5][1] ),
    .B2(_05659_),
    .X(_03638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12592_ (.A1(_05605_),
    .A2(_05644_),
    .B1(\design_top.core0.REG2[5][0] ),
    .B2(_05647_),
    .X(_03637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12593_ (.A(_08320_),
    .X(_05660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12594_ (.A(_05660_),
    .X(_05661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12595_ (.A(_05661_),
    .X(_05662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12596_ (.A(_05660_),
    .Y(_05663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12597_ (.A(_05663_),
    .X(_05664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12598_ (.A(_05664_),
    .X(_05665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12599_ (.A1(_05559_),
    .A2(_05662_),
    .B1(\design_top.core0.REG2[6][31] ),
    .B2(_05665_),
    .X(_03636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12600_ (.A1(_05566_),
    .A2(_05662_),
    .B1(\design_top.core0.REG2[6][30] ),
    .B2(_05665_),
    .X(_03635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12601_ (.A1(_05567_),
    .A2(_05662_),
    .B1(\design_top.core0.REG2[6][29] ),
    .B2(_05665_),
    .X(_03634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12602_ (.A1(_05568_),
    .A2(_05662_),
    .B1(\design_top.core0.REG2[6][28] ),
    .B2(_05665_),
    .X(_03633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12603_ (.A1(_05569_),
    .A2(_05662_),
    .B1(\design_top.core0.REG2[6][27] ),
    .B2(_05665_),
    .X(_03632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12604_ (.A(_05661_),
    .X(_05666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12605_ (.A(_05664_),
    .X(_05667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12606_ (.A1(_05570_),
    .A2(_05666_),
    .B1(\design_top.core0.REG2[6][26] ),
    .B2(_05667_),
    .X(_03631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12607_ (.A1(_05573_),
    .A2(_05666_),
    .B1(\design_top.core0.REG2[6][25] ),
    .B2(_05667_),
    .X(_03630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12608_ (.A1(_05574_),
    .A2(_05666_),
    .B1(\design_top.core0.REG2[6][24] ),
    .B2(_05667_),
    .X(_03629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12609_ (.A1(_05575_),
    .A2(_05666_),
    .B1(\design_top.core0.REG2[6][23] ),
    .B2(_05667_),
    .X(_03628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12610_ (.A1(_05576_),
    .A2(_05666_),
    .B1(\design_top.core0.REG2[6][22] ),
    .B2(_05667_),
    .X(_03627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12611_ (.A(_05661_),
    .X(_05668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12612_ (.A(_05664_),
    .X(_05669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12613_ (.A1(_05577_),
    .A2(_05668_),
    .B1(\design_top.core0.REG2[6][21] ),
    .B2(_05669_),
    .X(_03626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12614_ (.A1(_05580_),
    .A2(_05668_),
    .B1(\design_top.core0.REG2[6][20] ),
    .B2(_05669_),
    .X(_03625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12615_ (.A1(_05581_),
    .A2(_05668_),
    .B1(\design_top.core0.REG2[6][19] ),
    .B2(_05669_),
    .X(_03624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12616_ (.A1(_05582_),
    .A2(_05668_),
    .B1(\design_top.core0.REG2[6][18] ),
    .B2(_05669_),
    .X(_03623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12617_ (.A1(_05583_),
    .A2(_05668_),
    .B1(\design_top.core0.REG2[6][17] ),
    .B2(_05669_),
    .X(_03622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12618_ (.A(_05660_),
    .X(_05670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12619_ (.A(_05663_),
    .X(_05671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12620_ (.A1(_05584_),
    .A2(_05670_),
    .B1(\design_top.core0.REG2[6][16] ),
    .B2(_05671_),
    .X(_03621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12621_ (.A1(_05587_),
    .A2(_05670_),
    .B1(\design_top.core0.REG2[6][15] ),
    .B2(_05671_),
    .X(_03620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12622_ (.A1(_05588_),
    .A2(_05670_),
    .B1(\design_top.core0.REG2[6][14] ),
    .B2(_05671_),
    .X(_03619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12623_ (.A1(\design_top.core0.REG2[6][13] ),
    .A2(_05661_),
    .B1(_05655_),
    .B2(_05664_),
    .X(_03618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12624_ (.A1(_05589_),
    .A2(_05670_),
    .B1(\design_top.core0.REG2[6][12] ),
    .B2(_05671_),
    .X(_03617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12625_ (.A1(_05590_),
    .A2(_05670_),
    .B1(\design_top.core0.REG2[6][11] ),
    .B2(_05671_),
    .X(_03616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12626_ (.A(_05660_),
    .X(_05672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12627_ (.A(_05663_),
    .X(_05673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12628_ (.A1(_05591_),
    .A2(_05672_),
    .B1(\design_top.core0.REG2[6][10] ),
    .B2(_05673_),
    .X(_03615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12629_ (.A1(_05594_),
    .A2(_05672_),
    .B1(\design_top.core0.REG2[6][9] ),
    .B2(_05673_),
    .X(_03614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12630_ (.A1(_05595_),
    .A2(_05672_),
    .B1(\design_top.core0.REG2[6][8] ),
    .B2(_05673_),
    .X(_03613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12631_ (.A1(_05596_),
    .A2(_05672_),
    .B1(\design_top.core0.REG2[6][7] ),
    .B2(_05673_),
    .X(_03612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12632_ (.A1(_05597_),
    .A2(_05672_),
    .B1(\design_top.core0.REG2[6][6] ),
    .B2(_05673_),
    .X(_03611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12633_ (.A(_05660_),
    .X(_05674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12634_ (.A(_05663_),
    .X(_05675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12635_ (.A1(_05598_),
    .A2(_05674_),
    .B1(\design_top.core0.REG2[6][5] ),
    .B2(_05675_),
    .X(_03610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12636_ (.A1(_05601_),
    .A2(_05674_),
    .B1(\design_top.core0.REG2[6][4] ),
    .B2(_05675_),
    .X(_03609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12637_ (.A1(_05602_),
    .A2(_05674_),
    .B1(\design_top.core0.REG2[6][3] ),
    .B2(_05675_),
    .X(_03608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12638_ (.A1(_05603_),
    .A2(_05674_),
    .B1(\design_top.core0.REG2[6][2] ),
    .B2(_05675_),
    .X(_03607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12639_ (.A1(_05604_),
    .A2(_05674_),
    .B1(\design_top.core0.REG2[6][1] ),
    .B2(_05675_),
    .X(_03606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12640_ (.A1(_05605_),
    .A2(_05661_),
    .B1(\design_top.core0.REG2[6][0] ),
    .B2(_05664_),
    .X(_03605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12641_ (.A(_08174_),
    .X(_05676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12642_ (.A(_08368_),
    .X(_05677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12643_ (.A(_05677_),
    .X(_05678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12644_ (.A(_05678_),
    .X(_05679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12645_ (.A(_05677_),
    .Y(_05680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12646_ (.A(_05680_),
    .X(_05681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12647_ (.A(_05681_),
    .X(_05682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12648_ (.A1(_05676_),
    .A2(_05679_),
    .B1(\design_top.core0.REG2[7][31] ),
    .B2(_05682_),
    .X(_03604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12649_ (.A(_08179_),
    .X(_05683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12650_ (.A1(_05683_),
    .A2(_05679_),
    .B1(\design_top.core0.REG2[7][30] ),
    .B2(_05682_),
    .X(_03603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12651_ (.A(_08181_),
    .X(_05684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12652_ (.A1(_05684_),
    .A2(_05679_),
    .B1(\design_top.core0.REG2[7][29] ),
    .B2(_05682_),
    .X(_03602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12653_ (.A(_08183_),
    .X(_05685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12654_ (.A1(_05685_),
    .A2(_05679_),
    .B1(\design_top.core0.REG2[7][28] ),
    .B2(_05682_),
    .X(_03601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12655_ (.A(_08186_),
    .X(_05686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12656_ (.A1(_05686_),
    .A2(_05679_),
    .B1(\design_top.core0.REG2[7][27] ),
    .B2(_05682_),
    .X(_03600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12657_ (.A(_08188_),
    .X(_05687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12658_ (.A(_05678_),
    .X(_05688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12659_ (.A(_05681_),
    .X(_05689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12660_ (.A1(_05687_),
    .A2(_05688_),
    .B1(\design_top.core0.REG2[7][26] ),
    .B2(_05689_),
    .X(_03599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12661_ (.A(_08191_),
    .X(_05690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12662_ (.A1(_05690_),
    .A2(_05688_),
    .B1(\design_top.core0.REG2[7][25] ),
    .B2(_05689_),
    .X(_03598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12663_ (.A(_08193_),
    .X(_05691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12664_ (.A1(_05691_),
    .A2(_05688_),
    .B1(\design_top.core0.REG2[7][24] ),
    .B2(_05689_),
    .X(_03597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12665_ (.A(_08195_),
    .X(_05692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12666_ (.A1(_05692_),
    .A2(_05688_),
    .B1(\design_top.core0.REG2[7][23] ),
    .B2(_05689_),
    .X(_03596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12667_ (.A(_08198_),
    .X(_05693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12668_ (.A1(_05693_),
    .A2(_05688_),
    .B1(\design_top.core0.REG2[7][22] ),
    .B2(_05689_),
    .X(_03595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12669_ (.A(_08200_),
    .X(_05694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12670_ (.A(_05678_),
    .X(_05695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12671_ (.A(_05681_),
    .X(_05696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12672_ (.A1(_05694_),
    .A2(_05695_),
    .B1(\design_top.core0.REG2[7][21] ),
    .B2(_05696_),
    .X(_03594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12673_ (.A(_08203_),
    .X(_05697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12674_ (.A1(_05697_),
    .A2(_05695_),
    .B1(\design_top.core0.REG2[7][20] ),
    .B2(_05696_),
    .X(_03593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12675_ (.A(_08205_),
    .X(_05698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12676_ (.A1(_05698_),
    .A2(_05695_),
    .B1(\design_top.core0.REG2[7][19] ),
    .B2(_05696_),
    .X(_03592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12677_ (.A(_08207_),
    .X(_05699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12678_ (.A1(_05699_),
    .A2(_05695_),
    .B1(\design_top.core0.REG2[7][18] ),
    .B2(_05696_),
    .X(_03591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12679_ (.A(_08210_),
    .X(_05700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12680_ (.A1(_05700_),
    .A2(_05695_),
    .B1(\design_top.core0.REG2[7][17] ),
    .B2(_05696_),
    .X(_03590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12681_ (.A(_08212_),
    .X(_05701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12682_ (.A(_05677_),
    .X(_05702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12683_ (.A(_05680_),
    .X(_05703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12684_ (.A1(_05701_),
    .A2(_05702_),
    .B1(\design_top.core0.REG2[7][16] ),
    .B2(_05703_),
    .X(_03589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12685_ (.A(_08215_),
    .X(_05704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12686_ (.A1(_05704_),
    .A2(_05702_),
    .B1(\design_top.core0.REG2[7][15] ),
    .B2(_05703_),
    .X(_03588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12687_ (.A(_08217_),
    .X(_05705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12688_ (.A1(_05705_),
    .A2(_05702_),
    .B1(\design_top.core0.REG2[7][14] ),
    .B2(_05703_),
    .X(_03587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12689_ (.A1(\design_top.core0.REG2[7][13] ),
    .A2(_05678_),
    .B1(_05655_),
    .B2(_05681_),
    .X(_03586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12690_ (.A(_08219_),
    .X(_05706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12691_ (.A1(_05706_),
    .A2(_05702_),
    .B1(\design_top.core0.REG2[7][12] ),
    .B2(_05703_),
    .X(_03585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12692_ (.A(_08222_),
    .X(_05707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12693_ (.A1(_05707_),
    .A2(_05702_),
    .B1(\design_top.core0.REG2[7][11] ),
    .B2(_05703_),
    .X(_03584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12694_ (.A(_08224_),
    .X(_05708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12695_ (.A(_05677_),
    .X(_05709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12696_ (.A(_05680_),
    .X(_05710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12697_ (.A1(_05708_),
    .A2(_05709_),
    .B1(\design_top.core0.REG2[7][10] ),
    .B2(_05710_),
    .X(_03583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12698_ (.A(_08227_),
    .X(_05711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12699_ (.A1(_05711_),
    .A2(_05709_),
    .B1(\design_top.core0.REG2[7][9] ),
    .B2(_05710_),
    .X(_03582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12700_ (.A(_08229_),
    .X(_05712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12701_ (.A1(_05712_),
    .A2(_05709_),
    .B1(\design_top.core0.REG2[7][8] ),
    .B2(_05710_),
    .X(_03581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12702_ (.A(_08231_),
    .X(_05713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12703_ (.A1(_05713_),
    .A2(_05709_),
    .B1(\design_top.core0.REG2[7][7] ),
    .B2(_05710_),
    .X(_03580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12704_ (.A(_08234_),
    .X(_05714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12705_ (.A1(_05714_),
    .A2(_05709_),
    .B1(\design_top.core0.REG2[7][6] ),
    .B2(_05710_),
    .X(_03579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12706_ (.A(_08236_),
    .X(_05715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12707_ (.A(_05677_),
    .X(_05716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12708_ (.A(_05680_),
    .X(_05717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12709_ (.A1(_05715_),
    .A2(_05716_),
    .B1(\design_top.core0.REG2[7][5] ),
    .B2(_05717_),
    .X(_03578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12710_ (.A(_08239_),
    .X(_05718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12711_ (.A1(_05718_),
    .A2(_05716_),
    .B1(\design_top.core0.REG2[7][4] ),
    .B2(_05717_),
    .X(_03577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12712_ (.A(_08241_),
    .X(_05719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12713_ (.A1(_05719_),
    .A2(_05716_),
    .B1(\design_top.core0.REG2[7][3] ),
    .B2(_05717_),
    .X(_03576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12714_ (.A(_08243_),
    .X(_05720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12715_ (.A1(_05720_),
    .A2(_05716_),
    .B1(\design_top.core0.REG2[7][2] ),
    .B2(_05717_),
    .X(_03575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12716_ (.A(_08245_),
    .X(_05721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12717_ (.A1(_05721_),
    .A2(_05716_),
    .B1(\design_top.core0.REG2[7][1] ),
    .B2(_05717_),
    .X(_03574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12718_ (.A(_08247_),
    .X(_05722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12719_ (.A1(_05722_),
    .A2(_05678_),
    .B1(\design_top.core0.REG2[7][0] ),
    .B2(_05681_),
    .X(_03573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12720_ (.A(_08390_),
    .X(_05723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12721_ (.A(_05723_),
    .X(_05724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12722_ (.A(_05724_),
    .X(_05725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12723_ (.A(_05723_),
    .Y(_05726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12724_ (.A(_05726_),
    .X(_05727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12725_ (.A(_05727_),
    .X(_05728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12726_ (.A1(_05676_),
    .A2(_05725_),
    .B1(\design_top.core0.REG2[8][31] ),
    .B2(_05728_),
    .X(_03572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12727_ (.A1(_05683_),
    .A2(_05725_),
    .B1(\design_top.core0.REG2[8][30] ),
    .B2(_05728_),
    .X(_03571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12728_ (.A1(_05684_),
    .A2(_05725_),
    .B1(\design_top.core0.REG2[8][29] ),
    .B2(_05728_),
    .X(_03570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12729_ (.A1(_05685_),
    .A2(_05725_),
    .B1(\design_top.core0.REG2[8][28] ),
    .B2(_05728_),
    .X(_03569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12730_ (.A1(_05686_),
    .A2(_05725_),
    .B1(\design_top.core0.REG2[8][27] ),
    .B2(_05728_),
    .X(_03568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12731_ (.A(_05724_),
    .X(_05729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12732_ (.A(_05727_),
    .X(_05730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12733_ (.A1(_05687_),
    .A2(_05729_),
    .B1(\design_top.core0.REG2[8][26] ),
    .B2(_05730_),
    .X(_03567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12734_ (.A1(_05690_),
    .A2(_05729_),
    .B1(\design_top.core0.REG2[8][25] ),
    .B2(_05730_),
    .X(_03566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12735_ (.A1(_05691_),
    .A2(_05729_),
    .B1(\design_top.core0.REG2[8][24] ),
    .B2(_05730_),
    .X(_03565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12736_ (.A1(_05692_),
    .A2(_05729_),
    .B1(\design_top.core0.REG2[8][23] ),
    .B2(_05730_),
    .X(_03564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12737_ (.A1(_05693_),
    .A2(_05729_),
    .B1(\design_top.core0.REG2[8][22] ),
    .B2(_05730_),
    .X(_03563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12738_ (.A(_05724_),
    .X(_05731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12739_ (.A(_05727_),
    .X(_05732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12740_ (.A1(_05694_),
    .A2(_05731_),
    .B1(\design_top.core0.REG2[8][21] ),
    .B2(_05732_),
    .X(_03562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12741_ (.A1(_05697_),
    .A2(_05731_),
    .B1(\design_top.core0.REG2[8][20] ),
    .B2(_05732_),
    .X(_03561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12742_ (.A1(_05698_),
    .A2(_05731_),
    .B1(\design_top.core0.REG2[8][19] ),
    .B2(_05732_),
    .X(_03560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12743_ (.A1(_05699_),
    .A2(_05731_),
    .B1(\design_top.core0.REG2[8][18] ),
    .B2(_05732_),
    .X(_03559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12744_ (.A1(_05700_),
    .A2(_05731_),
    .B1(\design_top.core0.REG2[8][17] ),
    .B2(_05732_),
    .X(_03558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12745_ (.A(_05723_),
    .X(_05733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12746_ (.A(_05726_),
    .X(_05734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12747_ (.A1(_05701_),
    .A2(_05733_),
    .B1(\design_top.core0.REG2[8][16] ),
    .B2(_05734_),
    .X(_03557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12748_ (.A1(_05704_),
    .A2(_05733_),
    .B1(\design_top.core0.REG2[8][15] ),
    .B2(_05734_),
    .X(_03556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12749_ (.A1(_05705_),
    .A2(_05733_),
    .B1(\design_top.core0.REG2[8][14] ),
    .B2(_05734_),
    .X(_03555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12750_ (.A1(\design_top.core0.REG2[8][13] ),
    .A2(_05724_),
    .B1(_05655_),
    .B2(_05727_),
    .X(_03554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12751_ (.A1(_05706_),
    .A2(_05733_),
    .B1(\design_top.core0.REG2[8][12] ),
    .B2(_05734_),
    .X(_03553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12752_ (.A1(_05707_),
    .A2(_05733_),
    .B1(\design_top.core0.REG2[8][11] ),
    .B2(_05734_),
    .X(_03552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12753_ (.A(_05723_),
    .X(_05735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12754_ (.A(_05726_),
    .X(_05736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12755_ (.A1(_05708_),
    .A2(_05735_),
    .B1(\design_top.core0.REG2[8][10] ),
    .B2(_05736_),
    .X(_03551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12756_ (.A1(_05711_),
    .A2(_05735_),
    .B1(\design_top.core0.REG2[8][9] ),
    .B2(_05736_),
    .X(_03550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12757_ (.A1(_05712_),
    .A2(_05735_),
    .B1(\design_top.core0.REG2[8][8] ),
    .B2(_05736_),
    .X(_03549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12758_ (.A1(_05713_),
    .A2(_05735_),
    .B1(\design_top.core0.REG2[8][7] ),
    .B2(_05736_),
    .X(_03548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12759_ (.A1(_05714_),
    .A2(_05735_),
    .B1(\design_top.core0.REG2[8][6] ),
    .B2(_05736_),
    .X(_03547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12760_ (.A(_05723_),
    .X(_05737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12761_ (.A(_05726_),
    .X(_05738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12762_ (.A1(_05715_),
    .A2(_05737_),
    .B1(\design_top.core0.REG2[8][5] ),
    .B2(_05738_),
    .X(_03546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12763_ (.A1(_05718_),
    .A2(_05737_),
    .B1(\design_top.core0.REG2[8][4] ),
    .B2(_05738_),
    .X(_03545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12764_ (.A1(_05719_),
    .A2(_05737_),
    .B1(\design_top.core0.REG2[8][3] ),
    .B2(_05738_),
    .X(_03544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12765_ (.A1(_05720_),
    .A2(_05737_),
    .B1(\design_top.core0.REG2[8][2] ),
    .B2(_05738_),
    .X(_03543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12766_ (.A1(_05721_),
    .A2(_05737_),
    .B1(\design_top.core0.REG2[8][1] ),
    .B2(_05738_),
    .X(_03542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12767_ (.A1(_05722_),
    .A2(_05724_),
    .B1(\design_top.core0.REG2[8][0] ),
    .B2(_05727_),
    .X(_03541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12768_ (.A1(_05503_),
    .A2(_07368_),
    .B1(_07364_),
    .B2(_05638_),
    .X(_05739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12769_ (.A(_05739_),
    .Y(_05740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12770_ (.A(_05740_),
    .X(_05741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12771_ (.A(_05739_),
    .X(_05742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12772_ (.A1(_00276_),
    .A2(_05741_),
    .B1(\design_top.MEM[20][7] ),
    .B2(_05742_),
    .X(_03540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12773_ (.A1(_00275_),
    .A2(_05741_),
    .B1(\design_top.MEM[20][6] ),
    .B2(_05742_),
    .X(_03539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12774_ (.A1(_00274_),
    .A2(_05741_),
    .B1(\design_top.MEM[20][5] ),
    .B2(_05742_),
    .X(_03538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12775_ (.A1(_00273_),
    .A2(_05741_),
    .B1(\design_top.MEM[20][4] ),
    .B2(_05742_),
    .X(_03537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12776_ (.A1(_00272_),
    .A2(_05741_),
    .B1(\design_top.MEM[20][3] ),
    .B2(_05742_),
    .X(_03536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12777_ (.A1(_00271_),
    .A2(_05740_),
    .B1(\design_top.MEM[20][2] ),
    .B2(_05739_),
    .X(_03535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12778_ (.A1(_00270_),
    .A2(_05740_),
    .B1(\design_top.MEM[20][1] ),
    .B2(_05739_),
    .X(_03534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12779_ (.A1(_00269_),
    .A2(_05740_),
    .B1(\design_top.MEM[20][0] ),
    .B2(_05739_),
    .X(_03533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12780_ (.A1(_05521_),
    .A2(_07367_),
    .B1(_07381_),
    .B2(_05638_),
    .X(_05743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12781_ (.A(_05743_),
    .Y(_05744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12782_ (.A(_05744_),
    .X(_05745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12783_ (.A(_05743_),
    .X(_05746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12784_ (.A1(_00284_),
    .A2(_05745_),
    .B1(\design_top.MEM[21][7] ),
    .B2(_05746_),
    .X(_03532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12785_ (.A1(_00283_),
    .A2(_05745_),
    .B1(\design_top.MEM[21][6] ),
    .B2(_05746_),
    .X(_03531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12786_ (.A1(_00282_),
    .A2(_05745_),
    .B1(\design_top.MEM[21][5] ),
    .B2(_05746_),
    .X(_03530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12787_ (.A1(_00281_),
    .A2(_05745_),
    .B1(\design_top.MEM[21][4] ),
    .B2(_05746_),
    .X(_03529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12788_ (.A1(_00280_),
    .A2(_05745_),
    .B1(\design_top.MEM[21][3] ),
    .B2(_05746_),
    .X(_03528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12789_ (.A1(_00279_),
    .A2(_05744_),
    .B1(\design_top.MEM[21][2] ),
    .B2(_05743_),
    .X(_03527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12790_ (.A1(_00278_),
    .A2(_05744_),
    .B1(\design_top.MEM[21][1] ),
    .B2(_05743_),
    .X(_03526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12791_ (.A1(_00277_),
    .A2(_05744_),
    .B1(\design_top.MEM[21][0] ),
    .B2(_05743_),
    .X(_03525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12792_ (.A1(_08021_),
    .A2(_07367_),
    .B1(_07404_),
    .B2(_05638_),
    .X(_05747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12793_ (.A(_05747_),
    .Y(_05748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12794_ (.A(_05748_),
    .X(_05749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12795_ (.A(_05747_),
    .X(_05750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12796_ (.A1(_00292_),
    .A2(_05749_),
    .B1(\design_top.MEM[22][7] ),
    .B2(_05750_),
    .X(_03524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12797_ (.A1(_00291_),
    .A2(_05749_),
    .B1(\design_top.MEM[22][6] ),
    .B2(_05750_),
    .X(_03523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12798_ (.A1(_00290_),
    .A2(_05749_),
    .B1(\design_top.MEM[22][5] ),
    .B2(_05750_),
    .X(_03522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12799_ (.A1(_00289_),
    .A2(_05749_),
    .B1(\design_top.MEM[22][4] ),
    .B2(_05750_),
    .X(_03521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12800_ (.A1(_00288_),
    .A2(_05749_),
    .B1(\design_top.MEM[22][3] ),
    .B2(_05750_),
    .X(_03520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12801_ (.A1(_00287_),
    .A2(_05748_),
    .B1(\design_top.MEM[22][2] ),
    .B2(_05747_),
    .X(_03519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12802_ (.A1(_00286_),
    .A2(_05748_),
    .B1(\design_top.MEM[22][1] ),
    .B2(_05747_),
    .X(_03518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12803_ (.A1(_00285_),
    .A2(_05748_),
    .B1(\design_top.MEM[22][0] ),
    .B2(_05747_),
    .X(_03517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12804_ (.A(_08407_),
    .X(_05751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12805_ (.A(_05751_),
    .X(_05752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12806_ (.A(\design_top.core0.REG2[0][31] ),
    .B(_05752_),
    .X(_03516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12807_ (.A(\design_top.core0.REG2[0][30] ),
    .B(_05752_),
    .X(_03515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12808_ (.A(\design_top.core0.REG2[0][29] ),
    .B(_05752_),
    .X(_03514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12809_ (.A(\design_top.core0.REG2[0][28] ),
    .B(_05752_),
    .X(_03513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12810_ (.A(\design_top.core0.REG2[0][27] ),
    .B(_05752_),
    .X(_03512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12811_ (.A(_05751_),
    .X(_05753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12812_ (.A(\design_top.core0.REG2[0][26] ),
    .B(_05753_),
    .X(_03511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12813_ (.A(\design_top.core0.REG2[0][25] ),
    .B(_05753_),
    .X(_03510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12814_ (.A(\design_top.core0.REG2[0][24] ),
    .B(_05753_),
    .X(_03509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12815_ (.A(\design_top.core0.REG2[0][23] ),
    .B(_05753_),
    .X(_03508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12816_ (.A(\design_top.core0.REG2[0][22] ),
    .B(_05753_),
    .X(_03507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12817_ (.A(_05751_),
    .X(_05754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12818_ (.A(\design_top.core0.REG2[0][21] ),
    .B(_05754_),
    .X(_03506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12819_ (.A(\design_top.core0.REG2[0][20] ),
    .B(_05754_),
    .X(_03505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12820_ (.A(\design_top.core0.REG2[0][19] ),
    .B(_05754_),
    .X(_03504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12821_ (.A(\design_top.core0.REG2[0][18] ),
    .B(_05754_),
    .X(_03503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12822_ (.A(\design_top.core0.REG2[0][17] ),
    .B(_05754_),
    .X(_03502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12823_ (.A(_08407_),
    .X(_05755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12824_ (.A(\design_top.core0.REG2[0][16] ),
    .B(_05755_),
    .X(_03501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12825_ (.A(\design_top.core0.REG2[0][15] ),
    .B(_05755_),
    .X(_03500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12826_ (.A(\design_top.core0.REG2[0][14] ),
    .B(_05755_),
    .X(_03499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12827_ (.A1(\design_top.core0.REG2[0][13] ),
    .A2(_05751_),
    .B1(_05655_),
    .B2(_08076_),
    .X(_03498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12828_ (.A(\design_top.core0.REG2[0][12] ),
    .B(_05755_),
    .X(_03497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12829_ (.A(\design_top.core0.REG2[0][11] ),
    .B(_05755_),
    .X(_03496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12830_ (.A(_08407_),
    .X(_05756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12831_ (.A(\design_top.core0.REG2[0][10] ),
    .B(_05756_),
    .X(_03495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12832_ (.A(\design_top.core0.REG2[0][9] ),
    .B(_05756_),
    .X(_03494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12833_ (.A(\design_top.core0.REG2[0][8] ),
    .B(_05756_),
    .X(_03493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12834_ (.A(\design_top.core0.REG2[0][7] ),
    .B(_05756_),
    .X(_03492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12835_ (.A(\design_top.core0.REG2[0][6] ),
    .B(_05756_),
    .X(_03491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12836_ (.A(_08407_),
    .X(_05757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12837_ (.A(\design_top.core0.REG2[0][5] ),
    .B(_05757_),
    .X(_03490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12838_ (.A(\design_top.core0.REG2[0][4] ),
    .B(_05757_),
    .X(_03489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12839_ (.A(\design_top.core0.REG2[0][3] ),
    .B(_05757_),
    .X(_03488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12840_ (.A(\design_top.core0.REG2[0][2] ),
    .B(_05757_),
    .X(_03487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12841_ (.A(\design_top.core0.REG2[0][1] ),
    .B(_05757_),
    .X(_03486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _12842_ (.A(\design_top.core0.REG2[0][0] ),
    .B(_05751_),
    .X(_03485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12843_ (.A(_08418_),
    .X(_05758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12844_ (.A(_05758_),
    .X(_05759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12845_ (.A(_05759_),
    .X(_05760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12846_ (.A(_05758_),
    .Y(_05761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12847_ (.A(_05761_),
    .X(_05762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12848_ (.A(_05762_),
    .X(_05763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12849_ (.A1(_05676_),
    .A2(_05760_),
    .B1(\design_top.core0.REG2[10][31] ),
    .B2(_05763_),
    .X(_03484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12850_ (.A1(_05683_),
    .A2(_05760_),
    .B1(\design_top.core0.REG2[10][30] ),
    .B2(_05763_),
    .X(_03483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12851_ (.A1(_05684_),
    .A2(_05760_),
    .B1(\design_top.core0.REG2[10][29] ),
    .B2(_05763_),
    .X(_03482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12852_ (.A1(_05685_),
    .A2(_05760_),
    .B1(\design_top.core0.REG2[10][28] ),
    .B2(_05763_),
    .X(_03481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12853_ (.A1(_05686_),
    .A2(_05760_),
    .B1(\design_top.core0.REG2[10][27] ),
    .B2(_05763_),
    .X(_03480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12854_ (.A(_05759_),
    .X(_05764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12855_ (.A(_05762_),
    .X(_05765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12856_ (.A1(_05687_),
    .A2(_05764_),
    .B1(\design_top.core0.REG2[10][26] ),
    .B2(_05765_),
    .X(_03479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12857_ (.A1(_05690_),
    .A2(_05764_),
    .B1(\design_top.core0.REG2[10][25] ),
    .B2(_05765_),
    .X(_03478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12858_ (.A1(_05691_),
    .A2(_05764_),
    .B1(\design_top.core0.REG2[10][24] ),
    .B2(_05765_),
    .X(_03477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12859_ (.A1(_05692_),
    .A2(_05764_),
    .B1(\design_top.core0.REG2[10][23] ),
    .B2(_05765_),
    .X(_03476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12860_ (.A1(_05693_),
    .A2(_05764_),
    .B1(\design_top.core0.REG2[10][22] ),
    .B2(_05765_),
    .X(_03475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12861_ (.A(_05759_),
    .X(_05766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12862_ (.A(_05762_),
    .X(_05767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12863_ (.A1(_05694_),
    .A2(_05766_),
    .B1(\design_top.core0.REG2[10][21] ),
    .B2(_05767_),
    .X(_03474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12864_ (.A1(_05697_),
    .A2(_05766_),
    .B1(\design_top.core0.REG2[10][20] ),
    .B2(_05767_),
    .X(_03473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12865_ (.A1(_05698_),
    .A2(_05766_),
    .B1(\design_top.core0.REG2[10][19] ),
    .B2(_05767_),
    .X(_03472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12866_ (.A1(_05699_),
    .A2(_05766_),
    .B1(\design_top.core0.REG2[10][18] ),
    .B2(_05767_),
    .X(_03471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12867_ (.A1(_05700_),
    .A2(_05766_),
    .B1(\design_top.core0.REG2[10][17] ),
    .B2(_05767_),
    .X(_03470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12868_ (.A(_05758_),
    .X(_05768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12869_ (.A(_05761_),
    .X(_05769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12870_ (.A1(_05701_),
    .A2(_05768_),
    .B1(\design_top.core0.REG2[10][16] ),
    .B2(_05769_),
    .X(_03469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12871_ (.A1(_05704_),
    .A2(_05768_),
    .B1(\design_top.core0.REG2[10][15] ),
    .B2(_05769_),
    .X(_03468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12872_ (.A1(_05705_),
    .A2(_05768_),
    .B1(\design_top.core0.REG2[10][14] ),
    .B2(_05769_),
    .X(_03467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12873_ (.A(_08531_),
    .X(_05770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12874_ (.A1(\design_top.core0.REG2[10][13] ),
    .A2(_05759_),
    .B1(_05770_),
    .B2(_05762_),
    .X(_03466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12875_ (.A1(_05706_),
    .A2(_05768_),
    .B1(\design_top.core0.REG2[10][12] ),
    .B2(_05769_),
    .X(_03465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12876_ (.A1(_05707_),
    .A2(_05768_),
    .B1(\design_top.core0.REG2[10][11] ),
    .B2(_05769_),
    .X(_03464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12877_ (.A(_05758_),
    .X(_05771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12878_ (.A(_05761_),
    .X(_05772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12879_ (.A1(_05708_),
    .A2(_05771_),
    .B1(\design_top.core0.REG2[10][10] ),
    .B2(_05772_),
    .X(_03463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12880_ (.A1(_05711_),
    .A2(_05771_),
    .B1(\design_top.core0.REG2[10][9] ),
    .B2(_05772_),
    .X(_03462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12881_ (.A1(_05712_),
    .A2(_05771_),
    .B1(\design_top.core0.REG2[10][8] ),
    .B2(_05772_),
    .X(_03461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12882_ (.A1(_05713_),
    .A2(_05771_),
    .B1(\design_top.core0.REG2[10][7] ),
    .B2(_05772_),
    .X(_03460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12883_ (.A1(_05714_),
    .A2(_05771_),
    .B1(\design_top.core0.REG2[10][6] ),
    .B2(_05772_),
    .X(_03459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12884_ (.A(_05758_),
    .X(_05773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12885_ (.A(_05761_),
    .X(_05774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12886_ (.A1(_05715_),
    .A2(_05773_),
    .B1(\design_top.core0.REG2[10][5] ),
    .B2(_05774_),
    .X(_03458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12887_ (.A1(_05718_),
    .A2(_05773_),
    .B1(\design_top.core0.REG2[10][4] ),
    .B2(_05774_),
    .X(_03457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12888_ (.A1(_05719_),
    .A2(_05773_),
    .B1(\design_top.core0.REG2[10][3] ),
    .B2(_05774_),
    .X(_03456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12889_ (.A1(_05720_),
    .A2(_05773_),
    .B1(\design_top.core0.REG2[10][2] ),
    .B2(_05774_),
    .X(_03455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12890_ (.A1(_05721_),
    .A2(_05773_),
    .B1(\design_top.core0.REG2[10][1] ),
    .B2(_05774_),
    .X(_03454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12891_ (.A1(_05722_),
    .A2(_05759_),
    .B1(\design_top.core0.REG2[10][0] ),
    .B2(_05762_),
    .X(_03453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12892_ (.A(_08436_),
    .X(_05775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12893_ (.A(_05775_),
    .X(_05776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12894_ (.A(_05776_),
    .X(_05777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12895_ (.A(_05775_),
    .Y(_05778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12896_ (.A(_05778_),
    .X(_05779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12897_ (.A(_05779_),
    .X(_05780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12898_ (.A1(_05676_),
    .A2(_05777_),
    .B1(\design_top.core0.REG2[11][31] ),
    .B2(_05780_),
    .X(_03452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12899_ (.A1(_05683_),
    .A2(_05777_),
    .B1(\design_top.core0.REG2[11][30] ),
    .B2(_05780_),
    .X(_03451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12900_ (.A1(_05684_),
    .A2(_05777_),
    .B1(\design_top.core0.REG2[11][29] ),
    .B2(_05780_),
    .X(_03450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12901_ (.A1(_05685_),
    .A2(_05777_),
    .B1(\design_top.core0.REG2[11][28] ),
    .B2(_05780_),
    .X(_03449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12902_ (.A1(_05686_),
    .A2(_05777_),
    .B1(\design_top.core0.REG2[11][27] ),
    .B2(_05780_),
    .X(_03448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12903_ (.A(_05776_),
    .X(_05781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12904_ (.A(_05779_),
    .X(_05782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12905_ (.A1(_05687_),
    .A2(_05781_),
    .B1(\design_top.core0.REG2[11][26] ),
    .B2(_05782_),
    .X(_03447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12906_ (.A1(_05690_),
    .A2(_05781_),
    .B1(\design_top.core0.REG2[11][25] ),
    .B2(_05782_),
    .X(_03446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12907_ (.A1(_05691_),
    .A2(_05781_),
    .B1(\design_top.core0.REG2[11][24] ),
    .B2(_05782_),
    .X(_03445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12908_ (.A1(_05692_),
    .A2(_05781_),
    .B1(\design_top.core0.REG2[11][23] ),
    .B2(_05782_),
    .X(_03444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12909_ (.A1(_05693_),
    .A2(_05781_),
    .B1(\design_top.core0.REG2[11][22] ),
    .B2(_05782_),
    .X(_03443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12910_ (.A(_05776_),
    .X(_05783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12911_ (.A(_05779_),
    .X(_05784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12912_ (.A1(_05694_),
    .A2(_05783_),
    .B1(\design_top.core0.REG2[11][21] ),
    .B2(_05784_),
    .X(_03442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12913_ (.A1(_05697_),
    .A2(_05783_),
    .B1(\design_top.core0.REG2[11][20] ),
    .B2(_05784_),
    .X(_03441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12914_ (.A1(_05698_),
    .A2(_05783_),
    .B1(\design_top.core0.REG2[11][19] ),
    .B2(_05784_),
    .X(_03440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12915_ (.A1(_05699_),
    .A2(_05783_),
    .B1(\design_top.core0.REG2[11][18] ),
    .B2(_05784_),
    .X(_03439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12916_ (.A1(_05700_),
    .A2(_05783_),
    .B1(\design_top.core0.REG2[11][17] ),
    .B2(_05784_),
    .X(_03438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12917_ (.A(_05775_),
    .X(_05785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12918_ (.A(_05778_),
    .X(_05786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12919_ (.A1(_05701_),
    .A2(_05785_),
    .B1(\design_top.core0.REG2[11][16] ),
    .B2(_05786_),
    .X(_03437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12920_ (.A1(_05704_),
    .A2(_05785_),
    .B1(\design_top.core0.REG2[11][15] ),
    .B2(_05786_),
    .X(_03436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12921_ (.A1(_05705_),
    .A2(_05785_),
    .B1(\design_top.core0.REG2[11][14] ),
    .B2(_05786_),
    .X(_03435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12922_ (.A1(\design_top.core0.REG2[11][13] ),
    .A2(_05776_),
    .B1(_05770_),
    .B2(_05779_),
    .X(_03434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12923_ (.A1(_05706_),
    .A2(_05785_),
    .B1(\design_top.core0.REG2[11][12] ),
    .B2(_05786_),
    .X(_03433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12924_ (.A1(_05707_),
    .A2(_05785_),
    .B1(\design_top.core0.REG2[11][11] ),
    .B2(_05786_),
    .X(_03432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12925_ (.A(_05775_),
    .X(_05787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12926_ (.A(_05778_),
    .X(_05788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12927_ (.A1(_05708_),
    .A2(_05787_),
    .B1(\design_top.core0.REG2[11][10] ),
    .B2(_05788_),
    .X(_03431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12928_ (.A1(_05711_),
    .A2(_05787_),
    .B1(\design_top.core0.REG2[11][9] ),
    .B2(_05788_),
    .X(_03430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12929_ (.A1(_05712_),
    .A2(_05787_),
    .B1(\design_top.core0.REG2[11][8] ),
    .B2(_05788_),
    .X(_03429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12930_ (.A1(_05713_),
    .A2(_05787_),
    .B1(\design_top.core0.REG2[11][7] ),
    .B2(_05788_),
    .X(_03428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12931_ (.A1(_05714_),
    .A2(_05787_),
    .B1(\design_top.core0.REG2[11][6] ),
    .B2(_05788_),
    .X(_03427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12932_ (.A(_05775_),
    .X(_05789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12933_ (.A(_05778_),
    .X(_05790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12934_ (.A1(_05715_),
    .A2(_05789_),
    .B1(\design_top.core0.REG2[11][5] ),
    .B2(_05790_),
    .X(_03426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12935_ (.A1(_05718_),
    .A2(_05789_),
    .B1(\design_top.core0.REG2[11][4] ),
    .B2(_05790_),
    .X(_03425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12936_ (.A1(_05719_),
    .A2(_05789_),
    .B1(\design_top.core0.REG2[11][3] ),
    .B2(_05790_),
    .X(_03424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12937_ (.A1(_05720_),
    .A2(_05789_),
    .B1(\design_top.core0.REG2[11][2] ),
    .B2(_05790_),
    .X(_03423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12938_ (.A1(_05721_),
    .A2(_05789_),
    .B1(\design_top.core0.REG2[11][1] ),
    .B2(_05790_),
    .X(_03422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12939_ (.A1(_05722_),
    .A2(_05776_),
    .B1(\design_top.core0.REG2[11][0] ),
    .B2(_05779_),
    .X(_03421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12940_ (.A(_08453_),
    .X(_05791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12941_ (.A(_05791_),
    .X(_05792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12942_ (.A(_05792_),
    .X(_05793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12943_ (.A(_05791_),
    .Y(_05794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12944_ (.A(_05794_),
    .X(_05795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12945_ (.A(_05795_),
    .X(_05796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12946_ (.A1(_05676_),
    .A2(_05793_),
    .B1(\design_top.core0.REG2[12][31] ),
    .B2(_05796_),
    .X(_03420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12947_ (.A1(_05683_),
    .A2(_05793_),
    .B1(\design_top.core0.REG2[12][30] ),
    .B2(_05796_),
    .X(_03419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12948_ (.A1(_05684_),
    .A2(_05793_),
    .B1(\design_top.core0.REG2[12][29] ),
    .B2(_05796_),
    .X(_03418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12949_ (.A1(_05685_),
    .A2(_05793_),
    .B1(\design_top.core0.REG2[12][28] ),
    .B2(_05796_),
    .X(_03417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12950_ (.A1(_05686_),
    .A2(_05793_),
    .B1(\design_top.core0.REG2[12][27] ),
    .B2(_05796_),
    .X(_03416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12951_ (.A(_05792_),
    .X(_05797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12952_ (.A(_05795_),
    .X(_05798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12953_ (.A1(_05687_),
    .A2(_05797_),
    .B1(\design_top.core0.REG2[12][26] ),
    .B2(_05798_),
    .X(_03415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12954_ (.A1(_05690_),
    .A2(_05797_),
    .B1(\design_top.core0.REG2[12][25] ),
    .B2(_05798_),
    .X(_03414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12955_ (.A1(_05691_),
    .A2(_05797_),
    .B1(\design_top.core0.REG2[12][24] ),
    .B2(_05798_),
    .X(_03413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12956_ (.A1(_05692_),
    .A2(_05797_),
    .B1(\design_top.core0.REG2[12][23] ),
    .B2(_05798_),
    .X(_03412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12957_ (.A1(_05693_),
    .A2(_05797_),
    .B1(\design_top.core0.REG2[12][22] ),
    .B2(_05798_),
    .X(_03411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12958_ (.A(_05792_),
    .X(_05799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12959_ (.A(_05795_),
    .X(_05800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12960_ (.A1(_05694_),
    .A2(_05799_),
    .B1(\design_top.core0.REG2[12][21] ),
    .B2(_05800_),
    .X(_03410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12961_ (.A1(_05697_),
    .A2(_05799_),
    .B1(\design_top.core0.REG2[12][20] ),
    .B2(_05800_),
    .X(_03409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12962_ (.A1(_05698_),
    .A2(_05799_),
    .B1(\design_top.core0.REG2[12][19] ),
    .B2(_05800_),
    .X(_03408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12963_ (.A1(_05699_),
    .A2(_05799_),
    .B1(\design_top.core0.REG2[12][18] ),
    .B2(_05800_),
    .X(_03407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12964_ (.A1(_05700_),
    .A2(_05799_),
    .B1(\design_top.core0.REG2[12][17] ),
    .B2(_05800_),
    .X(_03406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12965_ (.A(_05791_),
    .X(_05801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12966_ (.A(_05794_),
    .X(_05802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12967_ (.A1(_05701_),
    .A2(_05801_),
    .B1(\design_top.core0.REG2[12][16] ),
    .B2(_05802_),
    .X(_03405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12968_ (.A1(_05704_),
    .A2(_05801_),
    .B1(\design_top.core0.REG2[12][15] ),
    .B2(_05802_),
    .X(_03404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12969_ (.A1(_05705_),
    .A2(_05801_),
    .B1(\design_top.core0.REG2[12][14] ),
    .B2(_05802_),
    .X(_03403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _12970_ (.A1(\design_top.core0.REG2[12][13] ),
    .A2(_05792_),
    .B1(_05770_),
    .B2(_05795_),
    .X(_03402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12971_ (.A1(_05706_),
    .A2(_05801_),
    .B1(\design_top.core0.REG2[12][12] ),
    .B2(_05802_),
    .X(_03401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12972_ (.A1(_05707_),
    .A2(_05801_),
    .B1(\design_top.core0.REG2[12][11] ),
    .B2(_05802_),
    .X(_03400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12973_ (.A(_05791_),
    .X(_05803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12974_ (.A(_05794_),
    .X(_05804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12975_ (.A1(_05708_),
    .A2(_05803_),
    .B1(\design_top.core0.REG2[12][10] ),
    .B2(_05804_),
    .X(_03399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12976_ (.A1(_05711_),
    .A2(_05803_),
    .B1(\design_top.core0.REG2[12][9] ),
    .B2(_05804_),
    .X(_03398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12977_ (.A1(_05712_),
    .A2(_05803_),
    .B1(\design_top.core0.REG2[12][8] ),
    .B2(_05804_),
    .X(_03397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12978_ (.A1(_05713_),
    .A2(_05803_),
    .B1(\design_top.core0.REG2[12][7] ),
    .B2(_05804_),
    .X(_03396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12979_ (.A1(_05714_),
    .A2(_05803_),
    .B1(\design_top.core0.REG2[12][6] ),
    .B2(_05804_),
    .X(_03395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12980_ (.A(_05791_),
    .X(_05805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12981_ (.A(_05794_),
    .X(_05806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12982_ (.A1(_05715_),
    .A2(_05805_),
    .B1(\design_top.core0.REG2[12][5] ),
    .B2(_05806_),
    .X(_03394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12983_ (.A1(_05718_),
    .A2(_05805_),
    .B1(\design_top.core0.REG2[12][4] ),
    .B2(_05806_),
    .X(_03393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12984_ (.A1(_05719_),
    .A2(_05805_),
    .B1(\design_top.core0.REG2[12][3] ),
    .B2(_05806_),
    .X(_03392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12985_ (.A1(_05720_),
    .A2(_05805_),
    .B1(\design_top.core0.REG2[12][2] ),
    .B2(_05806_),
    .X(_03391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12986_ (.A1(_05721_),
    .A2(_05805_),
    .B1(\design_top.core0.REG2[12][1] ),
    .B2(_05806_),
    .X(_03390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12987_ (.A1(_05722_),
    .A2(_05792_),
    .B1(\design_top.core0.REG2[12][0] ),
    .B2(_05795_),
    .X(_03389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12988_ (.A(_08501_),
    .X(_05807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12989_ (.A(_05807_),
    .X(_05808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12990_ (.A(_05808_),
    .X(_05809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _12991_ (.A(_05807_),
    .Y(_05810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12992_ (.A(_05810_),
    .X(_05811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12993_ (.A(_05811_),
    .X(_05812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12994_ (.A1(_08089_),
    .A2(_05809_),
    .B1(\design_top.core0.REG2[13][31] ),
    .B2(_05812_),
    .X(_03388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12995_ (.A1(_08091_),
    .A2(_05809_),
    .B1(\design_top.core0.REG2[13][30] ),
    .B2(_05812_),
    .X(_03387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12996_ (.A1(_08093_),
    .A2(_05809_),
    .B1(\design_top.core0.REG2[13][29] ),
    .B2(_05812_),
    .X(_03386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12997_ (.A1(_08095_),
    .A2(_05809_),
    .B1(\design_top.core0.REG2[13][28] ),
    .B2(_05812_),
    .X(_03385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _12998_ (.A1(_08098_),
    .A2(_05809_),
    .B1(\design_top.core0.REG2[13][27] ),
    .B2(_05812_),
    .X(_03384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _12999_ (.A(_05808_),
    .X(_05813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13000_ (.A(_05811_),
    .X(_05814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13001_ (.A1(_08102_),
    .A2(_05813_),
    .B1(\design_top.core0.REG2[13][26] ),
    .B2(_05814_),
    .X(_03383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13002_ (.A1(_08104_),
    .A2(_05813_),
    .B1(\design_top.core0.REG2[13][25] ),
    .B2(_05814_),
    .X(_03382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13003_ (.A1(_08106_),
    .A2(_05813_),
    .B1(\design_top.core0.REG2[13][24] ),
    .B2(_05814_),
    .X(_03381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13004_ (.A1(_08108_),
    .A2(_05813_),
    .B1(\design_top.core0.REG2[13][23] ),
    .B2(_05814_),
    .X(_03380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13005_ (.A1(_08111_),
    .A2(_05813_),
    .B1(\design_top.core0.REG2[13][22] ),
    .B2(_05814_),
    .X(_03379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13006_ (.A(_05808_),
    .X(_05815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13007_ (.A(_05811_),
    .X(_05816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13008_ (.A1(_08115_),
    .A2(_05815_),
    .B1(\design_top.core0.REG2[13][21] ),
    .B2(_05816_),
    .X(_03378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13009_ (.A1(_08117_),
    .A2(_05815_),
    .B1(\design_top.core0.REG2[13][20] ),
    .B2(_05816_),
    .X(_03377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13010_ (.A1(_08119_),
    .A2(_05815_),
    .B1(\design_top.core0.REG2[13][19] ),
    .B2(_05816_),
    .X(_03376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13011_ (.A1(_08121_),
    .A2(_05815_),
    .B1(\design_top.core0.REG2[13][18] ),
    .B2(_05816_),
    .X(_03375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13012_ (.A1(_08124_),
    .A2(_05815_),
    .B1(\design_top.core0.REG2[13][17] ),
    .B2(_05816_),
    .X(_03374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13013_ (.A(_05807_),
    .X(_05817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13014_ (.A(_05810_),
    .X(_05818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13015_ (.A1(_08128_),
    .A2(_05817_),
    .B1(\design_top.core0.REG2[13][16] ),
    .B2(_05818_),
    .X(_03373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13016_ (.A1(_08130_),
    .A2(_05817_),
    .B1(\design_top.core0.REG2[13][15] ),
    .B2(_05818_),
    .X(_03372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13017_ (.A1(_08132_),
    .A2(_05817_),
    .B1(\design_top.core0.REG2[13][14] ),
    .B2(_05818_),
    .X(_03371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13018_ (.A1(\design_top.core0.REG2[13][13] ),
    .A2(_05808_),
    .B1(_05770_),
    .B2(_05811_),
    .X(_03370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13019_ (.A1(_08135_),
    .A2(_05817_),
    .B1(\design_top.core0.REG2[13][12] ),
    .B2(_05818_),
    .X(_03369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13020_ (.A1(_08138_),
    .A2(_05817_),
    .B1(\design_top.core0.REG2[13][11] ),
    .B2(_05818_),
    .X(_03368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13021_ (.A(_05807_),
    .X(_05819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13022_ (.A(_05810_),
    .X(_05820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13023_ (.A1(_08142_),
    .A2(_05819_),
    .B1(\design_top.core0.REG2[13][10] ),
    .B2(_05820_),
    .X(_03367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13024_ (.A1(_08144_),
    .A2(_05819_),
    .B1(\design_top.core0.REG2[13][9] ),
    .B2(_05820_),
    .X(_03366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13025_ (.A1(_08146_),
    .A2(_05819_),
    .B1(\design_top.core0.REG2[13][8] ),
    .B2(_05820_),
    .X(_03365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13026_ (.A1(_08148_),
    .A2(_05819_),
    .B1(\design_top.core0.REG2[13][7] ),
    .B2(_05820_),
    .X(_03364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13027_ (.A1(_08151_),
    .A2(_05819_),
    .B1(\design_top.core0.REG2[13][6] ),
    .B2(_05820_),
    .X(_03363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13028_ (.A(_05807_),
    .X(_05821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13029_ (.A(_05810_),
    .X(_05822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13030_ (.A1(_08155_),
    .A2(_05821_),
    .B1(\design_top.core0.REG2[13][5] ),
    .B2(_05822_),
    .X(_03362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13031_ (.A1(_08157_),
    .A2(_05821_),
    .B1(\design_top.core0.REG2[13][4] ),
    .B2(_05822_),
    .X(_03361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13032_ (.A1(_08159_),
    .A2(_05821_),
    .B1(\design_top.core0.REG2[13][3] ),
    .B2(_05822_),
    .X(_03360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13033_ (.A1(_08161_),
    .A2(_05821_),
    .B1(\design_top.core0.REG2[13][2] ),
    .B2(_05822_),
    .X(_03359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13034_ (.A1(_08163_),
    .A2(_05821_),
    .B1(\design_top.core0.REG2[13][1] ),
    .B2(_05822_),
    .X(_03358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13035_ (.A1(_08165_),
    .A2(_05808_),
    .B1(\design_top.core0.REG2[13][0] ),
    .B2(_05811_),
    .X(_03357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13036_ (.A(_08518_),
    .X(_05823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13037_ (.A(_05823_),
    .X(_05824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13038_ (.A(_05824_),
    .X(_05825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13039_ (.A(_05823_),
    .Y(_05826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13040_ (.A(_05826_),
    .X(_05827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13041_ (.A(_05827_),
    .X(_05828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13042_ (.A1(_08089_),
    .A2(_05825_),
    .B1(\design_top.core0.REG2[14][31] ),
    .B2(_05828_),
    .X(_03356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13043_ (.A1(_08091_),
    .A2(_05825_),
    .B1(\design_top.core0.REG2[14][30] ),
    .B2(_05828_),
    .X(_03355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13044_ (.A1(_08093_),
    .A2(_05825_),
    .B1(\design_top.core0.REG2[14][29] ),
    .B2(_05828_),
    .X(_03354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13045_ (.A1(_08095_),
    .A2(_05825_),
    .B1(\design_top.core0.REG2[14][28] ),
    .B2(_05828_),
    .X(_03353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13046_ (.A1(_08098_),
    .A2(_05825_),
    .B1(\design_top.core0.REG2[14][27] ),
    .B2(_05828_),
    .X(_03352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13047_ (.A(_05824_),
    .X(_05829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13048_ (.A(_05827_),
    .X(_05830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13049_ (.A1(_08102_),
    .A2(_05829_),
    .B1(\design_top.core0.REG2[14][26] ),
    .B2(_05830_),
    .X(_03351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13050_ (.A1(_08104_),
    .A2(_05829_),
    .B1(\design_top.core0.REG2[14][25] ),
    .B2(_05830_),
    .X(_03350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13051_ (.A1(_08106_),
    .A2(_05829_),
    .B1(\design_top.core0.REG2[14][24] ),
    .B2(_05830_),
    .X(_03349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13052_ (.A1(_08108_),
    .A2(_05829_),
    .B1(\design_top.core0.REG2[14][23] ),
    .B2(_05830_),
    .X(_03348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13053_ (.A1(_08111_),
    .A2(_05829_),
    .B1(\design_top.core0.REG2[14][22] ),
    .B2(_05830_),
    .X(_03347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13054_ (.A(_05824_),
    .X(_05831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13055_ (.A(_05827_),
    .X(_05832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13056_ (.A1(_08115_),
    .A2(_05831_),
    .B1(\design_top.core0.REG2[14][21] ),
    .B2(_05832_),
    .X(_03346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13057_ (.A1(_08117_),
    .A2(_05831_),
    .B1(\design_top.core0.REG2[14][20] ),
    .B2(_05832_),
    .X(_03345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13058_ (.A1(_08119_),
    .A2(_05831_),
    .B1(\design_top.core0.REG2[14][19] ),
    .B2(_05832_),
    .X(_03344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13059_ (.A1(_08121_),
    .A2(_05831_),
    .B1(\design_top.core0.REG2[14][18] ),
    .B2(_05832_),
    .X(_03343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13060_ (.A1(_08124_),
    .A2(_05831_),
    .B1(\design_top.core0.REG2[14][17] ),
    .B2(_05832_),
    .X(_03342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13061_ (.A(_05823_),
    .X(_05833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13062_ (.A(_05826_),
    .X(_05834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13063_ (.A1(_08128_),
    .A2(_05833_),
    .B1(\design_top.core0.REG2[14][16] ),
    .B2(_05834_),
    .X(_03341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13064_ (.A1(_08130_),
    .A2(_05833_),
    .B1(\design_top.core0.REG2[14][15] ),
    .B2(_05834_),
    .X(_03340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13065_ (.A1(_08132_),
    .A2(_05833_),
    .B1(\design_top.core0.REG2[14][14] ),
    .B2(_05834_),
    .X(_03339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13066_ (.A1(\design_top.core0.REG2[14][13] ),
    .A2(_05824_),
    .B1(_05770_),
    .B2(_05827_),
    .X(_03338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13067_ (.A1(_08135_),
    .A2(_05833_),
    .B1(\design_top.core0.REG2[14][12] ),
    .B2(_05834_),
    .X(_03337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13068_ (.A1(_08138_),
    .A2(_05833_),
    .B1(\design_top.core0.REG2[14][11] ),
    .B2(_05834_),
    .X(_03336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13069_ (.A(_05823_),
    .X(_05835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13070_ (.A(_05826_),
    .X(_05836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13071_ (.A1(_08142_),
    .A2(_05835_),
    .B1(\design_top.core0.REG2[14][10] ),
    .B2(_05836_),
    .X(_03335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13072_ (.A1(_08144_),
    .A2(_05835_),
    .B1(\design_top.core0.REG2[14][9] ),
    .B2(_05836_),
    .X(_03334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13073_ (.A1(_08146_),
    .A2(_05835_),
    .B1(\design_top.core0.REG2[14][8] ),
    .B2(_05836_),
    .X(_03333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13074_ (.A1(_08148_),
    .A2(_05835_),
    .B1(\design_top.core0.REG2[14][7] ),
    .B2(_05836_),
    .X(_03332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13075_ (.A1(_08151_),
    .A2(_05835_),
    .B1(\design_top.core0.REG2[14][6] ),
    .B2(_05836_),
    .X(_03331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13076_ (.A(_05823_),
    .X(_05837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13077_ (.A(_05826_),
    .X(_05838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13078_ (.A1(_08155_),
    .A2(_05837_),
    .B1(\design_top.core0.REG2[14][5] ),
    .B2(_05838_),
    .X(_03330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13079_ (.A1(_08157_),
    .A2(_05837_),
    .B1(\design_top.core0.REG2[14][4] ),
    .B2(_05838_),
    .X(_03329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13080_ (.A1(_08159_),
    .A2(_05837_),
    .B1(\design_top.core0.REG2[14][3] ),
    .B2(_05838_),
    .X(_03328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13081_ (.A1(_08161_),
    .A2(_05837_),
    .B1(\design_top.core0.REG2[14][2] ),
    .B2(_05838_),
    .X(_03327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13082_ (.A1(_08163_),
    .A2(_05837_),
    .B1(\design_top.core0.REG2[14][1] ),
    .B2(_05838_),
    .X(_03326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13083_ (.A1(_08165_),
    .A2(_05824_),
    .B1(\design_top.core0.REG2[14][0] ),
    .B2(_05827_),
    .X(_03325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13084_ (.A1(_06868_),
    .A2(_06900_),
    .B1(_07414_),
    .B2(_05638_),
    .X(_05839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13085_ (.A(_05839_),
    .Y(_05840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13086_ (.A(_05840_),
    .X(_05841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13087_ (.A(_05839_),
    .X(_05842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13088_ (.A1(_00420_),
    .A2(_05841_),
    .B1(\design_top.MEM[8][7] ),
    .B2(_05842_),
    .X(_03324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13089_ (.A1(_00419_),
    .A2(_05841_),
    .B1(\design_top.MEM[8][6] ),
    .B2(_05842_),
    .X(_03323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13090_ (.A1(_00418_),
    .A2(_05841_),
    .B1(\design_top.MEM[8][5] ),
    .B2(_05842_),
    .X(_03322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13091_ (.A1(_00417_),
    .A2(_05841_),
    .B1(\design_top.MEM[8][4] ),
    .B2(_05842_),
    .X(_03321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13092_ (.A1(_00416_),
    .A2(_05841_),
    .B1(\design_top.MEM[8][3] ),
    .B2(_05842_),
    .X(_03320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13093_ (.A1(_00415_),
    .A2(_05840_),
    .B1(\design_top.MEM[8][2] ),
    .B2(_05839_),
    .X(_03319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13094_ (.A1(_00414_),
    .A2(_05840_),
    .B1(\design_top.MEM[8][1] ),
    .B2(_05839_),
    .X(_03318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13095_ (.A1(_00413_),
    .A2(_05840_),
    .B1(\design_top.MEM[8][0] ),
    .B2(_05839_),
    .X(_03317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13096_ (.A(_08015_),
    .X(_05843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13097_ (.A1(_05521_),
    .A2(_06868_),
    .B1(_06858_),
    .B2(_05843_),
    .X(_05844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13098_ (.A(_05844_),
    .Y(_05845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13099_ (.A(_05845_),
    .X(_05846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13100_ (.A(_05844_),
    .X(_05847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13101_ (.A1(_00428_),
    .A2(_05846_),
    .B1(\design_top.MEM[9][7] ),
    .B2(_05847_),
    .X(_03316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13102_ (.A1(_00427_),
    .A2(_05846_),
    .B1(\design_top.MEM[9][6] ),
    .B2(_05847_),
    .X(_03315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13103_ (.A1(_00426_),
    .A2(_05846_),
    .B1(\design_top.MEM[9][5] ),
    .B2(_05847_),
    .X(_03314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13104_ (.A1(_00425_),
    .A2(_05846_),
    .B1(\design_top.MEM[9][4] ),
    .B2(_05847_),
    .X(_03313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13105_ (.A1(_00424_),
    .A2(_05846_),
    .B1(\design_top.MEM[9][3] ),
    .B2(_05847_),
    .X(_03312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13106_ (.A1(_00423_),
    .A2(_05845_),
    .B1(\design_top.MEM[9][2] ),
    .B2(_05844_),
    .X(_03311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13107_ (.A1(_00422_),
    .A2(_05845_),
    .B1(\design_top.MEM[9][1] ),
    .B2(_05844_),
    .X(_03310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13108_ (.A1(_00421_),
    .A2(_05845_),
    .B1(\design_top.MEM[9][0] ),
    .B2(_05844_),
    .X(_03309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13109_ (.A1(_05503_),
    .A2(_07463_),
    .B1(_07459_),
    .B2(_05843_),
    .X(_05848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13110_ (.A(_05848_),
    .Y(_05849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13111_ (.A(_05849_),
    .X(_05850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13112_ (.A(_05848_),
    .X(_05851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13113_ (.A1(_00308_),
    .A2(_05850_),
    .B1(\design_top.MEM[24][7] ),
    .B2(_05851_),
    .X(_03308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13114_ (.A1(_00307_),
    .A2(_05850_),
    .B1(\design_top.MEM[24][6] ),
    .B2(_05851_),
    .X(_03307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13115_ (.A1(_00306_),
    .A2(_05850_),
    .B1(\design_top.MEM[24][5] ),
    .B2(_05851_),
    .X(_03306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13116_ (.A1(_00305_),
    .A2(_05850_),
    .B1(\design_top.MEM[24][4] ),
    .B2(_05851_),
    .X(_03305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13117_ (.A1(_00304_),
    .A2(_05850_),
    .B1(\design_top.MEM[24][3] ),
    .B2(_05851_),
    .X(_03304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13118_ (.A1(_00303_),
    .A2(_05849_),
    .B1(\design_top.MEM[24][2] ),
    .B2(_05848_),
    .X(_03303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13119_ (.A1(_00302_),
    .A2(_05849_),
    .B1(\design_top.MEM[24][1] ),
    .B2(_05848_),
    .X(_03302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13120_ (.A1(_00301_),
    .A2(_05849_),
    .B1(\design_top.MEM[24][0] ),
    .B2(_05848_),
    .X(_03301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13121_ (.A1(_05521_),
    .A2(_07462_),
    .B1(_07479_),
    .B2(_05843_),
    .X(_05852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13122_ (.A(_05852_),
    .Y(_05853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13123_ (.A(_05853_),
    .X(_05854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13124_ (.A(_05852_),
    .X(_05855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13125_ (.A1(_00316_),
    .A2(_05854_),
    .B1(\design_top.MEM[25][7] ),
    .B2(_05855_),
    .X(_03300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13126_ (.A1(_00315_),
    .A2(_05854_),
    .B1(\design_top.MEM[25][6] ),
    .B2(_05855_),
    .X(_03299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13127_ (.A1(_00314_),
    .A2(_05854_),
    .B1(\design_top.MEM[25][5] ),
    .B2(_05855_),
    .X(_03298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13128_ (.A1(_00313_),
    .A2(_05854_),
    .B1(\design_top.MEM[25][4] ),
    .B2(_05855_),
    .X(_03297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13129_ (.A1(_00312_),
    .A2(_05854_),
    .B1(\design_top.MEM[25][3] ),
    .B2(_05855_),
    .X(_03296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13130_ (.A1(_00311_),
    .A2(_05853_),
    .B1(\design_top.MEM[25][2] ),
    .B2(_05852_),
    .X(_03295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13131_ (.A1(_00310_),
    .A2(_05853_),
    .B1(\design_top.MEM[25][1] ),
    .B2(_05852_),
    .X(_03294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13132_ (.A1(_00309_),
    .A2(_05853_),
    .B1(\design_top.MEM[25][0] ),
    .B2(_05852_),
    .X(_03293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13133_ (.A1(_08021_),
    .A2(_07462_),
    .B1(_07493_),
    .B2(_05843_),
    .X(_05856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13134_ (.A(_05856_),
    .Y(_05857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13135_ (.A(_05857_),
    .X(_05858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13136_ (.A(_05856_),
    .X(_05859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13137_ (.A1(_00324_),
    .A2(_05858_),
    .B1(\design_top.MEM[26][7] ),
    .B2(_05859_),
    .X(_03292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13138_ (.A1(_00323_),
    .A2(_05858_),
    .B1(\design_top.MEM[26][6] ),
    .B2(_05859_),
    .X(_03291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13139_ (.A1(_00322_),
    .A2(_05858_),
    .B1(\design_top.MEM[26][5] ),
    .B2(_05859_),
    .X(_03290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13140_ (.A1(_00321_),
    .A2(_05858_),
    .B1(\design_top.MEM[26][4] ),
    .B2(_05859_),
    .X(_03289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13141_ (.A1(_00320_),
    .A2(_05858_),
    .B1(\design_top.MEM[26][3] ),
    .B2(_05859_),
    .X(_03288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13142_ (.A1(_00319_),
    .A2(_05857_),
    .B1(\design_top.MEM[26][2] ),
    .B2(_05856_),
    .X(_03287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13143_ (.A1(_00318_),
    .A2(_05857_),
    .B1(\design_top.MEM[26][1] ),
    .B2(_05856_),
    .X(_03286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13144_ (.A1(_00317_),
    .A2(_05857_),
    .B1(\design_top.MEM[26][0] ),
    .B2(_05856_),
    .X(_03285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13145_ (.A1(_08045_),
    .A2(_07462_),
    .B1(_07534_),
    .B2(_05843_),
    .X(_05860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13146_ (.A(_05860_),
    .Y(_05861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13147_ (.A(_05861_),
    .X(_05862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13148_ (.A(_05860_),
    .X(_05863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13149_ (.A1(_00332_),
    .A2(_05862_),
    .B1(\design_top.MEM[27][7] ),
    .B2(_05863_),
    .X(_03284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13150_ (.A1(_00331_),
    .A2(_05862_),
    .B1(\design_top.MEM[27][6] ),
    .B2(_05863_),
    .X(_03283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13151_ (.A1(_00330_),
    .A2(_05862_),
    .B1(\design_top.MEM[27][5] ),
    .B2(_05863_),
    .X(_03282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13152_ (.A1(_00329_),
    .A2(_05862_),
    .B1(\design_top.MEM[27][4] ),
    .B2(_05863_),
    .X(_03281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13153_ (.A1(_00328_),
    .A2(_05862_),
    .B1(\design_top.MEM[27][3] ),
    .B2(_05863_),
    .X(_03280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13154_ (.A1(_00327_),
    .A2(_05861_),
    .B1(\design_top.MEM[27][2] ),
    .B2(_05860_),
    .X(_03279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13155_ (.A1(_00326_),
    .A2(_05861_),
    .B1(\design_top.MEM[27][1] ),
    .B2(_05860_),
    .X(_03278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13156_ (.A1(_00325_),
    .A2(_05861_),
    .B1(\design_top.MEM[27][0] ),
    .B2(_05860_),
    .X(_03277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13157_ (.A(_08015_),
    .X(_05864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13158_ (.A1(_08045_),
    .A2(_07367_),
    .B1(_07437_),
    .B2(_05864_),
    .X(_05865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13159_ (.A(_05865_),
    .Y(_05866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13160_ (.A(_05866_),
    .X(_05867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13161_ (.A(_05865_),
    .X(_05868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13162_ (.A1(_00300_),
    .A2(_05867_),
    .B1(\design_top.MEM[23][7] ),
    .B2(_05868_),
    .X(_03276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13163_ (.A1(_00299_),
    .A2(_05867_),
    .B1(\design_top.MEM[23][6] ),
    .B2(_05868_),
    .X(_03275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13164_ (.A1(_00298_),
    .A2(_05867_),
    .B1(\design_top.MEM[23][5] ),
    .B2(_05868_),
    .X(_03274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13165_ (.A1(_00297_),
    .A2(_05867_),
    .B1(\design_top.MEM[23][4] ),
    .B2(_05868_),
    .X(_03273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13166_ (.A1(_00296_),
    .A2(_05867_),
    .B1(\design_top.MEM[23][3] ),
    .B2(_05868_),
    .X(_03272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13167_ (.A1(_00295_),
    .A2(_05866_),
    .B1(\design_top.MEM[23][2] ),
    .B2(_05865_),
    .X(_03271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13168_ (.A1(_00294_),
    .A2(_05866_),
    .B1(\design_top.MEM[23][1] ),
    .B2(_05865_),
    .X(_03270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13169_ (.A1(_00293_),
    .A2(_05866_),
    .B1(\design_top.MEM[23][0] ),
    .B2(_05865_),
    .X(_03269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13170_ (.A1(_05503_),
    .A2(_07066_),
    .B1(_07554_),
    .B2(_05864_),
    .X(_05869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13171_ (.A(_05869_),
    .Y(_05870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13172_ (.A(_05870_),
    .X(_05871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13173_ (.A(_05869_),
    .X(_05872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13174_ (.A1(_00340_),
    .A2(_05871_),
    .B1(\design_top.MEM[28][7] ),
    .B2(_05872_),
    .X(_03268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13175_ (.A1(_00339_),
    .A2(_05871_),
    .B1(\design_top.MEM[28][6] ),
    .B2(_05872_),
    .X(_03267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13176_ (.A1(_00338_),
    .A2(_05871_),
    .B1(\design_top.MEM[28][5] ),
    .B2(_05872_),
    .X(_03266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13177_ (.A1(_00337_),
    .A2(_05871_),
    .B1(\design_top.MEM[28][4] ),
    .B2(_05872_),
    .X(_03265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13178_ (.A1(_00336_),
    .A2(_05871_),
    .B1(\design_top.MEM[28][3] ),
    .B2(_05872_),
    .X(_03264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13179_ (.A1(_00335_),
    .A2(_05870_),
    .B1(\design_top.MEM[28][2] ),
    .B2(_05869_),
    .X(_03263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13180_ (.A1(_00334_),
    .A2(_05870_),
    .B1(\design_top.MEM[28][1] ),
    .B2(_05869_),
    .X(_03262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13181_ (.A1(_00333_),
    .A2(_05870_),
    .B1(\design_top.MEM[28][0] ),
    .B2(_05869_),
    .X(_03261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13182_ (.A1(_05521_),
    .A2(_07066_),
    .B1(_07568_),
    .B2(_05864_),
    .X(_05873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13183_ (.A(_05873_),
    .Y(_05874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13184_ (.A(_05874_),
    .X(_05875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13185_ (.A(_05873_),
    .X(_05876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13186_ (.A1(_00348_),
    .A2(_05875_),
    .B1(\design_top.MEM[29][7] ),
    .B2(_05876_),
    .X(_03260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13187_ (.A1(_00347_),
    .A2(_05875_),
    .B1(\design_top.MEM[29][6] ),
    .B2(_05876_),
    .X(_03259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13188_ (.A1(_00346_),
    .A2(_05875_),
    .B1(\design_top.MEM[29][5] ),
    .B2(_05876_),
    .X(_03258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13189_ (.A1(_00345_),
    .A2(_05875_),
    .B1(\design_top.MEM[29][4] ),
    .B2(_05876_),
    .X(_03257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13190_ (.A1(_00344_),
    .A2(_05875_),
    .B1(\design_top.MEM[29][3] ),
    .B2(_05876_),
    .X(_03256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13191_ (.A1(_00343_),
    .A2(_05874_),
    .B1(\design_top.MEM[29][2] ),
    .B2(_05873_),
    .X(_03255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13192_ (.A1(_00342_),
    .A2(_05874_),
    .B1(\design_top.MEM[29][1] ),
    .B2(_05873_),
    .X(_03254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13193_ (.A1(_00341_),
    .A2(_05874_),
    .B1(\design_top.MEM[29][0] ),
    .B2(_05873_),
    .X(_03253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13194_ (.A1(_06903_),
    .A2(_06976_),
    .B1(_07052_),
    .B2(_05864_),
    .X(_05877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13195_ (.A(_05877_),
    .Y(_05878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13196_ (.A(_05878_),
    .X(_05879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13197_ (.A(_05877_),
    .X(_05880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13198_ (.A1(_00356_),
    .A2(_05879_),
    .B1(\design_top.MEM[2][7] ),
    .B2(_05880_),
    .X(_03252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13199_ (.A1(_00355_),
    .A2(_05879_),
    .B1(\design_top.MEM[2][6] ),
    .B2(_05880_),
    .X(_03251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13200_ (.A1(_00354_),
    .A2(_05879_),
    .B1(\design_top.MEM[2][5] ),
    .B2(_05880_),
    .X(_03250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13201_ (.A1(_00353_),
    .A2(_05879_),
    .B1(\design_top.MEM[2][4] ),
    .B2(_05880_),
    .X(_03249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13202_ (.A1(_00352_),
    .A2(_05879_),
    .B1(\design_top.MEM[2][3] ),
    .B2(_05880_),
    .X(_03248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13203_ (.A1(_00351_),
    .A2(_05878_),
    .B1(\design_top.MEM[2][2] ),
    .B2(_05877_),
    .X(_03247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13204_ (.A1(_00350_),
    .A2(_05878_),
    .B1(\design_top.MEM[2][1] ),
    .B2(_05877_),
    .X(_03246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13205_ (.A1(_00349_),
    .A2(_05878_),
    .B1(\design_top.MEM[2][0] ),
    .B2(_05877_),
    .X(_03245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13206_ (.A1(_06864_),
    .A2(_07182_),
    .B1(_07179_),
    .B2(_05864_),
    .X(_05881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13207_ (.A(_05881_),
    .Y(_05882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13208_ (.A(_05882_),
    .X(_05883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13209_ (.A(_05881_),
    .X(_05884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13210_ (.A1(_00212_),
    .A2(_05883_),
    .B1(\design_top.MEM[13][7] ),
    .B2(_05884_),
    .X(_03244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13211_ (.A1(_00211_),
    .A2(_05883_),
    .B1(\design_top.MEM[13][6] ),
    .B2(_05884_),
    .X(_03243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13212_ (.A1(_00210_),
    .A2(_05883_),
    .B1(\design_top.MEM[13][5] ),
    .B2(_05884_),
    .X(_03242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13213_ (.A1(_00209_),
    .A2(_05883_),
    .B1(\design_top.MEM[13][4] ),
    .B2(_05884_),
    .X(_03241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13214_ (.A1(_00208_),
    .A2(_05883_),
    .B1(\design_top.MEM[13][3] ),
    .B2(_05884_),
    .X(_03240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13215_ (.A1(_00207_),
    .A2(_05882_),
    .B1(\design_top.MEM[13][2] ),
    .B2(_05881_),
    .X(_03239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13216_ (.A1(_00206_),
    .A2(_05882_),
    .B1(\design_top.MEM[13][1] ),
    .B2(_05881_),
    .X(_03238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13217_ (.A1(_00205_),
    .A2(_05882_),
    .B1(\design_top.MEM[13][0] ),
    .B2(_05881_),
    .X(_03237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13218_ (.A(_07601_),
    .Y(_05885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13219_ (.A(_06982_),
    .B(_05885_),
    .X(_05886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13220_ (.A(_06970_),
    .B(_06987_),
    .X(_05887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13221_ (.A(_05886_),
    .B(_05887_),
    .X(_05888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13222_ (.A(_05888_),
    .X(_05889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13223_ (.A(_05888_),
    .Y(_05890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13224_ (.A(_05890_),
    .X(_05891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13225_ (.A1(\design_top.GPIOFF[15] ),
    .A2(_05889_),
    .B1(\design_top.DATAO[31] ),
    .B2(_05891_),
    .X(_03236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13226_ (.A1(\design_top.GPIOFF[14] ),
    .A2(_05889_),
    .B1(\design_top.DATAO[30] ),
    .B2(_05891_),
    .X(_03235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13227_ (.A1(\design_top.GPIOFF[13] ),
    .A2(_05889_),
    .B1(\design_top.DATAO[29] ),
    .B2(_05891_),
    .X(_03234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13228_ (.A1(\design_top.GPIOFF[12] ),
    .A2(_05889_),
    .B1(\design_top.DATAO[28] ),
    .B2(_05891_),
    .X(_03233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13229_ (.A1(\design_top.GPIOFF[11] ),
    .A2(_05889_),
    .B1(\design_top.DATAO[27] ),
    .B2(_05891_),
    .X(_03232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13230_ (.A(_05888_),
    .X(_05892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13231_ (.A(_05890_),
    .X(_05893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13232_ (.A1(\design_top.GPIOFF[10] ),
    .A2(_05892_),
    .B1(\design_top.DATAO[26] ),
    .B2(_05893_),
    .X(_03231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13233_ (.A1(\design_top.GPIOFF[9] ),
    .A2(_05892_),
    .B1(\design_top.DATAO[25] ),
    .B2(_05893_),
    .X(_03230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13234_ (.A1(\design_top.GPIOFF[8] ),
    .A2(_05892_),
    .B1(\design_top.DATAO[24] ),
    .B2(_05893_),
    .X(_03229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13235_ (.A1(\design_top.GPIOFF[7] ),
    .A2(_05892_),
    .B1(\design_top.DATAO[23] ),
    .B2(_05893_),
    .X(_03228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13236_ (.A1(\design_top.GPIOFF[6] ),
    .A2(_05892_),
    .B1(\design_top.DATAO[22] ),
    .B2(_05893_),
    .X(_03227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13237_ (.A(_05888_),
    .X(_05894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13238_ (.A(_05890_),
    .X(_05895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13239_ (.A1(\design_top.GPIOFF[5] ),
    .A2(_05894_),
    .B1(\design_top.DATAO[21] ),
    .B2(_05895_),
    .X(_03226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13240_ (.A1(\design_top.GPIOFF[4] ),
    .A2(_05894_),
    .B1(\design_top.DATAO[20] ),
    .B2(_05895_),
    .X(_03225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13241_ (.A1(\design_top.GPIOFF[3] ),
    .A2(_05894_),
    .B1(\design_top.DATAO[19] ),
    .B2(_05895_),
    .X(_03224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13242_ (.A1(\design_top.GPIOFF[2] ),
    .A2(_05894_),
    .B1(\design_top.DATAO[18] ),
    .B2(_05895_),
    .X(_03223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13243_ (.A1(\design_top.GPIOFF[1] ),
    .A2(_05894_),
    .B1(\design_top.DATAO[17] ),
    .B2(_05895_),
    .X(_03222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13244_ (.A1(io_out[15]),
    .A2(_05888_),
    .B1(\design_top.DATAO[16] ),
    .B2(_05890_),
    .X(_03221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13245_ (.A(_01381_),
    .B(_05887_),
    .X(_05896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13246_ (.A(_05896_),
    .X(_05897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13247_ (.A(_05896_),
    .Y(_05898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13248_ (.A(_05898_),
    .X(_05899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13249_ (.A1(\design_top.LEDFF[15] ),
    .A2(_05897_),
    .B1(\design_top.DATAO[15] ),
    .B2(_05899_),
    .X(_03220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13250_ (.A1(\design_top.LEDFF[14] ),
    .A2(_05897_),
    .B1(\design_top.DATAO[14] ),
    .B2(_05899_),
    .X(_03219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13251_ (.A1(\design_top.LEDFF[13] ),
    .A2(_05897_),
    .B1(\design_top.DATAO[13] ),
    .B2(_05899_),
    .X(_03218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13252_ (.A1(\design_top.LEDFF[12] ),
    .A2(_05897_),
    .B1(\design_top.DATAO[12] ),
    .B2(_05899_),
    .X(_03217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13253_ (.A1(\design_top.LEDFF[11] ),
    .A2(_05897_),
    .B1(\design_top.DATAO[11] ),
    .B2(_05899_),
    .X(_03216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13254_ (.A(_05896_),
    .X(_05900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13255_ (.A(_05898_),
    .X(_05901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13256_ (.A1(\design_top.LEDFF[10] ),
    .A2(_05900_),
    .B1(\design_top.DATAO[10] ),
    .B2(_05901_),
    .X(_03215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13257_ (.A1(\design_top.LEDFF[9] ),
    .A2(_05900_),
    .B1(\design_top.DATAO[9] ),
    .B2(_05901_),
    .X(_03214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13258_ (.A1(\design_top.LEDFF[8] ),
    .A2(_05900_),
    .B1(\design_top.DATAO[8] ),
    .B2(_05901_),
    .X(_03213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13259_ (.A1(\design_top.LEDFF[7] ),
    .A2(_05900_),
    .B1(\design_top.DATAO[7] ),
    .B2(_05901_),
    .X(_03212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13260_ (.A1(\design_top.LEDFF[6] ),
    .A2(_05900_),
    .B1(\design_top.DATAO[6] ),
    .B2(_05901_),
    .X(_03211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13261_ (.A(_05896_),
    .X(_05902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13262_ (.A(_05898_),
    .X(_05903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13263_ (.A1(\design_top.LEDFF[5] ),
    .A2(_05902_),
    .B1(\design_top.DATAO[5] ),
    .B2(_05903_),
    .X(_03210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13264_ (.A1(\design_top.LEDFF[4] ),
    .A2(_05902_),
    .B1(\design_top.DATAO[4] ),
    .B2(_05903_),
    .X(_03209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13265_ (.A1(io_out[11]),
    .A2(_05902_),
    .B1(\design_top.DATAO[3] ),
    .B2(_05903_),
    .X(_03208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13266_ (.A1(io_out[10]),
    .A2(_05902_),
    .B1(\design_top.DATAO[2] ),
    .B2(_05903_),
    .X(_03207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13267_ (.A1(io_out[9]),
    .A2(_05902_),
    .B1(\design_top.DATAO[1] ),
    .B2(_05903_),
    .X(_03206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13268_ (.A1(io_out[8]),
    .A2(_05896_),
    .B1(\design_top.DATAO[0] ),
    .B2(_05898_),
    .X(_03205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13269_ (.A1(\design_top.ROMFF2[31] ),
    .A2(_07804_),
    .B1(\design_top.ROMFF[31] ),
    .B2(\design_top.HLT ),
    .X(_03204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13270_ (.A1(\design_top.ROMFF2[30] ),
    .A2(_07804_),
    .B1(\design_top.ROMFF[30] ),
    .B2(\design_top.HLT ),
    .X(_03203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13271_ (.A1(\design_top.ROMFF2[29] ),
    .A2(_07804_),
    .B1(\design_top.ROMFF[29] ),
    .B2(\design_top.HLT ),
    .X(_03202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13272_ (.A(_07751_),
    .X(_05904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13273_ (.A1(\design_top.ROMFF2[28] ),
    .A2(_07804_),
    .B1(\design_top.ROMFF[28] ),
    .B2(_05904_),
    .X(_03201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13274_ (.A(_07756_),
    .X(_05905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13275_ (.A1(\design_top.ROMFF2[27] ),
    .A2(_05905_),
    .B1(\design_top.ROMFF[27] ),
    .B2(_05904_),
    .X(_03200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13276_ (.A1(\design_top.ROMFF2[26] ),
    .A2(_05905_),
    .B1(\design_top.ROMFF[26] ),
    .B2(_05904_),
    .X(_03199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13277_ (.A1(\design_top.ROMFF2[25] ),
    .A2(_05905_),
    .B1(\design_top.ROMFF[25] ),
    .B2(_05904_),
    .X(_03198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13278_ (.A1(\design_top.ROMFF2[24] ),
    .A2(_05905_),
    .B1(\design_top.ROMFF[24] ),
    .B2(_05904_),
    .X(_03197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13279_ (.A(_07659_),
    .X(_05906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13280_ (.A(_05906_),
    .X(_05907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13281_ (.A1(\design_top.ROMFF2[23] ),
    .A2(_05905_),
    .B1(\design_top.ROMFF[23] ),
    .B2(_05907_),
    .X(_03196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13282_ (.A(_07726_),
    .X(_05908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13283_ (.A(_05908_),
    .X(_05909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13284_ (.A1(\design_top.ROMFF2[22] ),
    .A2(_05909_),
    .B1(\design_top.ROMFF[22] ),
    .B2(_05907_),
    .X(_03195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13285_ (.A1(\design_top.ROMFF2[21] ),
    .A2(_05909_),
    .B1(\design_top.ROMFF[21] ),
    .B2(_05907_),
    .X(_03194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13286_ (.A1(\design_top.ROMFF2[20] ),
    .A2(_05909_),
    .B1(\design_top.ROMFF[20] ),
    .B2(_05907_),
    .X(_03193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13287_ (.A1(\design_top.ROMFF2[19] ),
    .A2(_05909_),
    .B1(\design_top.ROMFF[19] ),
    .B2(_05907_),
    .X(_03192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13288_ (.A(_05906_),
    .X(_05910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13289_ (.A1(\design_top.ROMFF2[18] ),
    .A2(_05909_),
    .B1(\design_top.ROMFF[18] ),
    .B2(_05910_),
    .X(_03191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13290_ (.A(_05908_),
    .X(_05911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13291_ (.A1(\design_top.ROMFF2[17] ),
    .A2(_05911_),
    .B1(\design_top.ROMFF[17] ),
    .B2(_05910_),
    .X(_03190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13292_ (.A1(\design_top.ROMFF2[16] ),
    .A2(_05911_),
    .B1(\design_top.ROMFF[16] ),
    .B2(_05910_),
    .X(_03189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13293_ (.A1(\design_top.ROMFF2[15] ),
    .A2(_05911_),
    .B1(\design_top.ROMFF[15] ),
    .B2(_05910_),
    .X(_03188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13294_ (.A1(\design_top.ROMFF2[14] ),
    .A2(_05911_),
    .B1(\design_top.ROMFF[14] ),
    .B2(_05910_),
    .X(_03187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13295_ (.A(_05906_),
    .X(_05912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13296_ (.A1(\design_top.ROMFF2[13] ),
    .A2(_05911_),
    .B1(\design_top.ROMFF[13] ),
    .B2(_05912_),
    .X(_03186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13297_ (.A(_05908_),
    .X(_05913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13298_ (.A1(\design_top.ROMFF2[12] ),
    .A2(_05913_),
    .B1(\design_top.ROMFF[12] ),
    .B2(_05912_),
    .X(_03185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13299_ (.A1(\design_top.ROMFF2[11] ),
    .A2(_05913_),
    .B1(\design_top.ROMFF[11] ),
    .B2(_05912_),
    .X(_03184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13300_ (.A1(\design_top.ROMFF2[10] ),
    .A2(_05913_),
    .B1(\design_top.ROMFF[10] ),
    .B2(_05912_),
    .X(_03183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13301_ (.A1(\design_top.ROMFF2[9] ),
    .A2(_05913_),
    .B1(\design_top.ROMFF[9] ),
    .B2(_05912_),
    .X(_03182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13302_ (.A(_05906_),
    .X(_05914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13303_ (.A1(\design_top.ROMFF2[8] ),
    .A2(_05913_),
    .B1(\design_top.ROMFF[8] ),
    .B2(_05914_),
    .X(_03181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13304_ (.A(_05908_),
    .X(_05915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13305_ (.A1(\design_top.ROMFF2[7] ),
    .A2(_05915_),
    .B1(\design_top.ROMFF[7] ),
    .B2(_05914_),
    .X(_03180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13306_ (.A1(\design_top.ROMFF2[6] ),
    .A2(_05915_),
    .B1(\design_top.ROMFF[6] ),
    .B2(_05914_),
    .X(_03179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13307_ (.A1(\design_top.ROMFF2[5] ),
    .A2(_05915_),
    .B1(\design_top.ROMFF[5] ),
    .B2(_05914_),
    .X(_03178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13308_ (.A1(\design_top.ROMFF2[4] ),
    .A2(_05915_),
    .B1(\design_top.ROMFF[4] ),
    .B2(_05914_),
    .X(_03177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13309_ (.A(_05906_),
    .X(_05916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13310_ (.A1(\design_top.ROMFF2[3] ),
    .A2(_05915_),
    .B1(\design_top.ROMFF[3] ),
    .B2(_05916_),
    .X(_03176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13311_ (.A(_05908_),
    .X(_05917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13312_ (.A1(\design_top.ROMFF2[2] ),
    .A2(_05917_),
    .B1(\design_top.ROMFF[2] ),
    .B2(_05916_),
    .X(_03175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13313_ (.A1(\design_top.ROMFF2[1] ),
    .A2(_05917_),
    .B1(\design_top.ROMFF[1] ),
    .B2(_05916_),
    .X(_03174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13314_ (.A1(\design_top.ROMFF2[0] ),
    .A2(_05917_),
    .B1(\design_top.ROMFF[0] ),
    .B2(_05916_),
    .X(_03173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13315_ (.A1(\design_top.uart0.UART_XREQ ),
    .A2(_07952_),
    .B1(\design_top.uart0.UART_XACK ),
    .B2(_07960_),
    .X(_03172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13316_ (.A(\design_top.uart0.UART_RACK ),
    .Y(_05918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _13317_ (.A0(_05918_),
    .A1(\design_top.uart0.UART_RREQ ),
    .S(_07968_),
    .X(_03171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13318_ (.A(\design_top.uart0.UART_RXDFF[2] ),
    .X(_05919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _13319_ (.A(_07976_),
    .B(_07975_),
    .C(_07966_),
    .D(_07962_),
    .X(_05920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _13320_ (.A0(_05919_),
    .A1(\design_top.uart0.UART_RFIFO[7] ),
    .S(_05920_),
    .X(_03170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _13321_ (.A(_07976_),
    .B(_07978_),
    .C(_07966_),
    .D(_07899_),
    .X(_05921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _13322_ (.A0(_05919_),
    .A1(\design_top.uart0.UART_RFIFO[6] ),
    .S(_05921_),
    .X(_03169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13323_ (.A(_07965_),
    .X(_05922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _13324_ (.A(_07967_),
    .B(_07975_),
    .C(_05922_),
    .D(_07899_),
    .X(_05923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _13325_ (.A0(_05919_),
    .A1(\design_top.uart0.UART_RFIFO[5] ),
    .S(_05923_),
    .X(_03168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _13326_ (.A(_07966_),
    .B(_07962_),
    .C(_07967_),
    .D(_07978_),
    .X(_05924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _13327_ (.A0(_05919_),
    .A1(\design_top.uart0.UART_RFIFO[4] ),
    .S(_05924_),
    .X(_03167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _13328_ (.A(_07976_),
    .B(_07975_),
    .C(_05922_),
    .D(_07972_),
    .X(_05925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _13329_ (.A0(\design_top.uart0.UART_RXDFF[2] ),
    .A1(\design_top.uart0.UART_RFIFO[3] ),
    .S(_05925_),
    .X(_03166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _13330_ (.A(_07976_),
    .B(_07978_),
    .C(_05922_),
    .D(_07972_),
    .X(_05926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _13331_ (.A0(\design_top.uart0.UART_RXDFF[2] ),
    .A1(\design_top.uart0.UART_RFIFO[2] ),
    .S(_05926_),
    .X(_03165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _13332_ (.A(_07967_),
    .B(_07963_),
    .C(_05922_),
    .D(_07972_),
    .X(_05927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _13333_ (.A0(\design_top.uart0.UART_RXDFF[2] ),
    .A1(\design_top.uart0.UART_RFIFO[1] ),
    .S(_05927_),
    .X(_03164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _13334_ (.A(_07967_),
    .B(_07978_),
    .C(_05922_),
    .D(_07972_),
    .X(_05928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _13335_ (.A0(\design_top.uart0.UART_RXDFF[2] ),
    .A1(\design_top.uart0.UART_RFIFO[0] ),
    .S(_05928_),
    .X(_03163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13336_ (.A1(\design_top.core0.NXPC[31] ),
    .A2(_05917_),
    .B1(\design_top.core0.PC[31] ),
    .B2(_05916_),
    .X(_03162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13337_ (.A(_07659_),
    .X(_05929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13338_ (.A(_05929_),
    .X(_05930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13339_ (.A1(\design_top.core0.NXPC[30] ),
    .A2(_05917_),
    .B1(\design_top.core0.PC[30] ),
    .B2(_05930_),
    .X(_03161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13340_ (.A(_07726_),
    .X(_05931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13341_ (.A(_05931_),
    .X(_05932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13342_ (.A1(\design_top.core0.NXPC[29] ),
    .A2(_05932_),
    .B1(\design_top.core0.PC[29] ),
    .B2(_05930_),
    .X(_03160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13343_ (.A1(\design_top.core0.NXPC[28] ),
    .A2(_05932_),
    .B1(\design_top.core0.PC[28] ),
    .B2(_05930_),
    .X(_03159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13344_ (.A1(\design_top.core0.NXPC[27] ),
    .A2(_05932_),
    .B1(\design_top.core0.PC[27] ),
    .B2(_05930_),
    .X(_03158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13345_ (.A1(\design_top.core0.NXPC[26] ),
    .A2(_05932_),
    .B1(\design_top.core0.PC[26] ),
    .B2(_05930_),
    .X(_03157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13346_ (.A(_05929_),
    .X(_05933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13347_ (.A1(\design_top.core0.NXPC[25] ),
    .A2(_05932_),
    .B1(\design_top.core0.PC[25] ),
    .B2(_05933_),
    .X(_03156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13348_ (.A(_05931_),
    .X(_05934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13349_ (.A1(\design_top.core0.NXPC[24] ),
    .A2(_05934_),
    .B1(\design_top.core0.PC[24] ),
    .B2(_05933_),
    .X(_03155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13350_ (.A1(\design_top.core0.NXPC[23] ),
    .A2(_05934_),
    .B1(\design_top.core0.PC[23] ),
    .B2(_05933_),
    .X(_03154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13351_ (.A1(\design_top.core0.NXPC[22] ),
    .A2(_05934_),
    .B1(\design_top.core0.PC[22] ),
    .B2(_05933_),
    .X(_03153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13352_ (.A1(\design_top.core0.NXPC[21] ),
    .A2(_05934_),
    .B1(\design_top.core0.PC[21] ),
    .B2(_05933_),
    .X(_03152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13353_ (.A(_05929_),
    .X(_05935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13354_ (.A1(\design_top.core0.NXPC[20] ),
    .A2(_05934_),
    .B1(\design_top.core0.PC[20] ),
    .B2(_05935_),
    .X(_03151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13355_ (.A(_05931_),
    .X(_05936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13356_ (.A1(\design_top.core0.NXPC[19] ),
    .A2(_05936_),
    .B1(\design_top.core0.PC[19] ),
    .B2(_05935_),
    .X(_03150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13357_ (.A1(\design_top.core0.NXPC[18] ),
    .A2(_05936_),
    .B1(\design_top.core0.PC[18] ),
    .B2(_05935_),
    .X(_03149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13358_ (.A1(\design_top.core0.NXPC[17] ),
    .A2(_05936_),
    .B1(\design_top.core0.PC[17] ),
    .B2(_05935_),
    .X(_03148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13359_ (.A1(\design_top.core0.NXPC[16] ),
    .A2(_05936_),
    .B1(\design_top.core0.PC[16] ),
    .B2(_05935_),
    .X(_03147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13360_ (.A(_05929_),
    .X(_05937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13361_ (.A1(\design_top.core0.NXPC[15] ),
    .A2(_05936_),
    .B1(\design_top.core0.PC[15] ),
    .B2(_05937_),
    .X(_03146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13362_ (.A(_05931_),
    .X(_05938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13363_ (.A1(\design_top.core0.NXPC[14] ),
    .A2(_05938_),
    .B1(\design_top.core0.PC[14] ),
    .B2(_05937_),
    .X(_03145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13364_ (.A1(\design_top.core0.NXPC[13] ),
    .A2(_05938_),
    .B1(\design_top.core0.PC[13] ),
    .B2(_05937_),
    .X(_03144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13365_ (.A1(\design_top.core0.NXPC[12] ),
    .A2(_05938_),
    .B1(\design_top.core0.PC[12] ),
    .B2(_05937_),
    .X(_03143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13366_ (.A1(\design_top.core0.NXPC[11] ),
    .A2(_05938_),
    .B1(\design_top.core0.PC[11] ),
    .B2(_05937_),
    .X(_03142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13367_ (.A(_05929_),
    .X(_05939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13368_ (.A1(\design_top.core0.NXPC[10] ),
    .A2(_05938_),
    .B1(\design_top.core0.PC[10] ),
    .B2(_05939_),
    .X(_03141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13369_ (.A(_05931_),
    .X(_05940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13370_ (.A1(\design_top.core0.NXPC[9] ),
    .A2(_05940_),
    .B1(\design_top.core0.PC[9] ),
    .B2(_05939_),
    .X(_03140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13371_ (.A1(\design_top.core0.NXPC[8] ),
    .A2(_05940_),
    .B1(\design_top.core0.PC[8] ),
    .B2(_05939_),
    .X(_03139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13372_ (.A1(\design_top.core0.NXPC[7] ),
    .A2(_05940_),
    .B1(\design_top.core0.PC[7] ),
    .B2(_05939_),
    .X(_03138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13373_ (.A1(\design_top.core0.NXPC[6] ),
    .A2(_05940_),
    .B1(\design_top.core0.PC[6] ),
    .B2(_05939_),
    .X(_03137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13374_ (.A(_07659_),
    .X(_05941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13375_ (.A(_05941_),
    .X(_05942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13376_ (.A1(\design_top.core0.NXPC[5] ),
    .A2(_05940_),
    .B1(\design_top.core0.PC[5] ),
    .B2(_05942_),
    .X(_03136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13377_ (.A(_07726_),
    .X(_05943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13378_ (.A(_05943_),
    .X(_05944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13379_ (.A1(\design_top.core0.NXPC[4] ),
    .A2(_05944_),
    .B1(\design_top.core0.PC[4] ),
    .B2(_05942_),
    .X(_03135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13380_ (.A1(\design_top.core0.NXPC[3] ),
    .A2(_05944_),
    .B1(\design_top.core0.PC[3] ),
    .B2(_05942_),
    .X(_03134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13381_ (.A1(\design_top.core0.NXPC[2] ),
    .A2(_05944_),
    .B1(\design_top.core0.PC[2] ),
    .B2(_05942_),
    .X(_03133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13382_ (.A1(\design_top.core0.NXPC[1] ),
    .A2(_05944_),
    .B1(\design_top.core0.PC[1] ),
    .B2(_05942_),
    .X(_03132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13383_ (.A(_05941_),
    .X(_05945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13384_ (.A1(\design_top.core0.NXPC[0] ),
    .A2(_05944_),
    .B1(\design_top.core0.PC[0] ),
    .B2(_05945_),
    .X(_03131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13385_ (.A1(_05503_),
    .A2(_07182_),
    .B1(_07629_),
    .B2(_08022_),
    .X(_05946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13386_ (.A(_05946_),
    .Y(_05947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13387_ (.A(_05947_),
    .X(_05948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13388_ (.A(_05946_),
    .X(_05949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13389_ (.A1(_00204_),
    .A2(_05948_),
    .B1(\design_top.MEM[12][7] ),
    .B2(_05949_),
    .X(_03130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13390_ (.A1(_00203_),
    .A2(_05948_),
    .B1(\design_top.MEM[12][6] ),
    .B2(_05949_),
    .X(_03129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13391_ (.A1(_00202_),
    .A2(_05948_),
    .B1(\design_top.MEM[12][5] ),
    .B2(_05949_),
    .X(_03128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13392_ (.A1(_00201_),
    .A2(_05948_),
    .B1(\design_top.MEM[12][4] ),
    .B2(_05949_),
    .X(_03127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13393_ (.A1(_00200_),
    .A2(_05948_),
    .B1(\design_top.MEM[12][3] ),
    .B2(_05949_),
    .X(_03126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13394_ (.A1(_00199_),
    .A2(_05947_),
    .B1(\design_top.MEM[12][2] ),
    .B2(_05946_),
    .X(_03125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13395_ (.A1(_00198_),
    .A2(_05947_),
    .B1(\design_top.MEM[12][1] ),
    .B2(_05946_),
    .X(_03124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13396_ (.A1(_00197_),
    .A2(_05947_),
    .B1(\design_top.MEM[12][0] ),
    .B2(_05946_),
    .X(_03123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13397_ (.A(_05943_),
    .X(_05950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13398_ (.A1(\design_top.IADDR[31] ),
    .A2(_05950_),
    .B1(\design_top.core0.NXPC[31] ),
    .B2(_05945_),
    .X(_03122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13399_ (.A1(\design_top.IADDR[30] ),
    .A2(_05950_),
    .B1(\design_top.core0.NXPC[30] ),
    .B2(_05945_),
    .X(_03121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13400_ (.A1(\design_top.IADDR[29] ),
    .A2(_05950_),
    .B1(\design_top.core0.NXPC[29] ),
    .B2(_05945_),
    .X(_03120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13401_ (.A1(\design_top.IADDR[28] ),
    .A2(_05950_),
    .B1(\design_top.core0.NXPC[28] ),
    .B2(_05945_),
    .X(_03119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13402_ (.A(_05941_),
    .X(_05951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13403_ (.A1(\design_top.IADDR[27] ),
    .A2(_05950_),
    .B1(\design_top.core0.NXPC[27] ),
    .B2(_05951_),
    .X(_03118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13404_ (.A(_05943_),
    .X(_05952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13405_ (.A1(\design_top.IADDR[26] ),
    .A2(_05952_),
    .B1(\design_top.core0.NXPC[26] ),
    .B2(_05951_),
    .X(_03117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13406_ (.A1(\design_top.IADDR[25] ),
    .A2(_05952_),
    .B1(\design_top.core0.NXPC[25] ),
    .B2(_05951_),
    .X(_03116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13407_ (.A1(\design_top.IADDR[24] ),
    .A2(_05952_),
    .B1(\design_top.core0.NXPC[24] ),
    .B2(_05951_),
    .X(_03115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13408_ (.A1(\design_top.IADDR[23] ),
    .A2(_05952_),
    .B1(\design_top.core0.NXPC[23] ),
    .B2(_05951_),
    .X(_03114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13409_ (.A(_05941_),
    .X(_05953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13410_ (.A1(\design_top.IADDR[22] ),
    .A2(_05952_),
    .B1(\design_top.core0.NXPC[22] ),
    .B2(_05953_),
    .X(_03113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13411_ (.A(_05943_),
    .X(_05954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13412_ (.A1(\design_top.IADDR[21] ),
    .A2(_05954_),
    .B1(\design_top.core0.NXPC[21] ),
    .B2(_05953_),
    .X(_03112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13413_ (.A1(\design_top.IADDR[20] ),
    .A2(_05954_),
    .B1(\design_top.core0.NXPC[20] ),
    .B2(_05953_),
    .X(_03111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13414_ (.A1(\design_top.IADDR[19] ),
    .A2(_05954_),
    .B1(\design_top.core0.NXPC[19] ),
    .B2(_05953_),
    .X(_03110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13415_ (.A1(\design_top.IADDR[18] ),
    .A2(_05954_),
    .B1(\design_top.core0.NXPC[18] ),
    .B2(_05953_),
    .X(_03109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13416_ (.A(_05941_),
    .X(_05955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13417_ (.A1(\design_top.IADDR[17] ),
    .A2(_05954_),
    .B1(\design_top.core0.NXPC[17] ),
    .B2(_05955_),
    .X(_03108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13418_ (.A(_05943_),
    .X(_05956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13419_ (.A1(\design_top.IADDR[16] ),
    .A2(_05956_),
    .B1(\design_top.core0.NXPC[16] ),
    .B2(_05955_),
    .X(_03107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13420_ (.A1(\design_top.IADDR[15] ),
    .A2(_05956_),
    .B1(\design_top.core0.NXPC[15] ),
    .B2(_05955_),
    .X(_03106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13421_ (.A1(\design_top.IADDR[14] ),
    .A2(_05956_),
    .B1(\design_top.core0.NXPC[14] ),
    .B2(_05955_),
    .X(_03105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13422_ (.A1(\design_top.IADDR[13] ),
    .A2(_05956_),
    .B1(\design_top.core0.NXPC[13] ),
    .B2(_05955_),
    .X(_03104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13423_ (.A(_07642_),
    .X(_05957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13424_ (.A1(\design_top.IADDR[12] ),
    .A2(_05956_),
    .B1(\design_top.core0.NXPC[12] ),
    .B2(_05957_),
    .X(_03103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13425_ (.A(_07727_),
    .X(_05958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13426_ (.A1(\design_top.IADDR[11] ),
    .A2(_05958_),
    .B1(\design_top.core0.NXPC[11] ),
    .B2(_05957_),
    .X(_03102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13427_ (.A1(\design_top.IADDR[10] ),
    .A2(_05958_),
    .B1(\design_top.core0.NXPC[10] ),
    .B2(_05957_),
    .X(_03101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13428_ (.A1(\design_top.IADDR[9] ),
    .A2(_05958_),
    .B1(\design_top.core0.NXPC[9] ),
    .B2(_05957_),
    .X(_03100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13429_ (.A1(\design_top.IADDR[8] ),
    .A2(_05958_),
    .B1(\design_top.core0.NXPC[8] ),
    .B2(_05957_),
    .X(_03099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13430_ (.A(_07642_),
    .X(_05959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13431_ (.A1(\design_top.IADDR[7] ),
    .A2(_05958_),
    .B1(\design_top.core0.NXPC[7] ),
    .B2(_05959_),
    .X(_03098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13432_ (.A(_07727_),
    .X(_05960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13433_ (.A1(\design_top.IADDR[6] ),
    .A2(_05960_),
    .B1(\design_top.core0.NXPC[6] ),
    .B2(_05959_),
    .X(_03097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13434_ (.A1(\design_top.IADDR[5] ),
    .A2(_05960_),
    .B1(\design_top.core0.NXPC[5] ),
    .B2(_05959_),
    .X(_03096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13435_ (.A1(_07803_),
    .A2(_05960_),
    .B1(\design_top.core0.NXPC[4] ),
    .B2(_05959_),
    .X(_03095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13436_ (.A1(io_out[19]),
    .A2(_05960_),
    .B1(\design_top.core0.NXPC[3] ),
    .B2(_05959_),
    .X(_03094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13437_ (.A1(io_out[18]),
    .A2(_05960_),
    .B1(\design_top.core0.NXPC[2] ),
    .B2(_07767_),
    .X(_03093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13438_ (.A1(io_out[17]),
    .A2(_07720_),
    .B1(\design_top.core0.NXPC[1] ),
    .B2(_07767_),
    .X(_03092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13439_ (.A1(io_out[16]),
    .A2(_07720_),
    .B1(\design_top.core0.NXPC[0] ),
    .B2(_07767_),
    .X(_03091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13440_ (.A(_08544_),
    .X(_05961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13441_ (.A(_05961_),
    .X(_05962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13442_ (.A(_05962_),
    .X(_05963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13443_ (.A(_05961_),
    .Y(_05964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13444_ (.A(_05964_),
    .X(_05965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13445_ (.A(_05965_),
    .X(_05966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13446_ (.A1(_08089_),
    .A2(_05963_),
    .B1(\design_top.core0.REG2[9][31] ),
    .B2(_05966_),
    .X(_03090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13447_ (.A1(_08091_),
    .A2(_05963_),
    .B1(\design_top.core0.REG2[9][30] ),
    .B2(_05966_),
    .X(_03089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13448_ (.A1(_08093_),
    .A2(_05963_),
    .B1(\design_top.core0.REG2[9][29] ),
    .B2(_05966_),
    .X(_03088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13449_ (.A1(_08095_),
    .A2(_05963_),
    .B1(\design_top.core0.REG2[9][28] ),
    .B2(_05966_),
    .X(_03087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13450_ (.A1(_08098_),
    .A2(_05963_),
    .B1(\design_top.core0.REG2[9][27] ),
    .B2(_05966_),
    .X(_03086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13451_ (.A(_05962_),
    .X(_05967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13452_ (.A(_05965_),
    .X(_05968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13453_ (.A1(_08102_),
    .A2(_05967_),
    .B1(\design_top.core0.REG2[9][26] ),
    .B2(_05968_),
    .X(_03085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13454_ (.A1(_08104_),
    .A2(_05967_),
    .B1(\design_top.core0.REG2[9][25] ),
    .B2(_05968_),
    .X(_03084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13455_ (.A1(_08106_),
    .A2(_05967_),
    .B1(\design_top.core0.REG2[9][24] ),
    .B2(_05968_),
    .X(_03083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13456_ (.A1(_08108_),
    .A2(_05967_),
    .B1(\design_top.core0.REG2[9][23] ),
    .B2(_05968_),
    .X(_03082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13457_ (.A1(_08111_),
    .A2(_05967_),
    .B1(\design_top.core0.REG2[9][22] ),
    .B2(_05968_),
    .X(_03081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13458_ (.A(_05962_),
    .X(_05969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13459_ (.A(_05965_),
    .X(_05970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13460_ (.A1(_08115_),
    .A2(_05969_),
    .B1(\design_top.core0.REG2[9][21] ),
    .B2(_05970_),
    .X(_03080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13461_ (.A1(_08117_),
    .A2(_05969_),
    .B1(\design_top.core0.REG2[9][20] ),
    .B2(_05970_),
    .X(_03079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13462_ (.A1(_08119_),
    .A2(_05969_),
    .B1(\design_top.core0.REG2[9][19] ),
    .B2(_05970_),
    .X(_03078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13463_ (.A1(_08121_),
    .A2(_05969_),
    .B1(\design_top.core0.REG2[9][18] ),
    .B2(_05970_),
    .X(_03077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13464_ (.A1(_08124_),
    .A2(_05969_),
    .B1(\design_top.core0.REG2[9][17] ),
    .B2(_05970_),
    .X(_03076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13465_ (.A(_05961_),
    .X(_05971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13466_ (.A(_05964_),
    .X(_05972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13467_ (.A1(_08128_),
    .A2(_05971_),
    .B1(\design_top.core0.REG2[9][16] ),
    .B2(_05972_),
    .X(_03075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13468_ (.A1(_08130_),
    .A2(_05971_),
    .B1(\design_top.core0.REG2[9][15] ),
    .B2(_05972_),
    .X(_03074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13469_ (.A1(_08132_),
    .A2(_05971_),
    .B1(\design_top.core0.REG2[9][14] ),
    .B2(_05972_),
    .X(_03073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13470_ (.A1(\design_top.core0.REG2[9][13] ),
    .A2(_05962_),
    .B1(_08133_),
    .B2(_05965_),
    .X(_03072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13471_ (.A1(_08135_),
    .A2(_05971_),
    .B1(\design_top.core0.REG2[9][12] ),
    .B2(_05972_),
    .X(_03071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13472_ (.A1(_08138_),
    .A2(_05971_),
    .B1(\design_top.core0.REG2[9][11] ),
    .B2(_05972_),
    .X(_03070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13473_ (.A(_05961_),
    .X(_05973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13474_ (.A(_05964_),
    .X(_05974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13475_ (.A1(_08142_),
    .A2(_05973_),
    .B1(\design_top.core0.REG2[9][10] ),
    .B2(_05974_),
    .X(_03069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13476_ (.A1(_08144_),
    .A2(_05973_),
    .B1(\design_top.core0.REG2[9][9] ),
    .B2(_05974_),
    .X(_03068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13477_ (.A1(_08146_),
    .A2(_05973_),
    .B1(\design_top.core0.REG2[9][8] ),
    .B2(_05974_),
    .X(_03067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13478_ (.A1(_08148_),
    .A2(_05973_),
    .B1(\design_top.core0.REG2[9][7] ),
    .B2(_05974_),
    .X(_03066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13479_ (.A1(_08151_),
    .A2(_05973_),
    .B1(\design_top.core0.REG2[9][6] ),
    .B2(_05974_),
    .X(_03065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13480_ (.A(_05961_),
    .X(_05975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13481_ (.A(_05964_),
    .X(_05976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13482_ (.A1(_08155_),
    .A2(_05975_),
    .B1(\design_top.core0.REG2[9][5] ),
    .B2(_05976_),
    .X(_03064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13483_ (.A1(_08157_),
    .A2(_05975_),
    .B1(\design_top.core0.REG2[9][4] ),
    .B2(_05976_),
    .X(_03063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13484_ (.A1(_08159_),
    .A2(_05975_),
    .B1(\design_top.core0.REG2[9][3] ),
    .B2(_05976_),
    .X(_03062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13485_ (.A1(_08161_),
    .A2(_05975_),
    .B1(\design_top.core0.REG2[9][2] ),
    .B2(_05976_),
    .X(_03061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13486_ (.A1(_08163_),
    .A2(_05975_),
    .B1(\design_top.core0.REG2[9][1] ),
    .B2(_05976_),
    .X(_03060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13487_ (.A1(_08165_),
    .A2(_05962_),
    .B1(\design_top.core0.REG2[9][0] ),
    .B2(_05965_),
    .X(_03059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13488_ (.A(_06983_),
    .X(_05977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13489_ (.A(_05977_),
    .X(_01367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13490_ (.A(_05885_),
    .X(_05978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13491_ (.A(_05978_),
    .X(_01364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13492_ (.A(_06984_),
    .X(_05979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13493_ (.A(_05979_),
    .Y(_01372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13494_ (.A(_06984_),
    .X(_01373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13495_ (.A1_N(\design_top.IACK[7] ),
    .A2_N(\design_top.IREQ[7] ),
    .B1(\design_top.IACK[7] ),
    .B2(\design_top.IREQ[7] ),
    .X(_01376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13496_ (.A(\design_top.core0.FCT3[0] ),
    .Y(_05980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13497_ (.A(_07780_),
    .B(_05980_),
    .X(_05981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13498_ (.A(_05981_),
    .X(_01363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13499_ (.A(_05978_),
    .X(_05982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13500_ (.A(_05982_),
    .B(_01363_),
    .Y(_01377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _13501_ (.A1(_00802_),
    .A2(_06782_),
    .B1(_06783_),
    .C1(_06784_),
    .X(_05983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13502_ (.A(_05983_),
    .X(_05984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13503_ (.A(_05984_),
    .Y(_01378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13504_ (.A(_05983_),
    .X(_01379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13505_ (.A(_08016_),
    .X(_05985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13506_ (.A(_07052_),
    .B(_05985_),
    .Y(_01383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13507_ (.A(_07568_),
    .B(_05985_),
    .Y(_01384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13508_ (.A(_07554_),
    .B(_05985_),
    .Y(_01385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13509_ (.A(_07534_),
    .B(_05985_),
    .Y(_01386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13510_ (.A(_08016_),
    .X(_05986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13511_ (.A(_07493_),
    .B(_05986_),
    .Y(_01387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13512_ (.A(_07479_),
    .B(_05986_),
    .Y(_01388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13513_ (.A(_07459_),
    .B(_05986_),
    .Y(_01389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13514_ (.A(_06858_),
    .B(_05986_),
    .Y(_01390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13515_ (.A(_07414_),
    .B(_05986_),
    .Y(_01391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13516_ (.A(_07437_),
    .B(_05985_),
    .Y(_01392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13517_ (.A(_08016_),
    .X(_05987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13518_ (.A(_07404_),
    .B(_05987_),
    .Y(_01393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13519_ (.A(_07381_),
    .B(_05987_),
    .Y(_01394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13520_ (.A(_07364_),
    .B(_05987_),
    .Y(_01395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13521_ (.A(_07353_),
    .B(_05987_),
    .Y(_01396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13522_ (.A(_07319_),
    .B(_05987_),
    .Y(_01397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13523_ (.A(_08016_),
    .X(_05988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13524_ (.A(_05988_),
    .X(_05989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13525_ (.A(_07296_),
    .B(_05989_),
    .Y(_01398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13526_ (.A(_07281_),
    .B(_05989_),
    .Y(_01399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13527_ (.A(_07267_),
    .B(_05989_),
    .Y(_01400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13528_ (.A(_07251_),
    .B(_05989_),
    .Y(_01401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13529_ (.A(_07218_),
    .B(_05989_),
    .Y(_01402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13530_ (.A(_05988_),
    .X(_05990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13531_ (.A(_07194_),
    .B(_05990_),
    .Y(_01403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13532_ (.A(_07179_),
    .B(_05988_),
    .Y(_01404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13533_ (.A(_07169_),
    .B(_05990_),
    .Y(_01405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13534_ (.A(_07155_),
    .B(_05990_),
    .Y(_01406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13535_ (.A(_07128_),
    .B(_05990_),
    .Y(_01407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13536_ (.A(_07105_),
    .B(_05990_),
    .Y(_01408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13537_ (.A(_05988_),
    .X(_05991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13538_ (.A(_07080_),
    .B(_05991_),
    .Y(_01409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13539_ (.A(_07060_),
    .B(_05991_),
    .Y(_01410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13540_ (.A(_07044_),
    .B(_05991_),
    .Y(_01411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13541_ (.A(_01189_),
    .Y(_05992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13542_ (.A(_05992_),
    .X(_05993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13543_ (.A(_05993_),
    .B(_01373_),
    .Y(_01412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13544_ (.A(\design_top.core0.FCT3[2] ),
    .X(_05994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13545_ (.A(_05994_),
    .B(_01363_),
    .Y(_01362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13546_ (.A(_01080_),
    .Y(_05995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13547_ (.A(_05995_),
    .B(_01364_),
    .Y(_01413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13548_ (.A(_06664_),
    .Y(io_out[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13549_ (.A(_06972_),
    .B(_05991_),
    .Y(_01415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13550_ (.A(_06897_),
    .B(_05991_),
    .Y(_01416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13551_ (.A(\design_top.uart0.UART_XSTATE[0] ),
    .B(_07926_),
    .Y(_01417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13552_ (.A(_07629_),
    .B(_05988_),
    .Y(_01418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13553_ (.A(\design_top.DACK[1] ),
    .B(\design_top.DACK[0] ),
    .Y(_01419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13554_ (.A(_05886_),
    .X(_05996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13555_ (.A(_05996_),
    .Y(_01423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _13556_ (.A(_01260_),
    .B(_05982_),
    .C(_01367_),
    .X(_01424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13557_ (.A(_01260_),
    .Y(_05997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13558_ (.A(_05997_),
    .X(_05998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13559_ (.A(_07601_),
    .X(_05999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13560_ (.A(_05999_),
    .X(_06000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13561_ (.A(_05998_),
    .B(_06000_),
    .Y(_01425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _13562_ (.A(_01253_),
    .B(_05982_),
    .C(_01367_),
    .X(_01427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13563_ (.A(_01253_),
    .Y(_06001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13564_ (.A(_06001_),
    .X(_06002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13565_ (.A(_06002_),
    .B(_06000_),
    .Y(_01428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13566_ (.A(_05885_),
    .X(_06003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _13567_ (.A(_01245_),
    .B(_06003_),
    .C(_01367_),
    .X(_01430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13568_ (.A(_01245_),
    .Y(_06004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13569_ (.A(_06004_),
    .X(_06005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13570_ (.A(_06005_),
    .B(_06000_),
    .Y(_01431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _13571_ (.A(_01237_),
    .B(_06003_),
    .C(_01367_),
    .X(_01433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13572_ (.A(_01237_),
    .Y(_06006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13573_ (.A(_06006_),
    .X(_06007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13574_ (.A(_06007_),
    .B(_06000_),
    .Y(_01434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _13575_ (.A(_01229_),
    .B(_06003_),
    .C(_05977_),
    .X(_01436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13576_ (.A(_01229_),
    .Y(_06008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13577_ (.A(_06008_),
    .B(_06000_),
    .Y(_01437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _13578_ (.A(_01215_),
    .B(_06003_),
    .C(_05977_),
    .X(_01439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13579_ (.A(_01215_),
    .Y(_06009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13580_ (.A(_05999_),
    .X(_06010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13581_ (.A(_06009_),
    .B(_06010_),
    .Y(_01440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _13582_ (.A(_01203_),
    .B(_06003_),
    .C(_05977_),
    .X(_01442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13583_ (.A(_01203_),
    .Y(_06011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13584_ (.A(_06011_),
    .X(_06012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13585_ (.A(_06012_),
    .B(_06010_),
    .Y(_01443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _13586_ (.A(_01189_),
    .B(_05978_),
    .C(_05977_),
    .X(_01445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13587_ (.A(_05993_),
    .B(_06010_),
    .Y(_01446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13588_ (.A(_05998_),
    .B(_01379_),
    .Y(_01448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13589_ (.A(_01176_),
    .Y(_06013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13590_ (.A(_06013_),
    .B(_06010_),
    .Y(_01449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13591_ (.A(_06002_),
    .B(_01379_),
    .Y(_01451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13592_ (.A(_01161_),
    .Y(_06014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13593_ (.A(_06014_),
    .B(_06010_),
    .Y(_01452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13594_ (.A(_06005_),
    .B(_01379_),
    .Y(_01454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13595_ (.A(_01147_),
    .Y(_06015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13596_ (.A(_05999_),
    .X(_06016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13597_ (.A(_06015_),
    .B(_06016_),
    .Y(_01455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13598_ (.A(_06007_),
    .B(_01379_),
    .Y(_01457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13599_ (.A(_01133_),
    .Y(_06017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13600_ (.A(_06017_),
    .B(_06016_),
    .Y(_01458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13601_ (.A(_06008_),
    .B(_05984_),
    .Y(_01460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13602_ (.A(_01121_),
    .Y(_06018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13603_ (.A(_06018_),
    .B(_06016_),
    .Y(_01461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13604_ (.A(_06009_),
    .B(_05984_),
    .Y(_01463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13605_ (.A(_01107_),
    .Y(_06019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13606_ (.A(_06019_),
    .B(_06016_),
    .Y(_01464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13607_ (.A(_06012_),
    .B(_05984_),
    .Y(_01466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13608_ (.A(_01094_),
    .Y(_06020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13609_ (.A(_06020_),
    .B(_06016_),
    .Y(_01467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13610_ (.A(_05993_),
    .B(_05984_),
    .Y(_01469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13611_ (.A(_05995_),
    .B(_05999_),
    .Y(_01470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13612_ (.A(_05886_),
    .X(_01368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13613_ (.A(_05998_),
    .B(_01368_),
    .Y(_01472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13614_ (.A(_05998_),
    .B(_01364_),
    .Y(_01473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13615_ (.A(_06002_),
    .B(_01368_),
    .Y(_01475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13616_ (.A(_06002_),
    .B(_01364_),
    .Y(_01476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13617_ (.A(_06005_),
    .B(_01368_),
    .Y(_01478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13618_ (.A(_06005_),
    .B(_01364_),
    .Y(_01479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13619_ (.A(_06007_),
    .B(_01368_),
    .Y(_01481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13620_ (.A(_05978_),
    .X(_06021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13621_ (.A(_06007_),
    .B(_06021_),
    .Y(_01482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13622_ (.A(_06008_),
    .B(_05996_),
    .Y(_01484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13623_ (.A(_06008_),
    .B(_06021_),
    .Y(_01485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13624_ (.A(_06009_),
    .B(_05996_),
    .Y(_01487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13625_ (.A(_06009_),
    .B(_06021_),
    .Y(_01488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13626_ (.A(_06012_),
    .B(_05996_),
    .Y(_01490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13627_ (.A(_06012_),
    .B(_06021_),
    .Y(_01491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13628_ (.A(_05993_),
    .B(_05996_),
    .Y(_01493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13629_ (.A(_05993_),
    .B(_06021_),
    .Y(_01494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13630_ (.A(_05998_),
    .B(_01373_),
    .Y(_01496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13631_ (.A(_05978_),
    .X(_06022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13632_ (.A(_06013_),
    .B(_06022_),
    .Y(_01497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13633_ (.A(_06002_),
    .B(_01373_),
    .Y(_01499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13634_ (.A(_06014_),
    .B(_06022_),
    .Y(_01500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13635_ (.A(_06005_),
    .B(_01373_),
    .Y(_01502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13636_ (.A(_06015_),
    .B(_06022_),
    .Y(_01503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13637_ (.A(_06007_),
    .B(_05979_),
    .Y(_01505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13638_ (.A(_06017_),
    .B(_06022_),
    .Y(_01506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13639_ (.A(_06008_),
    .B(_05979_),
    .Y(_01508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13640_ (.A(_06018_),
    .B(_06022_),
    .Y(_01509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13641_ (.A(_06009_),
    .B(_05979_),
    .Y(_01511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13642_ (.A(_06019_),
    .B(_05982_),
    .Y(_01512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13643_ (.A(_06012_),
    .B(_05979_),
    .Y(_01514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13644_ (.A(_06020_),
    .B(_05982_),
    .Y(_01515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13645_ (.A(\design_top.core0.RESMODE[1] ),
    .Y(_06023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13646_ (.A(_07992_),
    .B(_06023_),
    .Y(_01517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13647_ (.A(_06658_),
    .B(_06659_),
    .Y(_01519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13648_ (.A(\design_top.core0.NXPC[0] ),
    .Y(_01520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13649_ (.A1(_06786_),
    .A2(_00805_),
    .B1(_06787_),
    .B2(_00808_),
    .X(_06024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13650_ (.A(_06024_),
    .Y(_01290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13651_ (.A(_01261_),
    .Y(_06025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13652_ (.A(_06025_),
    .B(_01290_),
    .X(_06026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13653_ (.A(_06026_),
    .X(_01521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13654_ (.A(_01261_),
    .X(_06027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13655_ (.A(_06027_),
    .B(_06024_),
    .Y(_01522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _13656_ (.A(\design_top.core0.FCT3[1] ),
    .B(\design_top.core0.FCT3[0] ),
    .C(_07809_),
    .X(_06028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13657_ (.A(_06028_),
    .X(_06029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13658_ (.A(_06029_),
    .X(_01523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _13659_ (.A(_07780_),
    .B(_05980_),
    .C(_07809_),
    .X(_06030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13660_ (.A(_06030_),
    .X(_06031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13661_ (.A(_06031_),
    .X(_01524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13662_ (.A(_07753_),
    .B(_07770_),
    .Y(_01525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13663_ (.A(_06027_),
    .B(_01290_),
    .X(_01526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13664_ (.A(_01254_),
    .X(_06032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13665_ (.A(_06032_),
    .B(_01526_),
    .X(_01527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13666_ (.A(_01246_),
    .X(_06033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13667_ (.A(_06033_),
    .X(_06034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13668_ (.A(_06034_),
    .B(_01527_),
    .X(_01528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13669_ (.A(_01238_),
    .X(_06035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13670_ (.A(_06035_),
    .X(_06036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13671_ (.A(_06036_),
    .B(_01528_),
    .X(_01529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13672_ (.A(_01230_),
    .X(_06037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13673_ (.A(_06037_),
    .X(_06038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13674_ (.A(_06038_),
    .B(_01529_),
    .X(_01530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13675_ (.A(_06773_),
    .X(_01534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13676_ (.A(_01563_),
    .X(_01564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13677_ (.A(\design_top.RAMFF[0] ),
    .Y(_01571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _13678_ (.A1_N(\design_top.uart0.UART_XREQ ),
    .A2_N(_08012_),
    .B1(\design_top.uart0.UART_XREQ ),
    .B2(_08012_),
    .X(_01572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13679_ (.A(\design_top.XADDR[2] ),
    .B(\design_top.XADDR[3] ),
    .Y(_01573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13680_ (.A(\design_top.IOMUX[3][0] ),
    .Y(_06039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13681_ (.A(\design_top.XADDR[2] ),
    .Y(_01582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13682_ (.A(\design_top.XADDR[3] ),
    .Y(_06040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13683_ (.A(_01582_),
    .B(_06040_),
    .X(_06041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13684_ (.A(_06041_),
    .X(_06042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13685_ (.A(io_out[8]),
    .Y(_06043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13686_ (.A(\design_top.XADDR[2] ),
    .B(_06040_),
    .X(_06044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13687_ (.A(_06044_),
    .X(_06045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _13688_ (.A(_01582_),
    .B(\design_top.XADDR[3] ),
    .C(_01572_),
    .X(_06046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _13689_ (.A1(_06039_),
    .A2(_06042_),
    .B1(_06043_),
    .B2(_06045_),
    .C1(_06046_),
    .X(_01574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13690_ (.A(\design_top.RAMFF[16] ),
    .Y(_01576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13691_ (.A(\design_top.IOMUX[3][16] ),
    .Y(_06047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13692_ (.A(_06041_),
    .X(_06048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13693_ (.A(_06048_),
    .X(_06049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13694_ (.A(io_out[15]),
    .Y(_06050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13695_ (.A(_06044_),
    .X(_06051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13696_ (.A(_06051_),
    .X(_06052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13697_ (.A1(_06047_),
    .A2(_06049_),
    .B1(_06050_),
    .B2(_06052_),
    .X(_01577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13698_ (.A(\design_top.RAMFF[24] ),
    .Y(_01581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13699_ (.A(\design_top.IOMUX[3][24] ),
    .Y(_06053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13700_ (.A(\design_top.GPIOFF[8] ),
    .Y(_06054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13701_ (.A1(_06053_),
    .A2(_06049_),
    .B1(_06054_),
    .B2(_06052_),
    .X(_01583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13702_ (.A(\design_top.RAMFF[8] ),
    .Y(_01586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13703_ (.A(\design_top.IOMUX[3][8] ),
    .Y(_06055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13704_ (.A(\design_top.LEDFF[8] ),
    .Y(_06056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13705_ (.A(_01582_),
    .B(\design_top.XADDR[3] ),
    .Y(_06057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13706_ (.A(_06057_),
    .X(_06058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _13707_ (.A(\design_top.uart0.UART_RFIFO[0] ),
    .B(_06058_),
    .Y(_06059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _13708_ (.A1(_06055_),
    .A2(_06042_),
    .B1(_06056_),
    .B2(_06045_),
    .C1(_06059_),
    .X(_01587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _13709_ (.A(_06658_),
    .B(_06659_),
    .C(\design_top.core0.XLUI ),
    .X(_01593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _13710_ (.A(_06658_),
    .B(_06659_),
    .C(\design_top.core0.XAUIPC ),
    .X(_01596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _13711_ (.A(\design_top.core0.SIMM[0] ),
    .B(\design_top.core0.PC[0] ),
    .Y(_06060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _13712_ (.A1(\design_top.core0.SIMM[0] ),
    .A2(\design_top.core0.PC[0] ),
    .B1(_06060_),
    .Y(_01597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13713_ (.A(\design_top.core0.NXPC[1] ),
    .Y(_01603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _13714_ (.A(_01254_),
    .B(_06781_),
    .Y(_01604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13715_ (.A(_07811_),
    .Y(_01248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13716_ (.A(_07812_),
    .Y(_01255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a32o_2 _13717_ (.A1(_06027_),
    .A2(_06024_),
    .A3(_07813_),
    .B1(_01255_),
    .B2(_01521_),
    .X(_01606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13718_ (.A(_06025_),
    .B(_00809_),
    .Y(_06061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13719_ (.A1_N(_07813_),
    .A2_N(_06061_),
    .B1(_07813_),
    .B2(_06061_),
    .X(_01607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13720_ (.A(_06032_),
    .B(_01608_),
    .X(_01609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13721_ (.A(_06034_),
    .B(_01609_),
    .X(_01610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13722_ (.A(_06036_),
    .B(_01610_),
    .X(_01611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13723_ (.A(_06038_),
    .B(_01611_),
    .X(_01612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13724_ (.A(_00843_),
    .X(_06062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13725_ (.A(_06027_),
    .B(_06062_),
    .X(_01639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _13726_ (.A(_01647_),
    .B(_01523_),
    .C(_01524_),
    .X(_01648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13727_ (.A(\design_top.RAMFF[1] ),
    .Y(_01651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13728_ (.A(\design_top.IOMUX[3][1] ),
    .Y(_06063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13729_ (.A(io_out[9]),
    .Y(_06064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _13730_ (.A1(\design_top.uart0.UART_RACK ),
    .A2(\design_top.uart0.UART_RREQ ),
    .B1(_06057_),
    .Y(_06065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _13731_ (.A1(\design_top.uart0.UART_RACK ),
    .A2(\design_top.uart0.UART_RREQ ),
    .B1(_06065_),
    .X(_06066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _13732_ (.A1(_06063_),
    .A2(_06042_),
    .B1(_06064_),
    .B2(_06045_),
    .C1(_06066_),
    .X(_01652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13733_ (.A(\design_top.RAMFF[17] ),
    .Y(_01654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13734_ (.A(\design_top.IOMUX[3][17] ),
    .Y(_06067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13735_ (.A(\design_top.GPIOFF[1] ),
    .Y(_06068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13736_ (.A1(_06067_),
    .A2(_06049_),
    .B1(_06068_),
    .B2(_06052_),
    .X(_01655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13737_ (.A(\design_top.RAMFF[25] ),
    .Y(_01659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13738_ (.A(\design_top.IOMUX[3][25] ),
    .Y(_06069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13739_ (.A(\design_top.GPIOFF[9] ),
    .Y(_06070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13740_ (.A1(_06069_),
    .A2(_06049_),
    .B1(_06070_),
    .B2(_06052_),
    .X(_01660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13741_ (.A(\design_top.RAMFF[9] ),
    .Y(_01663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13742_ (.A(\design_top.IOMUX[3][9] ),
    .Y(_06071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13743_ (.A(_06041_),
    .X(_06072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13744_ (.A(\design_top.LEDFF[9] ),
    .Y(_06073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13745_ (.A(_06044_),
    .X(_06074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _13746_ (.A(\design_top.uart0.UART_RFIFO[1] ),
    .B(_06058_),
    .Y(_06075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _13747_ (.A1(_06071_),
    .A2(_06072_),
    .B1(_06073_),
    .B2(_06074_),
    .C1(_06075_),
    .X(_01664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13748_ (.A(_06780_),
    .Y(_00801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13749_ (.A(\design_top.core0.PC[1] ),
    .Y(_06076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13750_ (.A1(_00801_),
    .A2(_06076_),
    .B1(_06780_),
    .B2(\design_top.core0.PC[1] ),
    .X(_06077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13751_ (.A(_06077_),
    .Y(_06078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a32o_2 _13752_ (.A1(\design_top.core0.SIMM[0] ),
    .A2(\design_top.core0.PC[0] ),
    .A3(_06077_),
    .B1(_06060_),
    .B2(_06078_),
    .X(_01672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13753_ (.A(\design_top.core0.NXPC[2] ),
    .Y(_01674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _13754_ (.A(_06033_),
    .B(_07826_),
    .Y(_01675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13755_ (.A(_07828_),
    .Y(_01292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _13756_ (.A1(_01255_),
    .A2(_01521_),
    .B1(_01604_),
    .Y(_06079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13757_ (.A(_06079_),
    .Y(_06080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13758_ (.A1(_07828_),
    .A2(_06079_),
    .B1(_01292_),
    .B2(_06080_),
    .X(_01676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13759_ (.A1(_06032_),
    .A2(_01248_),
    .B1(_07813_),
    .B2(_06061_),
    .X(_06081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13760_ (.A1_N(_07828_),
    .A2_N(_06081_),
    .B1(_07828_),
    .B2(_06081_),
    .X(_01677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13761_ (.A(_06034_),
    .B(_01679_),
    .X(_01680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13762_ (.A(_06036_),
    .B(_01680_),
    .X(_01681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13763_ (.A(_06038_),
    .B(_01681_),
    .X(_01682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13764_ (.A(_06032_),
    .B(_01559_),
    .X(_01694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13765_ (.A(_06841_),
    .X(_06082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _13766_ (.A(_06082_),
    .B(_00849_),
    .Y(_00851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _13767_ (.A(_01701_),
    .B(_01523_),
    .C(_01524_),
    .X(_01702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13768_ (.A(\design_top.RAMFF[2] ),
    .Y(_01705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13769_ (.A(\design_top.IOMUX[3][2] ),
    .Y(_06083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13770_ (.A(io_out[10]),
    .Y(_06084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13771_ (.A1(_06083_),
    .A2(_06049_),
    .B1(_06084_),
    .B2(_06052_),
    .X(_01706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13772_ (.A(\design_top.RAMFF[18] ),
    .Y(_01708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13773_ (.A(\design_top.IOMUX[3][18] ),
    .Y(_06085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13774_ (.A(_06048_),
    .X(_06086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13775_ (.A(\design_top.GPIOFF[2] ),
    .Y(_06087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13776_ (.A(_06051_),
    .X(_06088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13777_ (.A1(_06085_),
    .A2(_06086_),
    .B1(_06087_),
    .B2(_06088_),
    .X(_01709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13778_ (.A(\design_top.RAMFF[26] ),
    .Y(_01714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13779_ (.A(\design_top.IOMUX[3][26] ),
    .Y(_06089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13780_ (.A(\design_top.GPIOFF[10] ),
    .Y(_06090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13781_ (.A1(_06089_),
    .A2(_06086_),
    .B1(_06090_),
    .B2(_06088_),
    .X(_01715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13782_ (.A(\design_top.RAMFF[10] ),
    .Y(_01717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13783_ (.A(\design_top.IOMUX[3][10] ),
    .Y(_06091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13784_ (.A(\design_top.LEDFF[10] ),
    .Y(_06092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _13785_ (.A1(\design_top.uart0.UART_RFIFO[2] ),
    .A2(_06057_),
    .B1(_01573_),
    .Y(_06093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _13786_ (.A1(_06091_),
    .A2(_06072_),
    .B1(_06092_),
    .B2(_06074_),
    .C1(_06093_),
    .X(_01718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13787_ (.A1(_00801_),
    .A2(_06076_),
    .B1(_06060_),
    .B2(_06078_),
    .X(_06094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13788_ (.A(_06792_),
    .B(\design_top.core0.PC[2] ),
    .Y(_06095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _13789_ (.A1(_06792_),
    .A2(\design_top.core0.PC[2] ),
    .B1(_06095_),
    .X(_06096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _13790_ (.A1_N(_06094_),
    .A2_N(_06096_),
    .B1(_06094_),
    .B2(_06096_),
    .X(_02471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13791_ (.A(_02471_),
    .Y(_01726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13792_ (.A(\design_top.core0.NXPC[3] ),
    .Y(_01728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13793_ (.A(_07824_),
    .Y(_01293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _13794_ (.A1(_01675_),
    .A2(_06080_),
    .B1(_01247_),
    .X(_06097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13795_ (.A1_N(_01293_),
    .A2_N(_06097_),
    .B1(_01293_),
    .B2(_06097_),
    .X(_01729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13796_ (.A1(_07827_),
    .A2(_06081_),
    .B1(_01246_),
    .B2(_00793_),
    .X(_06098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _13797_ (.A(_01238_),
    .B(_06779_),
    .Y(_01240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13798_ (.A1(_01238_),
    .A2(_07823_),
    .B1(_01240_),
    .X(_06099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13799_ (.A1_N(_06098_),
    .A2_N(_06099_),
    .B1(_06098_),
    .B2(_06099_),
    .X(_01730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13800_ (.A(_06034_),
    .B(_01732_),
    .X(_01733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13801_ (.A(_06036_),
    .B(_01733_),
    .X(_01734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13802_ (.A(_06038_),
    .B(_01734_),
    .X(_01735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13803_ (.A(_06032_),
    .B(_01639_),
    .X(_01747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13804_ (.A(_01068_),
    .B(_06718_),
    .Y(_01069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _13805_ (.A(_01753_),
    .B(_01523_),
    .C(_01524_),
    .X(_01754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13806_ (.A(\design_top.RAMFF[3] ),
    .Y(_01757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13807_ (.A(\design_top.IOMUX[3][3] ),
    .Y(_06100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13808_ (.A(io_out[11]),
    .Y(_06101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13809_ (.A1(_06100_),
    .A2(_06086_),
    .B1(_06101_),
    .B2(_06088_),
    .X(_01758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13810_ (.A(\design_top.RAMFF[19] ),
    .Y(_01760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13811_ (.A(\design_top.IOMUX[3][19] ),
    .Y(_06102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13812_ (.A(\design_top.GPIOFF[3] ),
    .Y(_06103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13813_ (.A1(_06102_),
    .A2(_06086_),
    .B1(_06103_),
    .B2(_06088_),
    .X(_01761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13814_ (.A(\design_top.RAMFF[27] ),
    .Y(_01765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13815_ (.A(\design_top.IOMUX[3][27] ),
    .Y(_06104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13816_ (.A(\design_top.GPIOFF[11] ),
    .Y(_06105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13817_ (.A1(_06104_),
    .A2(_06086_),
    .B1(_06105_),
    .B2(_06088_),
    .X(_01766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13818_ (.A(\design_top.RAMFF[11] ),
    .Y(_01768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13819_ (.A(\design_top.IOMUX[3][11] ),
    .Y(_06106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13820_ (.A(\design_top.LEDFF[11] ),
    .Y(_06107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _13821_ (.A(\design_top.uart0.UART_RFIFO[3] ),
    .B(_06058_),
    .Y(_06108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _13822_ (.A1(_06106_),
    .A2(_06072_),
    .B1(_06107_),
    .B2(_06074_),
    .C1(_06108_),
    .X(_01769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13823_ (.A(_06815_),
    .X(_01062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _13824_ (.A1_N(_06792_),
    .A2_N(\design_top.core0.PC[2] ),
    .B1(_06094_),
    .B2(_06095_),
    .X(_06109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13825_ (.A(\design_top.core0.SIMM[3] ),
    .B(\design_top.core0.PC[3] ),
    .Y(_06110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _13826_ (.A1(_06847_),
    .A2(\design_top.core0.PC[3] ),
    .B1(_06110_),
    .X(_06111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _13827_ (.A1_N(_06109_),
    .A2_N(_06111_),
    .B1(_06109_),
    .B2(_06111_),
    .X(_02474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13828_ (.A(_02474_),
    .Y(_01777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13829_ (.A(\design_top.core0.NXPC[4] ),
    .Y(_01779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13830_ (.A(_07818_),
    .X(_01294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13831_ (.A1(_01293_),
    .A2(_06097_),
    .B1(_01240_),
    .X(_06112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13832_ (.A1_N(_01294_),
    .A2_N(_06112_),
    .B1(_01294_),
    .B2(_06112_),
    .X(_01781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13833_ (.A(_07823_),
    .Y(_01232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13834_ (.A1(_06035_),
    .A2(_01232_),
    .B1(_06098_),
    .B2(_06099_),
    .X(_06113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13835_ (.A1_N(_07819_),
    .A2_N(_06113_),
    .B1(_07819_),
    .B2(_06113_),
    .X(_01782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13836_ (.A(_06036_),
    .B(_01785_),
    .X(_01786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13837_ (.A(_06037_),
    .X(_06114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13838_ (.A(_06114_),
    .X(_06115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13839_ (.A(_06115_),
    .B(_01786_),
    .X(_01787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13840_ (.A(_06034_),
    .B(_01560_),
    .X(_01792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _13841_ (.A(_01797_),
    .B(_01523_),
    .C(_01524_),
    .X(_01798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13842_ (.A(\design_top.RAMFF[4] ),
    .Y(_01801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13843_ (.A(\design_top.IOMUX[3][4] ),
    .Y(_06116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13844_ (.A(_06048_),
    .X(_06117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13845_ (.A(\design_top.LEDFF[4] ),
    .Y(_06118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13846_ (.A(_06051_),
    .X(_06119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13847_ (.A1(_06116_),
    .A2(_06117_),
    .B1(_06118_),
    .B2(_06119_),
    .X(_01802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13848_ (.A(\design_top.RAMFF[20] ),
    .Y(_01804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13849_ (.A(\design_top.IOMUX[3][20] ),
    .Y(_06120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13850_ (.A(\design_top.GPIOFF[4] ),
    .Y(_06121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13851_ (.A1(_06120_),
    .A2(_06117_),
    .B1(_06121_),
    .B2(_06119_),
    .X(_01805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13852_ (.A(\design_top.RAMFF[28] ),
    .Y(_01809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13853_ (.A(\design_top.IOMUX[3][28] ),
    .Y(_06122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13854_ (.A(\design_top.GPIOFF[12] ),
    .Y(_06123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13855_ (.A1(_06122_),
    .A2(_06117_),
    .B1(_06123_),
    .B2(_06119_),
    .X(_01810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13856_ (.A(\design_top.RAMFF[12] ),
    .Y(_01812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13857_ (.A(\design_top.IOMUX[3][12] ),
    .Y(_06124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13858_ (.A(\design_top.LEDFF[12] ),
    .Y(_06125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _13859_ (.A(\design_top.uart0.UART_RFIFO[4] ),
    .B(_06058_),
    .Y(_06126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _13860_ (.A1(_06124_),
    .A2(_06072_),
    .B1(_06125_),
    .B2(_06074_),
    .C1(_06126_),
    .X(_01813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _13861_ (.A1_N(_06847_),
    .A2_N(\design_top.core0.PC[3] ),
    .B1(_06109_),
    .B2(_06110_),
    .X(_06127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13862_ (.A1_N(_06853_),
    .A2_N(\design_top.core0.PC[4] ),
    .B1(\design_top.core0.SIMM[4] ),
    .B2(\design_top.core0.PC[4] ),
    .X(_06128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13863_ (.A(_06127_),
    .Y(_06129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13864_ (.A(_06128_),
    .Y(_06130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13865_ (.A1(_06127_),
    .A2(_06128_),
    .B1(_06129_),
    .B2(_06130_),
    .X(_02477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13866_ (.A(_02477_),
    .Y(_01821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13867_ (.A(\design_top.core0.NXPC[5] ),
    .Y(_01823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13868_ (.A(_07817_),
    .Y(_01295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13869_ (.A1(_01294_),
    .A2(_06112_),
    .B1(_01780_),
    .X(_06131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13870_ (.A1_N(_01295_),
    .A2_N(_06131_),
    .B1(_01295_),
    .B2(_06131_),
    .X(_01824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13871_ (.A(_06776_),
    .X(_01224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13872_ (.A1(_07819_),
    .A2(_06113_),
    .B1(_01230_),
    .B2(_01224_),
    .X(_06132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13873_ (.A1_N(_07817_),
    .A2_N(_06132_),
    .B1(_07817_),
    .B2(_06132_),
    .X(_01825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13874_ (.A(_06035_),
    .X(_06133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13875_ (.A(_06133_),
    .B(_01828_),
    .X(_01829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13876_ (.A(_06115_),
    .B(_01829_),
    .X(_01830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13877_ (.A(_06033_),
    .B(_01640_),
    .X(_01835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13878_ (.A(_06029_),
    .X(_06134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13879_ (.A(_06031_),
    .X(_06135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _13880_ (.A(_01840_),
    .B(_06134_),
    .C(_06135_),
    .X(_01841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13881_ (.A(\design_top.RAMFF[5] ),
    .Y(_01844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13882_ (.A(\design_top.IOMUX[3][5] ),
    .Y(_06136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13883_ (.A(\design_top.LEDFF[5] ),
    .Y(_06137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13884_ (.A1(_06136_),
    .A2(_06117_),
    .B1(_06137_),
    .B2(_06119_),
    .X(_01845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13885_ (.A(\design_top.RAMFF[21] ),
    .Y(_01847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13886_ (.A(\design_top.IOMUX[3][21] ),
    .Y(_06138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13887_ (.A(\design_top.GPIOFF[5] ),
    .Y(_06139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13888_ (.A1(_06138_),
    .A2(_06117_),
    .B1(_06139_),
    .B2(_06119_),
    .X(_01848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13889_ (.A(\design_top.RAMFF[29] ),
    .Y(_01853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13890_ (.A(\design_top.IOMUX[3][29] ),
    .Y(_06140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13891_ (.A(_06041_),
    .X(_06141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13892_ (.A(\design_top.GPIOFF[13] ),
    .Y(_06142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13893_ (.A(_06044_),
    .X(_06143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13894_ (.A1(_06140_),
    .A2(_06141_),
    .B1(_06142_),
    .B2(_06143_),
    .X(_01854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13895_ (.A(\design_top.RAMFF[13] ),
    .Y(_01856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13896_ (.A(\design_top.IOMUX[3][13] ),
    .Y(_06144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13897_ (.A(\design_top.LEDFF[13] ),
    .Y(_06145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _13898_ (.A1(\design_top.uart0.UART_RFIFO[5] ),
    .A2(_06057_),
    .B1(_01573_),
    .Y(_06146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _13899_ (.A1(_06144_),
    .A2(_06072_),
    .B1(_06145_),
    .B2(_06074_),
    .C1(_06146_),
    .X(_01857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13900_ (.A(_06767_),
    .B(\design_top.core0.PC[5] ),
    .X(_06147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _13901_ (.A1(_06767_),
    .A2(\design_top.core0.PC[5] ),
    .B1_N(_06147_),
    .Y(_06148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13902_ (.A1(_06853_),
    .A2(\design_top.core0.PC[4] ),
    .B1(_06129_),
    .B2(_06130_),
    .X(_06149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _13903_ (.A1_N(_06148_),
    .A2_N(_06149_),
    .B1(_06148_),
    .B2(_06149_),
    .X(_02481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13904_ (.A(_02481_),
    .Y(_01865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13905_ (.A(\design_top.core0.NXPC[6] ),
    .Y(_01867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13906_ (.A(_07820_),
    .X(_01296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _13907_ (.A(_06768_),
    .B(_01216_),
    .Y(_01218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _13908_ (.A(_01295_),
    .B(_01294_),
    .C(_06112_),
    .X(_06150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _13909_ (.A1(_01218_),
    .A2(_01780_),
    .B1(_01217_),
    .X(_06151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _13910_ (.A(_06150_),
    .B(_06151_),
    .X(_06152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13911_ (.A1_N(_01296_),
    .A2_N(_06152_),
    .B1(_01296_),
    .B2(_06152_),
    .X(_01869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13912_ (.A1(_07817_),
    .A2(_06132_),
    .B1(_01534_),
    .B2(_01216_),
    .X(_06153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13913_ (.A1_N(_07821_),
    .A2_N(_06153_),
    .B1(_07821_),
    .B2(_06153_),
    .X(_01870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13914_ (.A(_06133_),
    .B(_01873_),
    .X(_01874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13915_ (.A(_06115_),
    .B(_01874_),
    .X(_01875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13916_ (.A(_06033_),
    .B(_01694_),
    .X(_01880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13917_ (.A(\design_top.core0.REG1[14][31] ),
    .Y(_00840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13918_ (.A(\design_top.core0.REG1[15][31] ),
    .Y(_00841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _13919_ (.A(_01885_),
    .B(_06134_),
    .C(_06135_),
    .X(_01886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13920_ (.A(\design_top.RAMFF[6] ),
    .Y(_01889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13921_ (.A(\design_top.IOMUX[3][6] ),
    .Y(_06154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13922_ (.A(\design_top.LEDFF[6] ),
    .Y(_06155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13923_ (.A1(_06154_),
    .A2(_06141_),
    .B1(_06155_),
    .B2(_06143_),
    .X(_01890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13924_ (.A(\design_top.RAMFF[22] ),
    .Y(_01892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13925_ (.A(\design_top.IOMUX[3][22] ),
    .Y(_06156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13926_ (.A(\design_top.GPIOFF[6] ),
    .Y(_06157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13927_ (.A1(_06156_),
    .A2(_06141_),
    .B1(_06157_),
    .B2(_06143_),
    .X(_01893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13928_ (.A(\design_top.RAMFF[30] ),
    .Y(_01898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13929_ (.A(\design_top.IOMUX[3][30] ),
    .Y(_06158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13930_ (.A(\design_top.GPIOFF[14] ),
    .Y(_06159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13931_ (.A1(_06158_),
    .A2(_06141_),
    .B1(_06159_),
    .B2(_06143_),
    .X(_01899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13932_ (.A(\design_top.RAMFF[14] ),
    .Y(_01901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13933_ (.A(\design_top.IOMUX[3][14] ),
    .Y(_06160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13934_ (.A(\design_top.LEDFF[14] ),
    .Y(_06161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _13935_ (.A1(\design_top.uart0.UART_RFIFO[6] ),
    .A2(_06057_),
    .B1(_01573_),
    .Y(_06162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _13936_ (.A1(_06160_),
    .A2(_06048_),
    .B1(_06161_),
    .B2(_06051_),
    .C1(_06162_),
    .X(_01902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13937_ (.A(\design_top.core0.REG1[13][31] ),
    .Y(_00839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a32o_2 _13938_ (.A1(_06853_),
    .A2(\design_top.core0.PC[4] ),
    .A3(_06147_),
    .B1(_06767_),
    .B2(\design_top.core0.PC[5] ),
    .X(_06163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _13939_ (.A1(_06130_),
    .A2(_06148_),
    .A3(_06129_),
    .B1(_06163_),
    .X(_06164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13940_ (.A(\design_top.core0.PC[6] ),
    .Y(_06165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13941_ (.A1(_06760_),
    .A2(\design_top.core0.PC[6] ),
    .B1(_01336_),
    .B2(_06165_),
    .X(_06166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _13942_ (.A1_N(_06164_),
    .A2_N(_06166_),
    .B1(_06164_),
    .B2(_06166_),
    .X(_02485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13943_ (.A(_02485_),
    .Y(_01910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13944_ (.A(\design_top.core0.NXPC[7] ),
    .Y(_01912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13945_ (.A(_07814_),
    .X(_01297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _13946_ (.A1(_01296_),
    .A2(_06152_),
    .B1(_01868_),
    .X(_06167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13947_ (.A1_N(_01297_),
    .A2_N(_06167_),
    .B1(_01297_),
    .B2(_06167_),
    .X(_01913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13948_ (.A(_06758_),
    .X(_01198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13949_ (.A1(_07821_),
    .A2(_06153_),
    .B1(_01198_),
    .B2(_01204_),
    .X(_06168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13950_ (.A(_06168_),
    .Y(_06169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13951_ (.A1(_01297_),
    .A2(_06168_),
    .B1(_07815_),
    .B2(_06169_),
    .X(_01914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13952_ (.A(_06133_),
    .B(_01917_),
    .X(_01918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13953_ (.A(_06115_),
    .B(_01918_),
    .X(_01919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13954_ (.A(_06033_),
    .B(_01747_),
    .X(_01924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13955_ (.A(\design_top.core0.REG1[11][31] ),
    .Y(_00836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13956_ (.A(\design_top.core0.REG1[12][31] ),
    .Y(_00838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _13957_ (.A(_01928_),
    .B(_06134_),
    .C(_06135_),
    .X(_01929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13958_ (.A(\design_top.RAMFF[7] ),
    .Y(_01932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13959_ (.A(\design_top.IOMUX[3][7] ),
    .Y(_06170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13960_ (.A(\design_top.LEDFF[7] ),
    .Y(_06171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13961_ (.A1(_06170_),
    .A2(_06141_),
    .B1(_06171_),
    .B2(_06143_),
    .X(_01933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13962_ (.A(\design_top.RAMFF[23] ),
    .Y(_01935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13963_ (.A(\design_top.IOMUX[3][23] ),
    .Y(_06172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13964_ (.A(\design_top.GPIOFF[7] ),
    .Y(_06173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13965_ (.A1(_06172_),
    .A2(_06042_),
    .B1(_06173_),
    .B2(_06045_),
    .X(_01936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13966_ (.A(\design_top.RAMFF[31] ),
    .Y(_01940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13967_ (.A(\design_top.IOMUX[3][31] ),
    .Y(_06174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13968_ (.A(\design_top.GPIOFF[15] ),
    .Y(_06175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13969_ (.A1(_06174_),
    .A2(_06042_),
    .B1(_06175_),
    .B2(_06045_),
    .X(_01941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13970_ (.A(\design_top.RAMFF[15] ),
    .Y(_01944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13971_ (.A(\design_top.IOMUX[3][15] ),
    .Y(_06176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13972_ (.A(\design_top.LEDFF[15] ),
    .Y(_06177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _13973_ (.A(\design_top.uart0.UART_RFIFO[7] ),
    .B(_06058_),
    .Y(_06178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _13974_ (.A1(_06176_),
    .A2(_06048_),
    .B1(_06177_),
    .B2(_06051_),
    .C1(_06178_),
    .X(_01945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13975_ (.A(_06763_),
    .B(\design_top.core0.PC[7] ),
    .X(_06179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _13976_ (.A1(_06763_),
    .A2(\design_top.core0.PC[7] ),
    .B1_N(_06179_),
    .Y(_06180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _13977_ (.A1(_06760_),
    .A2(\design_top.core0.PC[6] ),
    .B1(_06164_),
    .B2(_06166_),
    .X(_06181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _13978_ (.A1_N(_06180_),
    .A2_N(_06181_),
    .B1(_06180_),
    .B2(_06181_),
    .X(_02488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13979_ (.A(_02488_),
    .Y(_01953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13980_ (.A(\design_top.core0.REG1[10][31] ),
    .Y(_00835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13981_ (.A(\design_top.core0.NXPC[8] ),
    .Y(_01955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _13982_ (.A(_07844_),
    .X(_01298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13983_ (.A(_06764_),
    .B(_01190_),
    .Y(_01191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _13984_ (.A(_06761_),
    .B(_01204_),
    .Y(_01205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _13985_ (.A1(_01205_),
    .A2(_06151_),
    .B1(_01192_),
    .C1(_01868_),
    .X(_06182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _13986_ (.A1(_01297_),
    .A2(_01296_),
    .A3(_06150_),
    .B1(_01191_),
    .B2(_06182_),
    .X(_06183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13987_ (.A1_N(_01298_),
    .A2_N(_06183_),
    .B1(_01298_),
    .B2(_06183_),
    .X(_01957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _13988_ (.A1(_01230_),
    .A2(_06776_),
    .A3(_07816_),
    .B1(_01534_),
    .B2(_01216_),
    .X(_06184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _13989_ (.A1(_06758_),
    .A2(_01204_),
    .B1(_07821_),
    .B2(_06184_),
    .X(_06185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13990_ (.A(_07815_),
    .B(_06185_),
    .X(_06186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _13991_ (.A1(_01184_),
    .A2(_01190_),
    .B1(_07822_),
    .B2(_06113_),
    .C1(_06186_),
    .X(_06187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _13992_ (.A1_N(_07845_),
    .A2_N(_06187_),
    .B1(_07845_),
    .B2(_06187_),
    .X(_01958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13993_ (.A(\design_top.core0.REG1[8][31] ),
    .Y(_00833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13994_ (.A(_06115_),
    .B(_01962_),
    .X(_01963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _13995_ (.A(_06133_),
    .B(_01561_),
    .X(_01965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13996_ (.A(\design_top.core0.REG1[9][31] ),
    .Y(_00834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _13997_ (.A(_01968_),
    .B(_06134_),
    .C(_06135_),
    .X(_01969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _13998_ (.A(_05994_),
    .B(_01366_),
    .C(_01949_),
    .X(_01974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _13999_ (.A(\design_top.core0.REG1[7][31] ),
    .Y(_00831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a32o_2 _14000_ (.A1(_06760_),
    .A2(\design_top.core0.PC[6] ),
    .A3(_06179_),
    .B1(_06763_),
    .B2(\design_top.core0.PC[7] ),
    .X(_06188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31oi_2 _14001_ (.A1(_06166_),
    .A2(_06180_),
    .A3(_06164_),
    .B1(_06188_),
    .Y(_06189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14002_ (.A(\design_top.core0.PC[8] ),
    .Y(_06190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14003_ (.A1(_01360_),
    .A2(_06190_),
    .B1(_06750_),
    .B2(\design_top.core0.PC[8] ),
    .X(_06191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14004_ (.A1_N(_06189_),
    .A2_N(_06191_),
    .B1(_06189_),
    .B2(_06191_),
    .X(_01978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14005_ (.A(\design_top.core0.NXPC[9] ),
    .Y(_01980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14006_ (.A(_07839_),
    .Y(_06192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14007_ (.A(_06192_),
    .X(_01299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14008_ (.A1(_01298_),
    .A2(_06183_),
    .B1(_01956_),
    .X(_06193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14009_ (.A1_N(_01299_),
    .A2_N(_06193_),
    .B1(_01299_),
    .B2(_06193_),
    .X(_01981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14010_ (.A(_06749_),
    .B(_07837_),
    .Y(_01165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14011_ (.A1(_07837_),
    .A2(_07838_),
    .B1(_01165_),
    .X(_06194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14012_ (.A(_06798_),
    .X(_01171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14013_ (.A1(_07845_),
    .A2(_06187_),
    .B1(_01171_),
    .B2(_01177_),
    .X(_06195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14014_ (.A1_N(_06194_),
    .A2_N(_06195_),
    .B1(_06194_),
    .B2(_06195_),
    .X(_01982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14015_ (.A(_06114_),
    .X(_06196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14016_ (.A(_06196_),
    .B(_01986_),
    .X(_01987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14017_ (.A(_06133_),
    .B(_01641_),
    .X(_01989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14018_ (.A(\design_top.core0.REG1[4][31] ),
    .Y(_00828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14019_ (.A(\design_top.core0.REG1[5][31] ),
    .Y(_00829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14020_ (.A(\design_top.core0.REG1[6][31] ),
    .Y(_00830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14021_ (.A(_01992_),
    .B(_06134_),
    .C(_06135_),
    .X(_01993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14022_ (.A(_06748_),
    .Y(_01359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14023_ (.A(\design_top.core0.PC[9] ),
    .Y(_06197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14024_ (.A(_01359_),
    .B(_06197_),
    .Y(_06198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _14025_ (.A1(_01359_),
    .A2(_06197_),
    .B1(_06198_),
    .Y(_06199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _14026_ (.A1(_01360_),
    .A2(_06190_),
    .B1(_06189_),
    .B2(_06191_),
    .Y(_06200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14027_ (.A1_N(_06199_),
    .A2_N(_06200_),
    .B1(_06199_),
    .B2(_06200_),
    .X(_02001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14028_ (.A(\design_top.core0.NXPC[10] ),
    .Y(_02003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14029_ (.A(_07841_),
    .X(_01300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14030_ (.A1(_01299_),
    .A2(_06193_),
    .B1(_01165_),
    .X(_06201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14031_ (.A1_N(_01300_),
    .A2_N(_06201_),
    .B1(_01300_),
    .B2(_06201_),
    .X(_02005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14032_ (.A(_07838_),
    .Y(_01156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14033_ (.A1(_07837_),
    .A2(_01156_),
    .B1(_06194_),
    .B2(_06195_),
    .X(_06202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14034_ (.A1_N(_07842_),
    .A2_N(_06202_),
    .B1(_07842_),
    .B2(_06202_),
    .X(_02006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14035_ (.A(\design_top.core0.REG1[2][31] ),
    .Y(_00825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14036_ (.A(_06196_),
    .B(_02010_),
    .X(_02011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14037_ (.A(_06035_),
    .X(_06203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14038_ (.A(_06203_),
    .B(_01695_),
    .X(_02013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14039_ (.A(\design_top.core0.REG1[1][31] ),
    .Y(_00824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14040_ (.A(\design_top.core0.REG1[3][31] ),
    .Y(_00826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14041_ (.A(_06029_),
    .X(_06204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14042_ (.A(_06031_),
    .X(_06205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14043_ (.A(_02016_),
    .B(_06204_),
    .C(_06205_),
    .X(_02017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14044_ (.A(_06741_),
    .X(_01358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14045_ (.A(\design_top.core0.PC[10] ),
    .Y(_06206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14046_ (.A1(_01358_),
    .A2(_06206_),
    .B1(\design_top.core0.SIMM[10] ),
    .B2(\design_top.core0.PC[10] ),
    .X(_06207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _14047_ (.A1(_06748_),
    .A2(\design_top.core0.PC[9] ),
    .B1(_06198_),
    .B2(_06200_),
    .Y(_06208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14048_ (.A1_N(_06207_),
    .A2_N(_06208_),
    .B1(_06207_),
    .B2(_06208_),
    .X(_02025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14049_ (.A(\design_top.core0.NXPC[11] ),
    .Y(_02027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14050_ (.A(_07843_),
    .Y(_01301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14051_ (.A1(_01300_),
    .A2(_06201_),
    .B1(_02004_),
    .X(_06209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14052_ (.A1_N(_01301_),
    .A2_N(_06209_),
    .B1(_01301_),
    .B2(_06209_),
    .X(_02028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14053_ (.A1(_07842_),
    .A2(_06202_),
    .B1(_01142_),
    .B2(_01148_),
    .X(_06210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14054_ (.A(_06210_),
    .Y(_06211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14055_ (.A1(_01301_),
    .A2(_06210_),
    .B1(_07843_),
    .B2(_06211_),
    .X(_02029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14056_ (.A(_07764_),
    .B(_06663_),
    .Y(_00821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14057_ (.A(_06196_),
    .B(_02033_),
    .X(_02034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14058_ (.A(_06203_),
    .B(_01748_),
    .X(_02036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14059_ (.A(_02039_),
    .B(_06204_),
    .C(_06205_),
    .X(_02040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14060_ (.A(\design_top.core0.PC[11] ),
    .Y(_06212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14061_ (.A1(_01357_),
    .A2(_06212_),
    .B1(\design_top.core0.SIMM[11] ),
    .B2(\design_top.core0.PC[11] ),
    .X(_06213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14062_ (.A1(_01358_),
    .A2(_06206_),
    .B1(_06207_),
    .B2(_06208_),
    .X(_06214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14063_ (.A1_N(_06213_),
    .A2_N(_06214_),
    .B1(_06213_),
    .B2(_06214_),
    .X(_02048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14064_ (.A(\design_top.core0.NXPC[12] ),
    .Y(_02050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14065_ (.A(_07829_),
    .X(_01302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14066_ (.A(_06754_),
    .B(_01134_),
    .Y(_01136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _14067_ (.A(_01298_),
    .B(_01301_),
    .C(_01300_),
    .D(_01299_),
    .X(_06215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14068_ (.A(_07840_),
    .B(_01148_),
    .Y(_01149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _14069_ (.A1(_06192_),
    .A2(_01956_),
    .B1(_02004_),
    .C1(_01165_),
    .X(_06216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _14070_ (.A1(_01149_),
    .A2(_01135_),
    .A3(_06216_),
    .B1(_01136_),
    .X(_06217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14071_ (.A1(_06183_),
    .A2(_06215_),
    .B1(_06217_),
    .Y(_06218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14072_ (.A(_06218_),
    .Y(_06219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14073_ (.A1(_07830_),
    .A2(_06218_),
    .B1(_01302_),
    .B2(_06219_),
    .X(_02052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _14074_ (.A1(_01171_),
    .A2(_01177_),
    .A3(_06194_),
    .B1(_07837_),
    .B2(_01156_),
    .X(_06220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14075_ (.A1(_01142_),
    .A2(_01148_),
    .B1(_07842_),
    .B2(_06220_),
    .X(_06221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14076_ (.A(_07846_),
    .B(_06194_),
    .C(_06187_),
    .X(_06222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14077_ (.A1(_01540_),
    .A2(_01134_),
    .B1(_07843_),
    .B2(_06221_),
    .C1(_06222_),
    .X(_06223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14078_ (.A(_06724_),
    .X(_06224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14079_ (.A1_N(_06224_),
    .A2_N(_01285_),
    .B1(_06224_),
    .B2(_01285_),
    .X(_06225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14080_ (.A(_06223_),
    .B(_06225_),
    .X(_06226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14081_ (.A(_06226_),
    .Y(_06227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _14082_ (.A1(_06223_),
    .A2(_06225_),
    .B1(_06227_),
    .X(_02053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14083_ (.A(_06196_),
    .B(_02057_),
    .X(_02058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14084_ (.A(_06203_),
    .B(_01792_),
    .X(_02060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14085_ (.A(_02063_),
    .B(_06204_),
    .C(_06205_),
    .X(_02064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14086_ (.A(\design_top.core0.PC[12] ),
    .Y(_06228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14087_ (.A1(_01356_),
    .A2(_06228_),
    .B1(_06725_),
    .B2(\design_top.core0.PC[12] ),
    .X(_06229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14088_ (.A(_06207_),
    .B(_06213_),
    .X(_06230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4b_2 _14089_ (.A(_06191_),
    .B(_06189_),
    .C(_06230_),
    .D_N(_06199_),
    .X(_06231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _14090_ (.A1(_06750_),
    .A2(\design_top.core0.PC[8] ),
    .B1(_06198_),
    .X(_06232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14091_ (.A1(_06748_),
    .A2(\design_top.core0.PC[9] ),
    .B1(_06232_),
    .Y(_06233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _14092_ (.A1(_01357_),
    .A2(_06212_),
    .B1(_01358_),
    .C1(_06206_),
    .X(_06234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14093_ (.A1(_01357_),
    .A2(_06212_),
    .B1(_06233_),
    .B2(_06230_),
    .C1(_06234_),
    .X(_06235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _14094_ (.A(_06231_),
    .B(_06235_),
    .X(_06236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14095_ (.A1_N(_06229_),
    .A2_N(_06236_),
    .B1(_06229_),
    .B2(_06236_),
    .X(_02072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14096_ (.A(\design_top.core0.NXPC[13] ),
    .Y(_02074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14097_ (.A(_07831_),
    .Y(_01303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14098_ (.A1(_01302_),
    .A2(_06219_),
    .B1(_02051_),
    .X(_06237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14099_ (.A1_N(_01303_),
    .A2_N(_06237_),
    .B1(_01303_),
    .B2(_06237_),
    .X(_02075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14100_ (.A(_06729_),
    .X(_01102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14101_ (.A(_06805_),
    .X(_06238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14102_ (.A(_01284_),
    .Y(_06239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14103_ (.A1(_01102_),
    .A2(_01284_),
    .B1(_06238_),
    .B2(_06239_),
    .X(_06240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14104_ (.A(_06224_),
    .X(_01116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14105_ (.A1(_01116_),
    .A2(_01285_),
    .B1(_06226_),
    .Y(_06241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14106_ (.A1_N(_06240_),
    .A2_N(_06241_),
    .B1(_06240_),
    .B2(_06241_),
    .X(_02076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14107_ (.A(_06196_),
    .B(_02080_),
    .X(_02081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14108_ (.A(_06203_),
    .B(_01835_),
    .X(_02083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14109_ (.A(_02086_),
    .B(_06204_),
    .C(_06205_),
    .X(_02087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14110_ (.A(\design_top.core0.PC[13] ),
    .Y(_06242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14111_ (.A(_06730_),
    .B(\design_top.core0.PC[13] ),
    .X(_06243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14112_ (.A1(_01355_),
    .A2(_06242_),
    .B1(_06243_),
    .X(_06244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _14113_ (.A1(_01356_),
    .A2(_06228_),
    .B1(_06229_),
    .B2(_06236_),
    .Y(_06245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14114_ (.A1_N(_06244_),
    .A2_N(_06245_),
    .B1(_06244_),
    .B2(_06245_),
    .X(_02095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14115_ (.A(_02096_),
    .B(_08076_),
    .Y(_02097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor3_2 _14116_ (.A(\design_top.core0.RESMODE[0] ),
    .B(_06023_),
    .C(_01331_),
    .Y(_02098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14117_ (.A(\design_top.core0.NXPC[14] ),
    .Y(_02099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14118_ (.A(_07834_),
    .X(_01304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14119_ (.A(_06238_),
    .B(_01108_),
    .Y(_01110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _14120_ (.A1(_02051_),
    .A2(_01110_),
    .B1(_01109_),
    .X(_06246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _14121_ (.A1(_01302_),
    .A2(_01303_),
    .A3(_06219_),
    .B1(_06246_),
    .X(_06247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14122_ (.A1_N(_01304_),
    .A2_N(_06247_),
    .B1(_01304_),
    .B2(_06247_),
    .X(_02101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14123_ (.A(_06734_),
    .X(_06248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14124_ (.A1_N(_06248_),
    .A2_N(_01283_),
    .B1(_06248_),
    .B2(_01283_),
    .X(_06249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14125_ (.A1_N(_06724_),
    .A2_N(_01285_),
    .B1(_06238_),
    .B2(_06239_),
    .X(_06250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _14126_ (.A1(_06238_),
    .A2(_06239_),
    .B1(_06227_),
    .B2(_06250_),
    .Y(_06251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14127_ (.A1_N(_06249_),
    .A2_N(_06251_),
    .B1(_06249_),
    .B2(_06251_),
    .X(_02102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14128_ (.A(_06721_),
    .X(_01006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14129_ (.A(_06037_),
    .X(_06252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14130_ (.A(_06252_),
    .B(_02106_),
    .X(_02107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14131_ (.A(_06203_),
    .B(_01880_),
    .X(_02109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14132_ (.A(_02112_),
    .B(_06204_),
    .C(_06205_),
    .X(_02113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14133_ (.A(_06810_),
    .X(_01075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14134_ (.A(_06733_),
    .X(_01354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14135_ (.A(\design_top.core0.PC[14] ),
    .Y(_06253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14136_ (.A1(_01354_),
    .A2(_06253_),
    .B1(\design_top.core0.SIMM[14] ),
    .B2(\design_top.core0.PC[14] ),
    .X(_06254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14137_ (.A(_01355_),
    .B(_06242_),
    .Y(_06255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14138_ (.A1(_06255_),
    .A2(_06245_),
    .B1(_06243_),
    .Y(_06256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14139_ (.A1_N(_06254_),
    .A2_N(_06256_),
    .B1(_06254_),
    .B2(_06256_),
    .X(_02121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14140_ (.A(\design_top.core0.NXPC[15] ),
    .Y(_02123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14141_ (.A1(_01304_),
    .A2(_06247_),
    .B1(_02100_),
    .X(_06257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14142_ (.A1_N(_01305_),
    .A2_N(_06257_),
    .B1(_01305_),
    .B2(_06257_),
    .X(_02124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14143_ (.A(_01282_),
    .Y(_06258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14144_ (.A(_06809_),
    .B(_06258_),
    .Y(_06259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _14145_ (.A1(_06809_),
    .A2(_06258_),
    .B1(_06259_),
    .Y(_06260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14146_ (.A(_06248_),
    .X(_01089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _14147_ (.A1(_01089_),
    .A2(_01283_),
    .B1(_06249_),
    .B2(_06251_),
    .Y(_06261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14148_ (.A1_N(_06260_),
    .A2_N(_06261_),
    .B1(_06260_),
    .B2(_06261_),
    .X(_02125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14149_ (.A(_06252_),
    .B(_02129_),
    .X(_02130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14150_ (.A(_06035_),
    .B(_01924_),
    .X(_02132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14151_ (.A(_06028_),
    .X(_06262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14152_ (.A(_06030_),
    .X(_06263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14153_ (.A(_02134_),
    .B(_06262_),
    .C(_06263_),
    .X(_02135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14154_ (.A(_06808_),
    .B(\design_top.core0.PC[15] ),
    .Y(_06264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _14155_ (.A1(_06808_),
    .A2(\design_top.core0.PC[15] ),
    .B1(_06264_),
    .X(_06265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14156_ (.A1(_01354_),
    .A2(_06253_),
    .B1(_06254_),
    .B2(_06256_),
    .X(_06266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14157_ (.A1_N(_06265_),
    .A2_N(_06266_),
    .B1(_06265_),
    .B2(_06266_),
    .X(_02143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14158_ (.A(\design_top.core0.NXPC[16] ),
    .Y(_02145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _14159_ (.A(_01302_),
    .B(_01303_),
    .C(_01305_),
    .D(_01304_),
    .X(_06267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14160_ (.A(_07832_),
    .Y(_01082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14161_ (.A(_01088_),
    .B(_01095_),
    .Y(_01096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _14162_ (.A1(_02100_),
    .A2(_06246_),
    .B1(_01082_),
    .C1(_01096_),
    .X(_06268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _14163_ (.A1(_06217_),
    .A2(_06267_),
    .B1(_01083_),
    .C1(_06268_),
    .X(_06269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _14164_ (.A1(_06215_),
    .A2(_06267_),
    .A3(_06183_),
    .B1(_06269_),
    .X(_06270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14165_ (.A(_06270_),
    .Y(_06271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14166_ (.A1(_07854_),
    .A2(_06271_),
    .B1(_01306_),
    .B2(_06270_),
    .X(_02147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14167_ (.A1(_06248_),
    .A2(_01283_),
    .B1(_06810_),
    .B2(_01282_),
    .X(_06272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4bb_2 _14168_ (.A(_06249_),
    .B(_06225_),
    .C_N(_06260_),
    .D_N(_06240_),
    .X(_06273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14169_ (.A1(_06238_),
    .A2(_06239_),
    .B1(_06250_),
    .Y(_06274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _14170_ (.A(_06249_),
    .B(_06274_),
    .C_N(_06260_),
    .X(_06275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14171_ (.A1(_06259_),
    .A2(_06272_),
    .B1(_06223_),
    .B2(_06273_),
    .C1(_06275_),
    .X(_06276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14172_ (.A1_N(_06815_),
    .A2_N(_01281_),
    .B1(_06815_),
    .B2(_01281_),
    .X(_06277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14173_ (.A(_06276_),
    .B(_06277_),
    .X(_06278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14174_ (.A(_06278_),
    .Y(_06279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _14175_ (.A1(_06276_),
    .A2(_06277_),
    .B1(_06279_),
    .X(_02148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14176_ (.A(_06252_),
    .B(_01562_),
    .X(_02154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14177_ (.A(_02157_),
    .B(_06262_),
    .C(_06263_),
    .X(_02158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14178_ (.A(_05994_),
    .B(_05981_),
    .C(_02138_),
    .X(_02161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4b_2 _14179_ (.A(_06229_),
    .B(_06265_),
    .C(_06254_),
    .D_N(_06244_),
    .X(_06280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14180_ (.A(_06808_),
    .B(\design_top.core0.PC[15] ),
    .Y(_06281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31o_2 _14181_ (.A1(_06725_),
    .A2(\design_top.core0.PC[12] ),
    .A3(_06243_),
    .B1(_06255_),
    .X(_06282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _14182_ (.A(_06254_),
    .B(_06265_),
    .C_N(_06282_),
    .X(_06283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o311a_2 _14183_ (.A1(_01354_),
    .A2(_06253_),
    .A3(_06264_),
    .B1(_06281_),
    .C1(_06283_),
    .X(_06284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14184_ (.A1(_06235_),
    .A2(_06280_),
    .B1(_06231_),
    .B2(_06280_),
    .C1(_06284_),
    .X(_06285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14185_ (.A(\design_top.core0.PC[16] ),
    .Y(_06286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14186_ (.A1(_01352_),
    .A2(_06286_),
    .B1(_06717_),
    .B2(\design_top.core0.PC[16] ),
    .X(_06287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14187_ (.A1_N(_06285_),
    .A2_N(_06287_),
    .B1(_06285_),
    .B2(_06287_),
    .X(_02166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14188_ (.A(\design_top.core0.NXPC[17] ),
    .Y(_02168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14189_ (.A(_07855_),
    .Y(_01307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14190_ (.A1(_01306_),
    .A2(_06270_),
    .B1(_02146_),
    .X(_06288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14191_ (.A1_N(_01307_),
    .A2_N(_06288_),
    .B1(_01307_),
    .B2(_06288_),
    .X(_02169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14192_ (.A(_01048_),
    .X(_06289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14193_ (.A(_06716_),
    .X(_06290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14194_ (.A(_01280_),
    .Y(_06291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14195_ (.A1(_06289_),
    .A2(_01280_),
    .B1(_06290_),
    .B2(_06291_),
    .X(_06292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14196_ (.A1(_01062_),
    .A2(_01281_),
    .B1(_06278_),
    .Y(_06293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14197_ (.A1_N(_06292_),
    .A2_N(_06293_),
    .B1(_06292_),
    .B2(_06293_),
    .X(_02170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14198_ (.A(_06252_),
    .B(_01642_),
    .X(_02176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14199_ (.A(_02179_),
    .B(_06262_),
    .C(_06263_),
    .X(_02180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14200_ (.A(\design_top.core0.PC[17] ),
    .Y(_06294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14201_ (.A(_01351_),
    .B(_06294_),
    .Y(_06295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _14202_ (.A1(_01351_),
    .A2(_06294_),
    .B1(_06295_),
    .Y(_06296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _14203_ (.A1(_01352_),
    .A2(_06286_),
    .B1(_06285_),
    .B2(_06287_),
    .Y(_06297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14204_ (.A1_N(_06296_),
    .A2_N(_06297_),
    .B1(_06296_),
    .B2(_06297_),
    .X(_02187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14205_ (.A(\design_top.core0.NXPC[18] ),
    .Y(_02189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14206_ (.A(_07849_),
    .X(_01308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14207_ (.A(_06290_),
    .B(_01054_),
    .Y(_01056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _14208_ (.A1(_02146_),
    .A2(_01056_),
    .B1(_01055_),
    .Y(_06298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a31oi_2 _14209_ (.A1(_07854_),
    .A2(_07855_),
    .A3(_06271_),
    .B1(_06298_),
    .Y(_06299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14210_ (.A1_N(_01308_),
    .A2_N(_06299_),
    .B1(_01308_),
    .B2(_06299_),
    .X(_02191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14211_ (.A(_06711_),
    .X(_06300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14212_ (.A1_N(_06300_),
    .A2_N(_01279_),
    .B1(_06711_),
    .B2(_01279_),
    .X(_06301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14213_ (.A1_N(_06815_),
    .A2_N(_01281_),
    .B1(_06290_),
    .B2(_06291_),
    .X(_06302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _14214_ (.A1(_06290_),
    .A2(_06291_),
    .B1(_06279_),
    .B2(_06302_),
    .Y(_06303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14215_ (.A1_N(_06301_),
    .A2_N(_06303_),
    .B1(_06301_),
    .B2(_06303_),
    .X(_02192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14216_ (.A(_06252_),
    .B(_01696_),
    .X(_02198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14217_ (.A(_02201_),
    .B(_06262_),
    .C(_06263_),
    .X(_02202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14218_ (.A(_06710_),
    .X(_01350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14219_ (.A(\design_top.core0.PC[18] ),
    .Y(_06304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14220_ (.A1(\design_top.core0.SIMM[18] ),
    .A2(\design_top.core0.PC[18] ),
    .B1(_01350_),
    .B2(_06304_),
    .X(_06305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14221_ (.A(_06305_),
    .Y(_06306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _14222_ (.A1(_06714_),
    .A2(\design_top.core0.PC[17] ),
    .B1(_06295_),
    .B2(_06297_),
    .Y(_06307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14223_ (.A1_N(_06306_),
    .A2_N(_06307_),
    .B1(_06306_),
    .B2(_06307_),
    .X(_02209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14224_ (.A(\design_top.core0.NXPC[19] ),
    .Y(_02211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14225_ (.A1(_01308_),
    .A2(_06299_),
    .B1(_02190_),
    .X(_06308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14226_ (.A1_N(_01309_),
    .A2_N(_06308_),
    .B1(_01309_),
    .B2(_06308_),
    .X(_02212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14227_ (.A(_01278_),
    .Y(_06309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14228_ (.A(_07851_),
    .B(_06309_),
    .Y(_06310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _14229_ (.A1(_07851_),
    .A2(_06309_),
    .B1(_06310_),
    .Y(_06311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14230_ (.A(_06300_),
    .X(_01020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _14231_ (.A1(_01020_),
    .A2(_01279_),
    .B1(_06301_),
    .B2(_06303_),
    .Y(_06312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14232_ (.A1_N(_06311_),
    .A2_N(_06312_),
    .B1(_06311_),
    .B2(_06312_),
    .X(_02213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14233_ (.A(_06037_),
    .X(_06313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14234_ (.A(_06313_),
    .B(_01749_),
    .X(_02219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14235_ (.A(_02222_),
    .B(_06262_),
    .C(_06263_),
    .X(_02223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14236_ (.A(_00945_),
    .B(_06686_),
    .Y(_00946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14237_ (.A(\design_top.core0.PC[19] ),
    .Y(_06314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14238_ (.A1(\design_top.core0.SIMM[19] ),
    .A2(\design_top.core0.PC[19] ),
    .B1(_01349_),
    .B2(_06314_),
    .X(_06315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14239_ (.A(_06315_),
    .Y(_06316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14240_ (.A1(_01350_),
    .A2(_06304_),
    .B1(_06306_),
    .B2(_06307_),
    .X(_06317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14241_ (.A1_N(_06316_),
    .A2_N(_06317_),
    .B1(_06316_),
    .B2(_06317_),
    .X(_02230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14242_ (.A(\design_top.core0.NXPC[20] ),
    .Y(_02232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14243_ (.A(_07872_),
    .X(_01310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _14244_ (.A(_01306_),
    .B(_01307_),
    .C(_01308_),
    .D(_01309_),
    .X(_06318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14245_ (.A(_07852_),
    .Y(_01013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14246_ (.A(_07848_),
    .B(_06298_),
    .Y(_06319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _14247_ (.A1(_01027_),
    .A2(_01013_),
    .A3(_06319_),
    .B1(_01014_),
    .X(_06320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14248_ (.A1(_06270_),
    .A2(_06318_),
    .B1(_06320_),
    .Y(_06321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14249_ (.A(_06321_),
    .Y(_06322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14250_ (.A1(_07873_),
    .A2(_06321_),
    .B1(_01310_),
    .B2(_06322_),
    .X(_02234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14251_ (.A(_06689_),
    .X(_06323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14252_ (.A1_N(_06323_),
    .A2_N(_01277_),
    .B1(_06689_),
    .B2(_01277_),
    .X(_06324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14253_ (.A1(_06300_),
    .A2(_01279_),
    .B1(_01006_),
    .B2(_01278_),
    .X(_06325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4bb_2 _14254_ (.A(_06301_),
    .B(_06277_),
    .C_N(_06311_),
    .D_N(_06292_),
    .X(_06326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14255_ (.A1(_06290_),
    .A2(_06291_),
    .B1(_06302_),
    .Y(_06327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _14256_ (.A(_06301_),
    .B(_06327_),
    .C_N(_06311_),
    .X(_06328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14257_ (.A1(_06310_),
    .A2(_06325_),
    .B1(_06276_),
    .B2(_06326_),
    .C1(_06328_),
    .X(_06329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14258_ (.A(_06324_),
    .B(_06329_),
    .X(_06330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14259_ (.A1(_06324_),
    .A2(_06329_),
    .B1_N(_06330_),
    .X(_02235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14260_ (.A(_06313_),
    .B(_01793_),
    .X(_02241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14261_ (.A(_06827_),
    .X(_06331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14262_ (.A(_06331_),
    .X(_00939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14263_ (.A(_06028_),
    .X(_06332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14264_ (.A(_06030_),
    .X(_06333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14265_ (.A(_02244_),
    .B(_06332_),
    .C(_06333_),
    .X(_02245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14266_ (.A(\design_top.core0.PC[20] ),
    .Y(_06334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14267_ (.A1(_01348_),
    .A2(_06334_),
    .B1(_06690_),
    .B2(\design_top.core0.PC[20] ),
    .X(_06335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4b_2 _14268_ (.A(_06287_),
    .B(_06316_),
    .C(_06306_),
    .D_N(_06296_),
    .X(_06336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _14269_ (.A1(_01349_),
    .A2(_06314_),
    .B1(_01350_),
    .C1(_06304_),
    .X(_06337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _14270_ (.A1(_06717_),
    .A2(\design_top.core0.PC[16] ),
    .B1(_06295_),
    .X(_06338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2111ai_2 _14271_ (.A1(_06714_),
    .A2(\design_top.core0.PC[17] ),
    .B1(_06338_),
    .C1(_06305_),
    .D1(_06315_),
    .Y(_06339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _14272_ (.A1(_01349_),
    .A2(_06314_),
    .B1(_06337_),
    .C1(_06339_),
    .X(_06340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14273_ (.A1(_06285_),
    .A2(_06336_),
    .B1(_06340_),
    .X(_06341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14274_ (.A1_N(_06335_),
    .A2_N(_06341_),
    .B1(_06335_),
    .B2(_06341_),
    .X(_02252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14275_ (.A(\design_top.core0.NXPC[21] ),
    .Y(_02254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14276_ (.A(_07871_),
    .Y(_01311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14277_ (.A1(_01310_),
    .A2(_06322_),
    .B1(_02233_),
    .X(_06342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14278_ (.A1_N(_01311_),
    .A2_N(_06342_),
    .B1(_01311_),
    .B2(_06342_),
    .X(_02255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14279_ (.A(_06694_),
    .X(_06343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14280_ (.A1_N(_06343_),
    .A2_N(_01276_),
    .B1(_06343_),
    .B2(_01276_),
    .X(_06344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14281_ (.A(_06323_),
    .X(_00993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14282_ (.A1(_00993_),
    .A2(_01277_),
    .B1(_06330_),
    .Y(_06345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14283_ (.A1_N(_06344_),
    .A2_N(_06345_),
    .B1(_06344_),
    .B2(_06345_),
    .X(_02256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14284_ (.A(_06313_),
    .B(_01836_),
    .X(_02262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14285_ (.A(_02265_),
    .B(_06332_),
    .C(_06333_),
    .X(_02266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14286_ (.A(\design_top.core0.PC[21] ),
    .Y(_06346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14287_ (.A(_01347_),
    .B(_06346_),
    .Y(_06347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _14288_ (.A1(_01347_),
    .A2(_06346_),
    .B1(_06347_),
    .Y(_06348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _14289_ (.A1(_01348_),
    .A2(_06334_),
    .B1(_06335_),
    .B2(_06341_),
    .Y(_06349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14290_ (.A1_N(_06348_),
    .A2_N(_06349_),
    .B1(_06348_),
    .B2(_06349_),
    .X(_02273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14291_ (.A(\design_top.core0.NXPC[22] ),
    .Y(_02275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14292_ (.A(_07874_),
    .X(_01312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14293_ (.A(_06821_),
    .B(_00985_),
    .Y(_00987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _14294_ (.A1(_00987_),
    .A2(_02233_),
    .B1(_00986_),
    .X(_06350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _14295_ (.A1(_01311_),
    .A2(_01310_),
    .A3(_06322_),
    .B1(_06350_),
    .X(_06351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14296_ (.A1_N(_01312_),
    .A2_N(_06351_),
    .B1(_01312_),
    .B2(_06351_),
    .X(_02277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14297_ (.A(_06698_),
    .X(_06352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14298_ (.A1_N(_06352_),
    .A2_N(_01275_),
    .B1(_06352_),
    .B2(_01275_),
    .X(_06353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14299_ (.A(_06694_),
    .X(_00979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14300_ (.A1(_06323_),
    .A2(_01277_),
    .B1(_06343_),
    .B2(_01276_),
    .X(_06354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14301_ (.A1(_00979_),
    .A2(_01276_),
    .B1(_06330_),
    .B2(_06354_),
    .X(_06355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14302_ (.A1_N(_06353_),
    .A2_N(_06355_),
    .B1(_06353_),
    .B2(_06355_),
    .X(_02278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14303_ (.A(_06313_),
    .B(_01881_),
    .X(_02284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14304_ (.A(_02287_),
    .B(_06332_),
    .C(_06333_),
    .X(_02288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14305_ (.A(\design_top.core0.PC[22] ),
    .Y(_06356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14306_ (.A1(_01346_),
    .A2(_06356_),
    .B1(_06699_),
    .B2(\design_top.core0.PC[22] ),
    .X(_06357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _14307_ (.A1(_06820_),
    .A2(\design_top.core0.PC[21] ),
    .B1(_06347_),
    .B2(_06349_),
    .Y(_06358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14308_ (.A1_N(_06357_),
    .A2_N(_06358_),
    .B1(_06357_),
    .B2(_06358_),
    .X(_02295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14309_ (.A(\design_top.core0.NXPC[23] ),
    .Y(_02297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14310_ (.A1(_01312_),
    .A2(_06351_),
    .B1(_02276_),
    .X(_06359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14311_ (.A1_N(_01313_),
    .A2_N(_06359_),
    .B1(_01313_),
    .B2(_06359_),
    .X(_02298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14312_ (.A(_06702_),
    .X(_06360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14313_ (.A(_01274_),
    .Y(_06361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14314_ (.A(_06360_),
    .B(_06361_),
    .Y(_06362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _14315_ (.A1(_06360_),
    .A2(_06361_),
    .B1(_06362_),
    .Y(_06363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14316_ (.A(_06352_),
    .X(_00966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _14317_ (.A1(_00966_),
    .A2(_01275_),
    .B1(_06353_),
    .B2(_06355_),
    .Y(_06364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14318_ (.A1_N(_06363_),
    .A2_N(_06364_),
    .B1(_06363_),
    .B2(_06364_),
    .X(_02299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14319_ (.A(_06313_),
    .B(_01925_),
    .X(_02305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14320_ (.A(_02308_),
    .B(_06332_),
    .C(_06333_),
    .X(_02309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14321_ (.A1_N(_07743_),
    .A2_N(\design_top.core0.PC[23] ),
    .B1(_07743_),
    .B2(\design_top.core0.PC[23] ),
    .X(_06365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14322_ (.A1(_01346_),
    .A2(_06356_),
    .B1(_06357_),
    .B2(_06358_),
    .X(_06366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14323_ (.A1_N(_06365_),
    .A2_N(_06366_),
    .B1(_06365_),
    .B2(_06366_),
    .X(_02316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14324_ (.A(\design_top.core0.NXPC[24] ),
    .Y(_02318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14325_ (.A(_07862_),
    .X(_01314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _14326_ (.A(_01311_),
    .B(_01310_),
    .C(_01313_),
    .D(_01312_),
    .X(_06367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14327_ (.A(_07869_),
    .Y(_00959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14328_ (.A(_00965_),
    .B(_00972_),
    .Y(_00973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _14329_ (.A1(_02276_),
    .A2(_06350_),
    .B1(_00959_),
    .C1(_00973_),
    .X(_06368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _14330_ (.A1(_06320_),
    .A2(_06367_),
    .B1(_00960_),
    .C1(_06368_),
    .X(_06369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _14331_ (.A1(_06318_),
    .A2(_06367_),
    .A3(_06270_),
    .B1(_06369_),
    .X(_06370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14332_ (.A1_N(_01314_),
    .A2_N(_06370_),
    .B1(_01314_),
    .B2(_06370_),
    .X(_02320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14333_ (.A1_N(_06331_),
    .A2_N(_01273_),
    .B1(_06331_),
    .B2(_01273_),
    .X(_06371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14334_ (.A1(_06352_),
    .A2(_01275_),
    .B1(_00952_),
    .B2(_01274_),
    .X(_06372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14335_ (.A(_06363_),
    .Y(_06373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4b_2 _14336_ (.A(_06353_),
    .B(_06373_),
    .C(_06324_),
    .D_N(_06344_),
    .X(_06374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2111o_2 _14337_ (.A1(_00979_),
    .A2(_01276_),
    .B1(_06354_),
    .C1(_06353_),
    .D1(_06373_),
    .X(_06375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14338_ (.A1(_06362_),
    .A2(_06372_),
    .B1(_06329_),
    .B2(_06374_),
    .C1(_06375_),
    .X(_06376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14339_ (.A(_06371_),
    .B(_06376_),
    .X(_06377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14340_ (.A1(_06371_),
    .A2(_06376_),
    .B1_N(_06377_),
    .X(_02321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14341_ (.A(_06037_),
    .X(_06378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14342_ (.A(_06378_),
    .B(_01965_),
    .X(_02327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14343_ (.A(_02330_),
    .B(_06332_),
    .C(_06333_),
    .X(_02331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2b_2 _14344_ (.A(_06335_),
    .B_N(_06348_),
    .X(_06379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14345_ (.A(_06357_),
    .B(_06365_),
    .X(_06380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _14346_ (.A1(_06820_),
    .A2(\design_top.core0.PC[21] ),
    .B1(_06690_),
    .C1(\design_top.core0.PC[20] ),
    .X(_06381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14347_ (.A(_06340_),
    .B(_06379_),
    .Y(_06382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _14348_ (.A1(_06347_),
    .A2(_06381_),
    .A3(_06382_),
    .B1(_06699_),
    .B2(\design_top.core0.PC[22] ),
    .X(_06383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a221o_2 _14349_ (.A1(_06699_),
    .A2(\design_top.core0.PC[22] ),
    .B1(_07743_),
    .B2(\design_top.core0.PC[23] ),
    .C1(_06383_),
    .X(_06384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14350_ (.A1(_07743_),
    .A2(\design_top.core0.PC[23] ),
    .B1(_06384_),
    .Y(_06385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o41a_2 _14351_ (.A1(_06379_),
    .A2(_06380_),
    .A3(_06336_),
    .A4(_06285_),
    .B1(_06385_),
    .X(_06386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14352_ (.A(_06685_),
    .B(\design_top.core0.PC[24] ),
    .Y(_06387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14353_ (.A1(_06685_),
    .A2(\design_top.core0.PC[24] ),
    .B1(_06387_),
    .Y(_06388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14354_ (.A1_N(_06386_),
    .A2_N(_06388_),
    .B1(_06386_),
    .B2(_06388_),
    .X(_02338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14355_ (.A(\design_top.core0.NXPC[25] ),
    .Y(_02340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14356_ (.A(_07861_),
    .Y(_01315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14357_ (.A1(_01314_),
    .A2(_06370_),
    .B1(_02319_),
    .X(_06389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14358_ (.A1_N(_01315_),
    .A2_N(_06389_),
    .B1(_01315_),
    .B2(_06389_),
    .X(_02341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14359_ (.A(_06830_),
    .X(_06390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14360_ (.A1_N(_06390_),
    .A2_N(_01272_),
    .B1(_06390_),
    .B2(_01272_),
    .X(_06391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14361_ (.A1(_00939_),
    .A2(_01273_),
    .B1(_06377_),
    .Y(_06392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14362_ (.A1_N(_06391_),
    .A2_N(_06392_),
    .B1(_06391_),
    .B2(_06392_),
    .X(_02342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14363_ (.A(_06378_),
    .B(_01989_),
    .X(_02348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14364_ (.A(_06028_),
    .X(_06393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14365_ (.A(_06030_),
    .X(_06394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14366_ (.A(_02351_),
    .B(_06393_),
    .C(_06394_),
    .X(_02352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14367_ (.A(\design_top.core0.PC[25] ),
    .Y(_06395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14368_ (.A(_01343_),
    .B(_06395_),
    .X(_06396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14369_ (.A1(_06683_),
    .A2(\design_top.core0.PC[25] ),
    .B1(_06396_),
    .X(_06397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14370_ (.A1(_06386_),
    .A2(_06388_),
    .B1(_06387_),
    .Y(_06398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14371_ (.A1_N(_06397_),
    .A2_N(_06398_),
    .B1(_06397_),
    .B2(_06398_),
    .X(_02359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14372_ (.A(\design_top.core0.NXPC[26] ),
    .Y(_02361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14373_ (.A(_07859_),
    .X(_01316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14374_ (.A(_06684_),
    .B(_00931_),
    .Y(_00933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _14375_ (.A1(_02319_),
    .A2(_00933_),
    .B1(_00932_),
    .X(_06399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _14376_ (.A1(_01314_),
    .A2(_01315_),
    .A3(_06370_),
    .B1(_06399_),
    .X(_06400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14377_ (.A1_N(_01316_),
    .A2_N(_06400_),
    .B1(_01316_),
    .B2(_06400_),
    .X(_02363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14378_ (.A(_06678_),
    .X(_06401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14379_ (.A1_N(_06401_),
    .A2_N(_01271_),
    .B1(_06401_),
    .B2(_01271_),
    .X(_06402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14380_ (.A(_06390_),
    .X(_00925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14381_ (.A1(_06331_),
    .A2(_01273_),
    .B1(_06390_),
    .B2(_01272_),
    .X(_06403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14382_ (.A1(_00925_),
    .A2(_01272_),
    .B1(_06377_),
    .B2(_06403_),
    .X(_06404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14383_ (.A1_N(_06402_),
    .A2_N(_06404_),
    .B1(_06402_),
    .B2(_06404_),
    .X(_02364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14384_ (.A(_06378_),
    .B(_02013_),
    .X(_02370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14385_ (.A(_02373_),
    .B(_06393_),
    .C(_06394_),
    .X(_02374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14386_ (.A(_06677_),
    .X(_01342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14387_ (.A(\design_top.core0.PC[26] ),
    .Y(_06405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14388_ (.A1(_01342_),
    .A2(_06405_),
    .B1(\design_top.core0.SIMM[26] ),
    .B2(\design_top.core0.PC[26] ),
    .X(_06406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14389_ (.A(_06398_),
    .Y(_06407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14390_ (.A1(_01343_),
    .A2(_06395_),
    .B1(_06396_),
    .B2(_06407_),
    .X(_06408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14391_ (.A1_N(_06406_),
    .A2_N(_06408_),
    .B1(_06406_),
    .B2(_06408_),
    .X(_02381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14392_ (.A(\design_top.core0.NXPC[27] ),
    .Y(_02383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14393_ (.A(_07858_),
    .Y(_01317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14394_ (.A1(_01316_),
    .A2(_06400_),
    .B1(_02362_),
    .X(_06409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14395_ (.A1_N(_01317_),
    .A2_N(_06409_),
    .B1(_01317_),
    .B2(_06409_),
    .X(_02384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14396_ (.A(_01270_),
    .Y(_06410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14397_ (.A(_07857_),
    .B(_06410_),
    .Y(_06411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _14398_ (.A1(_07857_),
    .A2(_06410_),
    .B1(_06411_),
    .Y(_06412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14399_ (.A(_06401_),
    .X(_00912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _14400_ (.A1(_00912_),
    .A2(_01271_),
    .B1(_06402_),
    .B2(_06404_),
    .Y(_06413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14401_ (.A1_N(_06412_),
    .A2_N(_06413_),
    .B1(_06412_),
    .B2(_06413_),
    .X(_02385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14402_ (.A(_06378_),
    .B(_02036_),
    .X(_02391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14403_ (.A(_02394_),
    .B(_06393_),
    .C(_06394_),
    .X(_02395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14404_ (.A(\design_top.core0.PC[27] ),
    .Y(_06414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14405_ (.A1(_01341_),
    .A2(_06414_),
    .B1(\design_top.core0.SIMM[27] ),
    .B2(\design_top.core0.PC[27] ),
    .X(_06415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14406_ (.A1(_01342_),
    .A2(_06405_),
    .B1(_06406_),
    .B2(_06408_),
    .X(_06416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14407_ (.A1_N(_06415_),
    .A2_N(_06416_),
    .B1(_06415_),
    .B2(_06416_),
    .X(_02402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14408_ (.A(\design_top.core0.NXPC[28] ),
    .Y(_02404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14409_ (.A(_00884_),
    .B(_00891_),
    .Y(_02405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14410_ (.A(_07866_),
    .Y(_01318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14411_ (.A(_07857_),
    .B(_00904_),
    .Y(_00906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _14412_ (.A(_07862_),
    .B(_01315_),
    .C(_01317_),
    .D(_01316_),
    .X(_06417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14413_ (.A(_00911_),
    .B(_00918_),
    .Y(_00919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _14414_ (.A1(_00919_),
    .A2(_06399_),
    .B1(_00906_),
    .C1(_02362_),
    .X(_06418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14415_ (.A1(_06370_),
    .A2(_06417_),
    .B1(_00905_),
    .B2(_06418_),
    .X(_06419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14416_ (.A1_N(_01318_),
    .A2_N(_06419_),
    .B1(_01318_),
    .B2(_06419_),
    .X(_02406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14417_ (.A(_06834_),
    .X(_00898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14418_ (.A1(_00912_),
    .A2(_01271_),
    .B1(_00898_),
    .B2(_01270_),
    .X(_06420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14419_ (.A(_06412_),
    .Y(_06421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4b_2 _14420_ (.A(_06402_),
    .B(_06421_),
    .C(_06371_),
    .D_N(_06391_),
    .X(_06422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2111o_2 _14421_ (.A1(_00925_),
    .A2(_01272_),
    .B1(_06403_),
    .C1(_06402_),
    .D1(_06421_),
    .X(_06423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14422_ (.A1(_06411_),
    .A2(_06420_),
    .B1(_06376_),
    .B2(_06422_),
    .C1(_06423_),
    .X(_06424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14423_ (.A(_06424_),
    .Y(_06425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14424_ (.A(_06673_),
    .X(_06426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14425_ (.A(_06426_),
    .X(_00885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14426_ (.A1_N(_00885_),
    .A2_N(_01269_),
    .B1(_00885_),
    .B2(_01269_),
    .X(_06427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14427_ (.A(_06427_),
    .Y(_06428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14428_ (.A1(_06425_),
    .A2(_06428_),
    .B1(_06424_),
    .B2(_06427_),
    .X(_02407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14429_ (.A(_06378_),
    .B(_02060_),
    .X(_02413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14430_ (.A(_02416_),
    .B(_06393_),
    .C(_06394_),
    .X(_02417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a211o_2 _14431_ (.A1(_01341_),
    .A2(_06414_),
    .B1(_01342_),
    .C1(_06405_),
    .X(_06429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14432_ (.A(_06406_),
    .B(_06415_),
    .X(_06430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a221o_2 _14433_ (.A1(_01343_),
    .A2(_06395_),
    .B1(_06387_),
    .B2(_06396_),
    .C1(_06430_),
    .X(_06431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4b_2 _14434_ (.A(_06388_),
    .B(_06386_),
    .C(_06430_),
    .D_N(_06397_),
    .X(_06432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2111a_2 _14435_ (.A1(_01341_),
    .A2(_06414_),
    .B1(_06429_),
    .C1(_06431_),
    .D1(_06432_),
    .X(_06433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14436_ (.A(_06674_),
    .B(\design_top.core0.PC[28] ),
    .Y(_06434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _14437_ (.A1(_06674_),
    .A2(\design_top.core0.PC[28] ),
    .B1(_06434_),
    .X(_06435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14438_ (.A1_N(_06433_),
    .A2_N(_06435_),
    .B1(_06433_),
    .B2(_06435_),
    .X(_02572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14439_ (.A(_02572_),
    .Y(_02424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14440_ (.A(\design_top.core0.NXPC[29] ),
    .Y(_02426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14441_ (.A1(_00892_),
    .A2(_06419_),
    .B1(_02405_),
    .Y(_06436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14442_ (.A(_06436_),
    .Y(_06437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14443_ (.A1(_01319_),
    .A2(_06437_),
    .B1(_07865_),
    .B2(_06436_),
    .X(_02427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14444_ (.A(_06837_),
    .X(_00871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14445_ (.A(_01268_),
    .Y(_06438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14446_ (.A1(_00871_),
    .A2(_01268_),
    .B1(_06669_),
    .B2(_06438_),
    .X(_06439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14447_ (.A1_N(_00885_),
    .A2_N(_01269_),
    .B1(_06425_),
    .B2(_06428_),
    .X(_06440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14448_ (.A1_N(_06439_),
    .A2_N(_06440_),
    .B1(_06439_),
    .B2(_06440_),
    .X(_02428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14449_ (.A(_06114_),
    .B(_02083_),
    .X(_02434_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14450_ (.A(_02437_),
    .B(_06393_),
    .C(_06394_),
    .X(_02438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14451_ (.A1_N(_06674_),
    .A2_N(\design_top.core0.PC[28] ),
    .B1(_06433_),
    .B2(_06434_),
    .X(_06441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14452_ (.A(_06668_),
    .B(\design_top.core0.PC[29] ),
    .Y(_06442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _14453_ (.A1(_06668_),
    .A2(\design_top.core0.PC[29] ),
    .B1(_06442_),
    .X(_06443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14454_ (.A1_N(_06441_),
    .A2_N(_06443_),
    .B1(_06441_),
    .B2(_06443_),
    .X(_02576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14455_ (.A(_02576_),
    .Y(_02445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14456_ (.A(\design_top.core0.NXPC[30] ),
    .Y(_02447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14457_ (.A(_06669_),
    .B(_00877_),
    .Y(_00878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14458_ (.A1(_00878_),
    .A2(_06437_),
    .B1(_00879_),
    .X(_06444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14459_ (.A1_N(_01320_),
    .A2_N(_06444_),
    .B1(_01320_),
    .B2(_06444_),
    .X(_02448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14460_ (.A1_N(_06666_),
    .A2_N(_01267_),
    .B1(_06666_),
    .B2(_01267_),
    .X(_06445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14461_ (.A(_06439_),
    .Y(_06446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14462_ (.A1_N(_06426_),
    .A2_N(_01269_),
    .B1(_06669_),
    .B2(_06438_),
    .X(_06447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14463_ (.A1(_06669_),
    .A2(_06438_),
    .B1(_06447_),
    .Y(_06448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _14464_ (.A1(_06427_),
    .A2(_06446_),
    .A3(_06424_),
    .B1(_06448_),
    .X(_06449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14465_ (.A1_N(_06445_),
    .A2_N(_06449_),
    .B1(_06445_),
    .B2(_06449_),
    .X(_02449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14466_ (.A(_06114_),
    .B(_02109_),
    .X(_02455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14467_ (.A(_02458_),
    .B(_06029_),
    .C(_06031_),
    .X(_02459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14468_ (.A(\design_top.core0.PC[30] ),
    .Y(_06450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14469_ (.A1(\design_top.core0.SIMM[30] ),
    .A2(\design_top.core0.PC[30] ),
    .B1(_01338_),
    .B2(_06450_),
    .X(_06451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14470_ (.A1_N(_06668_),
    .A2_N(\design_top.core0.PC[29] ),
    .B1(_06441_),
    .B2(_06442_),
    .X(_06452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14471_ (.A1_N(_06451_),
    .A2_N(_06452_),
    .B1(_06451_),
    .B2(_06452_),
    .X(_02466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14472_ (.A(io_out[18]),
    .Y(_02470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14473_ (.A(io_out[19]),
    .B(io_out[18]),
    .Y(_06453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14474_ (.A1(io_out[19]),
    .A2(io_out[18]),
    .B1(_06453_),
    .X(_02473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14475_ (.A(_06453_),
    .Y(_06454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2bb2a_2 _14476_ (.A1_N(_07803_),
    .A2_N(_06454_),
    .B1(_07803_),
    .B2(_06454_),
    .X(_02476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _14477_ (.A(\design_top.IADDR[4] ),
    .B(_06454_),
    .C(\design_top.IADDR[5] ),
    .X(_06455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _14478_ (.A1(_07803_),
    .A2(_06454_),
    .B1(\design_top.IADDR[5] ),
    .Y(_06456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14479_ (.A(_06455_),
    .B(_06456_),
    .Y(_02479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14480_ (.A(\design_top.IADDR[6] ),
    .B(_06455_),
    .Y(_06457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14481_ (.A1(\design_top.IADDR[6] ),
    .A2(_06455_),
    .B1(_06457_),
    .X(_02483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14482_ (.A(_06457_),
    .Y(_06458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14483_ (.A(\design_top.IADDR[7] ),
    .B(_06458_),
    .Y(_06459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14484_ (.A1(\design_top.IADDR[7] ),
    .A2(_06458_),
    .B1(_06459_),
    .X(_02487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14485_ (.A1(_01336_),
    .A2(_01198_),
    .B1(_06762_),
    .B2(_06855_),
    .X(_06460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _14486_ (.A1_N(_06765_),
    .A2_N(_06460_),
    .B1(_06765_),
    .B2(_06460_),
    .Y(_02489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14487_ (.A(_06459_),
    .Y(_06461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14488_ (.A(\design_top.IADDR[8] ),
    .B(_06461_),
    .Y(_06462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14489_ (.A1(\design_top.IADDR[8] ),
    .A2(_06461_),
    .B1(_06462_),
    .X(_02491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14490_ (.A(_01978_),
    .Y(_02492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14491_ (.A(_06797_),
    .X(_06463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14492_ (.A(_06463_),
    .Y(_06464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14493_ (.A1(_06463_),
    .A2(_06800_),
    .B1(_06464_),
    .B2(_06799_),
    .X(_02493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14494_ (.A(_06462_),
    .Y(_06465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14495_ (.A(\design_top.IADDR[9] ),
    .B(_06465_),
    .Y(_06466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14496_ (.A1(\design_top.IADDR[9] ),
    .A2(_06465_),
    .B1(_06466_),
    .X(_02495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14497_ (.A(_02001_),
    .Y(_02496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14498_ (.A1(_01360_),
    .A2(_01171_),
    .B1(_06463_),
    .B2(_06800_),
    .X(_06467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14499_ (.A(_06467_),
    .Y(_06468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14500_ (.A1(_06802_),
    .A2(_06467_),
    .B1(_06801_),
    .B2(_06468_),
    .X(_02497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14501_ (.A(\design_top.IADDR[10] ),
    .Y(_06469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14502_ (.A(_06469_),
    .B(_06466_),
    .Y(_06470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _14503_ (.A1(_06469_),
    .A2(_06466_),
    .B1(_06470_),
    .Y(_02499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14504_ (.A(_02025_),
    .Y(_02500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _14505_ (.A1(_06800_),
    .A2(_06802_),
    .A3(_06463_),
    .B1(_06753_),
    .X(_06471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14506_ (.A(_06471_),
    .Y(_06472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14507_ (.A1(_06744_),
    .A2(_06471_),
    .B1(_06743_),
    .B2(_06472_),
    .X(_02501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _14508_ (.A(_06466_),
    .B(_06469_),
    .C_N(\design_top.IADDR[11] ),
    .X(_06473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14509_ (.A1(\design_top.IADDR[11] ),
    .A2(_06470_),
    .B1(_06473_),
    .X(_02503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14510_ (.A(_02048_),
    .Y(_02504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14511_ (.A1(_01358_),
    .A2(_01142_),
    .B1(_06744_),
    .B2(_06471_),
    .X(_06474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14512_ (.A(_06474_),
    .Y(_06475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14513_ (.A1(_06747_),
    .A2(_06474_),
    .B1(_06746_),
    .B2(_06475_),
    .X(_02505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14514_ (.A(_06473_),
    .Y(_06476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14515_ (.A(\design_top.IADDR[12] ),
    .B(_06476_),
    .Y(_06477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14516_ (.A1(\design_top.IADDR[12] ),
    .A2(_06476_),
    .B1(_06477_),
    .X(_02507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14517_ (.A(_02072_),
    .Y(_02508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14518_ (.A1(_06463_),
    .A2(_06803_),
    .B1(_06756_),
    .Y(_06478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14519_ (.A(_06478_),
    .Y(_06479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14520_ (.A1(_06728_),
    .A2(_06479_),
    .B1(_06727_),
    .B2(_06478_),
    .X(_02509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14521_ (.A(_06477_),
    .Y(_06480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14522_ (.A(\design_top.IADDR[13] ),
    .B(_06480_),
    .Y(_06481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14523_ (.A1(\design_top.IADDR[13] ),
    .A2(_06480_),
    .B1(_06481_),
    .X(_02511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14524_ (.A(_02095_),
    .Y(_02512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14525_ (.A1(_01356_),
    .A2(_01116_),
    .B1(_06728_),
    .B2(_06479_),
    .X(_06482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14526_ (.A(_06482_),
    .Y(_06483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14527_ (.A1(_06732_),
    .A2(_06482_),
    .B1(_06731_),
    .B2(_06483_),
    .X(_02513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14528_ (.A(_06481_),
    .Y(_06484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14529_ (.A(\design_top.IADDR[14] ),
    .B(_06484_),
    .Y(_06485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14530_ (.A1(\design_top.IADDR[14] ),
    .A2(_06484_),
    .B1(_06485_),
    .X(_02515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14531_ (.A(_02121_),
    .Y(_02516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _14532_ (.A1(_06728_),
    .A2(_06732_),
    .A3(_06479_),
    .B1(_06807_),
    .X(_06486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14533_ (.A(_06486_),
    .Y(_06487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14534_ (.A1(_06736_),
    .A2(_06486_),
    .B1(_06735_),
    .B2(_06487_),
    .X(_02517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14535_ (.A(_06485_),
    .Y(_06488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14536_ (.A(\design_top.IADDR[15] ),
    .B(_06488_),
    .Y(_06489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14537_ (.A1(\design_top.IADDR[15] ),
    .A2(_06488_),
    .B1(_06489_),
    .X(_02519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14538_ (.A(_02143_),
    .Y(_02520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14539_ (.A1(_01354_),
    .A2(_01089_),
    .B1(_06736_),
    .B2(_06486_),
    .X(_06490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14540_ (.A(_06490_),
    .Y(_06491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14541_ (.A1(_06739_),
    .A2(_06490_),
    .B1(_06738_),
    .B2(_06491_),
    .X(_02521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14542_ (.A(_06489_),
    .Y(_06492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14543_ (.A(\design_top.IADDR[16] ),
    .B(_06492_),
    .Y(_06493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14544_ (.A1(\design_top.IADDR[16] ),
    .A2(_06492_),
    .B1(_06493_),
    .X(_02523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14545_ (.A(_02166_),
    .Y(_02524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14546_ (.A(_06813_),
    .Y(_06494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14547_ (.A1(_06813_),
    .A2(_06817_),
    .B1(_06494_),
    .B2(_06816_),
    .X(_02525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14548_ (.A(_06493_),
    .Y(_06495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14549_ (.A(\design_top.IADDR[17] ),
    .B(_06495_),
    .Y(_06496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14550_ (.A1(\design_top.IADDR[17] ),
    .A2(_06495_),
    .B1(_06496_),
    .X(_02527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14551_ (.A(_02187_),
    .Y(_02528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14552_ (.A1(_06717_),
    .A2(_06718_),
    .B1(_06494_),
    .B2(_06816_),
    .X(_06497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14553_ (.A1_N(_06814_),
    .A2_N(_06497_),
    .B1(_06814_),
    .B2(_06497_),
    .X(_02529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14554_ (.A(\design_top.IADDR[18] ),
    .Y(_06498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14555_ (.A(_06498_),
    .B(_06496_),
    .Y(_06499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _14556_ (.A1(_06498_),
    .A2(_06496_),
    .B1(_06499_),
    .Y(_02531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14557_ (.A(_02209_),
    .Y(_02532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _14558_ (.A1(_06814_),
    .A2(_06817_),
    .A3(_06813_),
    .B1(_06720_),
    .X(_06500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14559_ (.A(_06500_),
    .Y(_06501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14560_ (.A1(_06713_),
    .A2(_06500_),
    .B1(_06712_),
    .B2(_06501_),
    .X(_02533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _14561_ (.A(_06496_),
    .B(_06498_),
    .C_N(\design_top.IADDR[19] ),
    .X(_06502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14562_ (.A1(\design_top.IADDR[19] ),
    .A2(_06499_),
    .B1(_06502_),
    .X(_02535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14563_ (.A(_02230_),
    .Y(_02536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14564_ (.A1(_01350_),
    .A2(_01020_),
    .B1(_06713_),
    .B2(_06500_),
    .X(_06503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14565_ (.A(_06503_),
    .Y(_06504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14566_ (.A1(_06709_),
    .A2(_06503_),
    .B1(_06708_),
    .B2(_06504_),
    .X(_02537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14567_ (.A(_06502_),
    .Y(_06505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14568_ (.A(\design_top.IADDR[20] ),
    .B(_06505_),
    .Y(_06506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14569_ (.A1(\design_top.IADDR[20] ),
    .A2(_06505_),
    .B1(_06506_),
    .X(_02539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14570_ (.A(_02252_),
    .Y(_02540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14571_ (.A1(_06813_),
    .A2(_06818_),
    .B1(_06723_),
    .Y(_06507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14572_ (.A(_06507_),
    .Y(_06508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14573_ (.A1(_06693_),
    .A2(_06508_),
    .B1(_06692_),
    .B2(_06507_),
    .X(_02541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14574_ (.A(_06506_),
    .Y(_06509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14575_ (.A(\design_top.IADDR[21] ),
    .B(_06509_),
    .Y(_06510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14576_ (.A1(\design_top.IADDR[21] ),
    .A2(_06509_),
    .B1(_06510_),
    .X(_02543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14577_ (.A(_02273_),
    .Y(_02544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14578_ (.A1(_01348_),
    .A2(_00993_),
    .B1(_06693_),
    .B2(_06508_),
    .X(_06511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14579_ (.A(_06511_),
    .Y(_06512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14580_ (.A1(_06696_),
    .A2(_06511_),
    .B1(_06695_),
    .B2(_06512_),
    .X(_02545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14581_ (.A(_06510_),
    .Y(_06513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14582_ (.A(\design_top.IADDR[22] ),
    .B(_06513_),
    .Y(_06514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14583_ (.A1(\design_top.IADDR[22] ),
    .A2(_06513_),
    .B1(_06514_),
    .X(_02547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14584_ (.A(_02295_),
    .Y(_02548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _14585_ (.A1(_06693_),
    .A2(_06696_),
    .A3(_06508_),
    .B1(_06823_),
    .X(_06515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14586_ (.A(_06515_),
    .Y(_06516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14587_ (.A1(_06701_),
    .A2(_06515_),
    .B1(_06700_),
    .B2(_06516_),
    .X(_02549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14588_ (.A(_06514_),
    .Y(_06517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14589_ (.A(\design_top.IADDR[23] ),
    .B(_06517_),
    .Y(_06518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14590_ (.A1(\design_top.IADDR[23] ),
    .A2(_06517_),
    .B1(_06518_),
    .X(_02551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14591_ (.A(_02316_),
    .Y(_02552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14592_ (.A1(_01346_),
    .A2(_00966_),
    .B1(_06701_),
    .B2(_06515_),
    .X(_06519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14593_ (.A(_06519_),
    .Y(_06520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14594_ (.A1(_06705_),
    .A2(_06519_),
    .B1(_06704_),
    .B2(_06520_),
    .X(_02553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14595_ (.A(_06518_),
    .Y(_06521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14596_ (.A(\design_top.IADDR[24] ),
    .B(_06521_),
    .Y(_06522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14597_ (.A1(\design_top.IADDR[24] ),
    .A2(_06521_),
    .B1(_06522_),
    .X(_02555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14598_ (.A(_02338_),
    .Y(_02556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14599_ (.A(_06826_),
    .Y(_06523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14600_ (.A1(_06826_),
    .A2(_06829_),
    .B1(_06523_),
    .B2(_06828_),
    .X(_02557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14601_ (.A(_06522_),
    .Y(_06524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14602_ (.A(\design_top.IADDR[25] ),
    .B(_06524_),
    .Y(_06525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14603_ (.A1(\design_top.IADDR[25] ),
    .A2(_06524_),
    .B1(_06525_),
    .X(_02559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14604_ (.A(_02359_),
    .Y(_02560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14605_ (.A1(_01344_),
    .A2(_00939_),
    .B1(_06826_),
    .B2(_06829_),
    .X(_06526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14606_ (.A(_06526_),
    .Y(_06527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14607_ (.A1(_06832_),
    .A2(_06526_),
    .B1(_06831_),
    .B2(_06527_),
    .X(_02561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14608_ (.A(\design_top.IADDR[26] ),
    .Y(_06528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14609_ (.A(_06528_),
    .B(_06525_),
    .Y(_06529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _14610_ (.A1(_06528_),
    .A2(_06525_),
    .B1(_06529_),
    .Y(_02563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14611_ (.A(_02381_),
    .Y(_02564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o31a_2 _14612_ (.A1(_06829_),
    .A2(_06832_),
    .A3(_06826_),
    .B1(_06688_),
    .X(_06530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _14613_ (.A1_N(_06679_),
    .A2_N(_06530_),
    .B1(_06679_),
    .B2(_06530_),
    .Y(_02565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3b_2 _14614_ (.A(_06525_),
    .B(_06528_),
    .C_N(\design_top.IADDR[27] ),
    .X(_06531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14615_ (.A1(\design_top.IADDR[27] ),
    .A2(_06529_),
    .B1(_06531_),
    .X(_02567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14616_ (.A(_02402_),
    .Y(_02568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14617_ (.A1(_01342_),
    .A2(_00912_),
    .B1(_06679_),
    .B2(_06530_),
    .X(_06532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _14618_ (.A1_N(_06681_),
    .A2_N(_06532_),
    .B1(_06681_),
    .B2(_06532_),
    .Y(_02569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14619_ (.A(_06531_),
    .Y(_06533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14620_ (.A(\design_top.IADDR[28] ),
    .B(_06533_),
    .Y(_06534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14621_ (.A1(\design_top.IADDR[28] ),
    .A2(_06533_),
    .B1(_06534_),
    .X(_02571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14622_ (.A(_06836_),
    .Y(_06535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14623_ (.A1(_06836_),
    .A2(_06676_),
    .B1(_06535_),
    .B2(_06675_),
    .X(_02573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14624_ (.A(_06534_),
    .Y(_06536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14625_ (.A(\design_top.IADDR[29] ),
    .B(_06536_),
    .Y(_06537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14626_ (.A1(\design_top.IADDR[29] ),
    .A2(_06536_),
    .B1(_06537_),
    .X(_02575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14627_ (.A1(_01340_),
    .A2(_00885_),
    .B1(_06836_),
    .B2(_06676_),
    .X(_06538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14628_ (.A(_06538_),
    .Y(_06539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14629_ (.A1(_06672_),
    .A2(_06538_),
    .B1(_06671_),
    .B2(_06539_),
    .X(_02577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14630_ (.A(_06537_),
    .Y(_06540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14631_ (.A(\design_top.IADDR[30] ),
    .B(_06540_),
    .Y(_06541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14632_ (.A1(\design_top.IADDR[30] ),
    .A2(_06540_),
    .B1(_06541_),
    .X(_02579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14633_ (.A(_02466_),
    .Y(_02580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2oi_2 _14634_ (.A1_N(_06667_),
    .A2_N(_06839_),
    .B1(_06667_),
    .B2(_06839_),
    .Y(_02581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14635_ (.A(\design_top.IADDR[31] ),
    .Y(_06542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a32o_2 _14636_ (.A1(\design_top.IADDR[30] ),
    .A2(_06540_),
    .A3(_06542_),
    .B1(\design_top.IADDR[31] ),
    .B2(_06541_),
    .X(_02583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _14637_ (.A1(_01338_),
    .A2(_06450_),
    .B1(_06451_),
    .B2(_06452_),
    .Y(_06543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14638_ (.A1_N(_00763_),
    .A2_N(\design_top.core0.PC[31] ),
    .B1(_00763_),
    .B2(\design_top.core0.PC[31] ),
    .X(_06544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14639_ (.A1_N(_06543_),
    .A2_N(_06544_),
    .B1(_06543_),
    .B2(_06544_),
    .X(_02584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14640_ (.A(_02584_),
    .Y(_02585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14641_ (.A(_07953_),
    .B(_07926_),
    .X(_02587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14642_ (.A(_05999_),
    .B(_01363_),
    .Y(_01365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14643_ (.A(_05994_),
    .B(_01366_),
    .Y(_01323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14644_ (.A(_07809_),
    .B(_01366_),
    .Y(_01263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14645_ (.A(_07809_),
    .B(_01363_),
    .Y(_01265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _14646_ (.A(_07780_),
    .B(_05980_),
    .C(_05994_),
    .X(_01287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and3_2 _14647_ (.A(_07780_),
    .B(\design_top.core0.FCT3[0] ),
    .C(\design_top.core0.FCT3[2] ),
    .X(_01289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14648_ (.A(_07864_),
    .Y(_01321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14649_ (.A1(_06027_),
    .A2(_06024_),
    .B1(_01521_),
    .Y(_01291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2b_2 _14650_ (.A_N(_07878_),
    .B(_01291_),
    .Y(_01322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14651_ (.A(_06666_),
    .X(_00857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14652_ (.A1(_00925_),
    .A2(_00930_),
    .B1(_00939_),
    .B2(_00944_),
    .X(_06545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _14653_ (.A1(_00857_),
    .A2(_00862_),
    .B1(_00871_),
    .B2(_00876_),
    .Y(_06546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14654_ (.A(_00862_),
    .Y(_06547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22oi_2 _14655_ (.A1(_00871_),
    .A2(_00876_),
    .B1(_06426_),
    .B2(_00890_),
    .Y(_06548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221ai_2 _14656_ (.A1(_00939_),
    .A2(_00944_),
    .B1(_06665_),
    .B2(_06547_),
    .C1(_06548_),
    .Y(_06549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14657_ (.A(_00843_),
    .B(_00848_),
    .Y(_06550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _14658_ (.A1(_06062_),
    .A2(_00848_),
    .B1(_06550_),
    .X(_06551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _14659_ (.A1(_00898_),
    .A2(_00903_),
    .B1(_06426_),
    .B2(_00890_),
    .Y(_06552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14660_ (.A1(_00898_),
    .A2(_00903_),
    .B1(_06401_),
    .B2(_00917_),
    .X(_06553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14661_ (.A1(_06401_),
    .A2(_00917_),
    .B1(_00925_),
    .B2(_00930_),
    .X(_06554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4b_2 _14662_ (.A(_06551_),
    .B(_06552_),
    .C(_06553_),
    .D_N(_06554_),
    .X(_06555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _14663_ (.A(_06545_),
    .B(_06546_),
    .C(_06549_),
    .D(_06555_),
    .X(_06556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14664_ (.A1(_05997_),
    .A2(_00809_),
    .B1(_06001_),
    .B2(_06781_),
    .X(_06557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14665_ (.A1(_01237_),
    .A2(_06848_),
    .B1(_06006_),
    .B2(_06779_),
    .X(_06558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14666_ (.A1(_01215_),
    .A2(_01534_),
    .B1(_01229_),
    .B2(_01224_),
    .X(_06559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14667_ (.A(_01215_),
    .B(_01534_),
    .X(_06560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14668_ (.A1(_01229_),
    .A2(_01224_),
    .B1(_05997_),
    .B2(_00809_),
    .X(_06561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _14669_ (.A1(_06001_),
    .A2(_06781_),
    .B1(_06560_),
    .C1(_06561_),
    .X(_06562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14670_ (.A(_01245_),
    .B(_00793_),
    .X(_06563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14671_ (.A1(_05992_),
    .A2(_06764_),
    .B1(_06011_),
    .B2(_06761_),
    .X(_06564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14672_ (.A1(_01203_),
    .A2(_01198_),
    .B1(_01189_),
    .B2(_01184_),
    .C1(_06564_),
    .X(_06565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2111ai_2 _14673_ (.A1(_06004_),
    .A2(_07826_),
    .B1(_06562_),
    .C1(_06563_),
    .D1(_06565_),
    .Y(_06566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _14674_ (.A(_06557_),
    .B(_06558_),
    .C(_06559_),
    .D(_06566_),
    .X(_06567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14675_ (.A1(_06343_),
    .A2(_00984_),
    .B1(_06323_),
    .B2(_00998_),
    .X(_06568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14676_ (.A1(_01062_),
    .A2(_01067_),
    .B1(_06289_),
    .B2(_01053_),
    .X(_06569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14677_ (.A1(_01062_),
    .A2(_01067_),
    .B1(_06289_),
    .B2(_01053_),
    .X(_06570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221ai_2 _14678_ (.A1(_00979_),
    .A2(_00984_),
    .B1(_00993_),
    .B2(_00998_),
    .C1(_06570_),
    .Y(_06571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14679_ (.A(_01011_),
    .Y(_06572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14680_ (.A(_01006_),
    .B(_01011_),
    .X(_06573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21boi_2 _14681_ (.A1(_06300_),
    .A2(_01025_),
    .B1_N(_06573_),
    .Y(_06574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14682_ (.A1(_07851_),
    .A2(_06572_),
    .B1(_06300_),
    .B2(_01025_),
    .C1(_06574_),
    .X(_06575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14683_ (.A(_00957_),
    .Y(_06576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22oi_2 _14684_ (.A1(_06360_),
    .A2(_06576_),
    .B1(_06698_),
    .B2(_00971_),
    .Y(_06577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14685_ (.A1(_06360_),
    .A2(_06576_),
    .B1(_06352_),
    .B2(_00971_),
    .C1(_06577_),
    .X(_06578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2_2 _14686_ (.A(_06575_),
    .B(_06578_),
    .Y(_06579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4_2 _14687_ (.A(_06568_),
    .B(_06569_),
    .C(_06571_),
    .D(_06579_),
    .X(_06580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14688_ (.A1(_01080_),
    .A2(_01075_),
    .B1(_01094_),
    .B2(_06248_),
    .X(_06581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14689_ (.A1(_06015_),
    .A2(_07840_),
    .B1(_06014_),
    .B2(_06749_),
    .X(_06582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14690_ (.A1(_01107_),
    .A2(_01102_),
    .B1(_01121_),
    .B2(_06224_),
    .X(_06583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14691_ (.A1(_01107_),
    .A2(_01102_),
    .B1(_01094_),
    .B2(_01089_),
    .X(_06584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4b_2 _14692_ (.A(_06581_),
    .B(_06582_),
    .C(_06583_),
    .D_N(_06584_),
    .X(_06585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14693_ (.A1(_06017_),
    .A2(_06754_),
    .B1(_06015_),
    .B2(_07840_),
    .X(_06586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14694_ (.A1(_01176_),
    .A2(_01171_),
    .B1(_01133_),
    .B2(_01540_),
    .X(_06587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14695_ (.A1(_01080_),
    .A2(_01075_),
    .B1(_01121_),
    .B2(_06224_),
    .C1(_06587_),
    .X(_06588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14696_ (.A1(_06013_),
    .A2(_06751_),
    .B1(_06014_),
    .B2(_06749_),
    .X(_06589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and4b_2 _14697_ (.A_N(_06585_),
    .B(_06586_),
    .C(_06588_),
    .D(_06589_),
    .X(_06590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or4b_2 _14698_ (.A(_06556_),
    .B(_06567_),
    .C(_06580_),
    .D_N(_06590_),
    .X(_06591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14699_ (.A(_00848_),
    .Y(_06592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211ai_2 _14700_ (.A1(_00952_),
    .A2(_00957_),
    .B1(_00966_),
    .C1(_00971_),
    .Y(_06593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o211a_2 _14701_ (.A1(_06289_),
    .A2(_01053_),
    .B1(_06569_),
    .C1(_06575_),
    .X(_06594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a32o_2 _14702_ (.A1(_01020_),
    .A2(_01025_),
    .A3(_06573_),
    .B1(_01006_),
    .B2(_01011_),
    .X(_06595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14703_ (.A1(_00993_),
    .A2(_00998_),
    .B1(_06594_),
    .B2(_06595_),
    .X(_06596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221ai_2 _14704_ (.A1(_00979_),
    .A2(_00984_),
    .B1(_06568_),
    .B2(_06596_),
    .C1(_06578_),
    .Y(_06597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14705_ (.A1(_06582_),
    .A2(_06589_),
    .B1(_06586_),
    .Y(_06598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14706_ (.A1(_01133_),
    .A2(_01540_),
    .B1(_01121_),
    .B2(_01116_),
    .C1(_06598_),
    .X(_06599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14707_ (.A1(_06583_),
    .A2(_06599_),
    .B1(_06584_),
    .X(_06600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14708_ (.A1(_01080_),
    .A2(_01075_),
    .B1(_06581_),
    .B2(_06600_),
    .X(_06601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14709_ (.A(_06564_),
    .Y(_06602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221ai_2 _14710_ (.A1(_06001_),
    .A2(_06781_),
    .B1(_06004_),
    .B2(_07826_),
    .C1(_06557_),
    .Y(_06603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a22o_2 _14711_ (.A1(_01237_),
    .A2(_06848_),
    .B1(_06563_),
    .B2(_06603_),
    .X(_06604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14712_ (.A1(_01237_),
    .A2(_06848_),
    .B1(_01229_),
    .B2(_01224_),
    .C1(_06604_),
    .X(_06605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14713_ (.A1(_01203_),
    .A2(_01198_),
    .B1(_06559_),
    .B2(_06605_),
    .C1(_06560_),
    .X(_06606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14714_ (.A1(_01189_),
    .A2(_01184_),
    .B1(_06602_),
    .B2(_06606_),
    .C1(_06590_),
    .X(_06607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21bai_2 _14715_ (.A1(_06601_),
    .A2(_06607_),
    .B1_N(_06580_),
    .Y(_06608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o2111a_2 _14716_ (.A1(_06360_),
    .A2(_06576_),
    .B1(_06593_),
    .C1(_06597_),
    .D1(_06608_),
    .X(_06609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21oi_2 _14717_ (.A1(_06545_),
    .A2(_06554_),
    .B1(_06553_),
    .Y(_06610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14718_ (.A1(_06552_),
    .A2(_06610_),
    .B1(_06548_),
    .X(_06611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22ai_2 _14719_ (.A1(_06665_),
    .A2(_06547_),
    .B1(_06546_),
    .B2(_06611_),
    .Y(_06612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14720_ (.A1(_06062_),
    .A2(_00848_),
    .B1(_06612_),
    .Y(_06613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221ai_2 _14721_ (.A1(_06082_),
    .A2(_06592_),
    .B1(_06556_),
    .B2(_06609_),
    .C1(_06613_),
    .Y(_06614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _14722_ (.A(_06591_),
    .B(_06614_),
    .X(_01288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14723_ (.A(_01266_),
    .Y(_06615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14724_ (.A(_06082_),
    .B(_06615_),
    .Y(_06616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _14725_ (.A1(_06082_),
    .A2(_06615_),
    .B1(_06616_),
    .X(_06617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14726_ (.A(_06445_),
    .B(_06617_),
    .X(_06618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14727_ (.A(_06427_),
    .B(_06446_),
    .C(_06618_),
    .X(_06619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _14728_ (.A1(_00857_),
    .A2(_01267_),
    .A3(_06616_),
    .B1(_06062_),
    .B2(_01266_),
    .X(_06620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221ai_2 _14729_ (.A1(_06448_),
    .A2(_06618_),
    .B1(_06424_),
    .B2(_06619_),
    .C1(_06620_),
    .Y(_01286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14730_ (.A1(_06082_),
    .A2(_06592_),
    .B1(_06550_),
    .B2(_06614_),
    .C1(_06591_),
    .X(_01264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14731_ (.A(\design_top.TIMER[0] ),
    .Y(_02912_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14732_ (.A1(\design_top.TIMER[1] ),
    .A2(\design_top.TIMER[0] ),
    .B1_N(_07005_),
    .X(_02913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14733_ (.A1(\design_top.TIMER[2] ),
    .A2(_07005_),
    .B1_N(_07006_),
    .X(_02914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14734_ (.A1(\design_top.TIMER[3] ),
    .A2(_07006_),
    .B1_N(_07007_),
    .X(_02915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14735_ (.A1(\design_top.TIMER[4] ),
    .A2(_07007_),
    .B1_N(_07008_),
    .X(_02916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14736_ (.A1(\design_top.TIMER[5] ),
    .A2(_07008_),
    .B1_N(_07009_),
    .X(_02917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14737_ (.A1(\design_top.TIMER[6] ),
    .A2(_07009_),
    .B1_N(_07010_),
    .X(_02918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14738_ (.A1(\design_top.TIMER[7] ),
    .A2(_07010_),
    .B1_N(_07011_),
    .X(_02919_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14739_ (.A1(\design_top.TIMER[8] ),
    .A2(_07011_),
    .B1_N(_07012_),
    .X(_02920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14740_ (.A1(\design_top.TIMER[9] ),
    .A2(_07012_),
    .B1_N(_07013_),
    .X(_02921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14741_ (.A1(\design_top.TIMER[10] ),
    .A2(_07013_),
    .B1_N(_07014_),
    .X(_02922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14742_ (.A1(\design_top.TIMER[11] ),
    .A2(_07014_),
    .B1_N(_07015_),
    .X(_02923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14743_ (.A1(\design_top.TIMER[12] ),
    .A2(_07015_),
    .B1_N(_07016_),
    .X(_02924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14744_ (.A1(\design_top.TIMER[13] ),
    .A2(_07016_),
    .B1_N(_07017_),
    .X(_02925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14745_ (.A1(\design_top.TIMER[14] ),
    .A2(_07017_),
    .B1_N(_07018_),
    .X(_02926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14746_ (.A1(\design_top.TIMER[15] ),
    .A2(_07018_),
    .B1_N(_07019_),
    .X(_02927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14747_ (.A(\design_top.TIMER[16] ),
    .B(_07019_),
    .X(_06621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14748_ (.A1(\design_top.TIMER[16] ),
    .A2(_07019_),
    .B1_N(_06621_),
    .X(_02928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14749_ (.A1(\design_top.TIMER[17] ),
    .A2(_06621_),
    .B1_N(_07020_),
    .X(_02929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14750_ (.A(\design_top.TIMER[18] ),
    .B(_07020_),
    .X(_06622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14751_ (.A1(\design_top.TIMER[18] ),
    .A2(_07020_),
    .B1_N(_06622_),
    .X(_02930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14752_ (.A1(\design_top.TIMER[19] ),
    .A2(_06622_),
    .B1_N(_07021_),
    .X(_02931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14753_ (.A(\design_top.TIMER[20] ),
    .B(_07021_),
    .X(_06623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14754_ (.A1(\design_top.TIMER[20] ),
    .A2(_07021_),
    .B1_N(_06623_),
    .X(_02932_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14755_ (.A1(\design_top.TIMER[21] ),
    .A2(_06623_),
    .B1_N(_07022_),
    .X(_02933_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14756_ (.A(\design_top.TIMER[22] ),
    .B(_07022_),
    .X(_06624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14757_ (.A1(\design_top.TIMER[22] ),
    .A2(_07022_),
    .B1_N(_06624_),
    .X(_02934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14758_ (.A1(\design_top.TIMER[23] ),
    .A2(_06624_),
    .B1_N(_07023_),
    .X(_02935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14759_ (.A(\design_top.TIMER[24] ),
    .B(_07023_),
    .Y(_06625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21o_2 _14760_ (.A1(\design_top.TIMER[24] ),
    .A2(_07023_),
    .B1(_06625_),
    .X(_02936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14761_ (.A(\design_top.TIMER[25] ),
    .Y(_06626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21ai_2 _14762_ (.A1(_06626_),
    .A2(_06625_),
    .B1(_07024_),
    .Y(_02937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14763_ (.A1(\design_top.TIMER[26] ),
    .A2(_07024_),
    .B1_N(_07025_),
    .X(_02938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14764_ (.A1(\design_top.TIMER[27] ),
    .A2(_07025_),
    .B1_N(_07026_),
    .X(_02939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14765_ (.A(\design_top.TIMER[28] ),
    .B(_07026_),
    .X(_06627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14766_ (.A1(\design_top.TIMER[28] ),
    .A2(_07026_),
    .B1_N(_06627_),
    .X(_02940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14767_ (.A(\design_top.TIMER[29] ),
    .B(_06627_),
    .X(_06628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a21bo_2 _14768_ (.A1(\design_top.TIMER[29] ),
    .A2(_06627_),
    .B1_N(_06628_),
    .X(_02941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14769_ (.A1_N(\design_top.TIMER[30] ),
    .A2_N(_06628_),
    .B1(\design_top.TIMER[30] ),
    .B2(_06628_),
    .X(_02942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14770_ (.A1(\design_top.TIMER[30] ),
    .A2(_06628_),
    .B1(\design_top.TIMER[31] ),
    .X(_06629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14771_ (.A(_01375_),
    .B(_06629_),
    .X(_02943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14772_ (.A1(_01116_),
    .A2(_01122_),
    .B1(_07830_),
    .B2(_06223_),
    .X(_06630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14773_ (.A1(_01102_),
    .A2(_01108_),
    .B1(_07831_),
    .B2(_06630_),
    .X(_06631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14774_ (.A1(_01089_),
    .A2(_01095_),
    .B1(_07835_),
    .B2(_06631_),
    .X(_06632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14775_ (.A1(_01075_),
    .A2(_01081_),
    .B1(_07833_),
    .B2(_06632_),
    .X(_06633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _14776_ (.A1(_01068_),
    .A2(_01062_),
    .A3(_07855_),
    .B1(_06289_),
    .B2(_01054_),
    .X(_06634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14777_ (.A1(_01020_),
    .A2(_01026_),
    .B1(_07850_),
    .B2(_06634_),
    .X(_06635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14778_ (.A1(_01006_),
    .A2(_01012_),
    .B1(_07853_),
    .B2(_06635_),
    .X(_06636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _14779_ (.A1(_06323_),
    .A2(_00999_),
    .A3(_07871_),
    .B1(_06343_),
    .B2(_00985_),
    .X(_06637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14780_ (.A1(_00966_),
    .A2(_00972_),
    .B1(_07875_),
    .B2(_06637_),
    .X(_06638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14781_ (.A(_07870_),
    .B(_06638_),
    .X(_06639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14782_ (.A1(_00952_),
    .A2(_00958_),
    .B1(_07876_),
    .B2(_06636_),
    .C1(_06639_),
    .X(_06640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _14783_ (.A1(_00945_),
    .A2(_06331_),
    .A3(_07861_),
    .B1(_06390_),
    .B2(_00931_),
    .X(_06641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14784_ (.A1(_00912_),
    .A2(_00918_),
    .B1(_07860_),
    .B2(_06641_),
    .X(_06642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14785_ (.A(_07858_),
    .B(_06642_),
    .X(_06643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14786_ (.A1(_00898_),
    .A2(_00904_),
    .B1(_07863_),
    .B2(_06640_),
    .C1(_06643_),
    .X(_06644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o32a_2 _14787_ (.A1(_06426_),
    .A2(_00891_),
    .A3(_07865_),
    .B1(_00871_),
    .B2(_00877_),
    .X(_06645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14788_ (.A1(_00857_),
    .A2(_00863_),
    .B1(_07867_),
    .B2(_06645_),
    .X(_06646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o221a_2 _14789_ (.A1(_07877_),
    .A2(_06633_),
    .B1(_07868_),
    .B2(_06644_),
    .C1(_06646_),
    .X(_06647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14790_ (.A1_N(_07864_),
    .A2_N(_06647_),
    .B1(_06062_),
    .B2(_00849_),
    .X(_01262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14791_ (.A(_06665_),
    .B(_00863_),
    .Y(_00864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14792_ (.A(_06038_),
    .B(_06769_),
    .Y(_01231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14793_ (.A(_06691_),
    .B(_00999_),
    .Y(_01000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14794_ (.A(\design_top.core0.REG1[12][17] ),
    .Y(_01043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14795_ (.A(\design_top.core0.REG1[13][17] ),
    .Y(_01044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14796_ (.A(_06751_),
    .B(_01177_),
    .Y(_01178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14797_ (.A(\design_top.core0.REG1[10][17] ),
    .Y(_01040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14798_ (.A(\design_top.core0.REG1[11][17] ),
    .Y(_01041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14799_ (.A(\design_top.core0.REG1[14][17] ),
    .Y(_01045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14800_ (.A(\design_top.core0.REG1[15][17] ),
    .Y(_01046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14801_ (.A(\design_top.core0.REG1[4][17] ),
    .Y(_01033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14802_ (.A(\design_top.core0.REG1[5][17] ),
    .Y(_01034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14803_ (.A(\design_top.core0.REG1[6][17] ),
    .Y(_01035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14804_ (.A(\design_top.core0.REG1[7][17] ),
    .Y(_01036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14805_ (.A(\design_top.core0.REG1[8][17] ),
    .Y(_01038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14806_ (.A(\design_top.core0.REG1[9][17] ),
    .Y(_01039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14807_ (.A(\design_top.core0.REG1[1][17] ),
    .Y(_01029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14808_ (.A(\design_top.core0.REG1[2][17] ),
    .Y(_01030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14809_ (.A(\design_top.core0.REG1[3][17] ),
    .Y(_01031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14810_ (.A(_06726_),
    .B(_01122_),
    .Y(_01123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14811_ (.A(\design_top.IDATA[20] ),
    .Y(_06648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14812_ (.A(_07651_),
    .X(_06649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor4_2 _14813_ (.A(_06648_),
    .B(_00009_),
    .C(_00008_),
    .D(_06649_),
    .Y(_00708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14814_ (.A(_07651_),
    .X(_06650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14815_ (.A(_07691_),
    .B(_06650_),
    .Y(_00709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14816_ (.A(_07686_),
    .B(_06650_),
    .Y(_00712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14817_ (.A(_07683_),
    .B(_06650_),
    .Y(_00715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14818_ (.A(_07681_),
    .B(_06650_),
    .Y(_00719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14819_ (.A(_07679_),
    .B(_06650_),
    .Y(_00722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14820_ (.A(_07651_),
    .X(_06651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14821_ (.A(_07677_),
    .B(_06651_),
    .Y(_00725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14822_ (.A(_07672_),
    .B(_06651_),
    .Y(_00728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14823_ (.A(_07670_),
    .B(_06651_),
    .Y(_00731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14824_ (.A(_07666_),
    .B(_06651_),
    .Y(_00734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14825_ (.A(_07661_),
    .B(_06651_),
    .Y(_00737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_1 _14826_ (.A(_07651_),
    .X(_06652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14827_ (.A(_07640_),
    .B(_06652_),
    .Y(_00740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _14828_ (.A(\design_top.IDATA[12] ),
    .B(_06652_),
    .X(_00743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _14829_ (.A(\design_top.IDATA[13] ),
    .B(_06652_),
    .X(_00746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _14830_ (.A(\design_top.IDATA[14] ),
    .B(_06652_),
    .X(_00748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _14831_ (.A(\design_top.IDATA[15] ),
    .B(_06652_),
    .X(_00750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _14832_ (.A(\design_top.IDATA[16] ),
    .B(_06649_),
    .X(_00752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _14833_ (.A(\design_top.IDATA[17] ),
    .B(_06649_),
    .X(_00754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _14834_ (.A(\design_top.IDATA[18] ),
    .B(_06649_),
    .X(_00756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__and2_2 _14835_ (.A(_00665_),
    .B(_06649_),
    .X(_00758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nor2_2 _14836_ (.A(_06648_),
    .B(_00643_),
    .Y(_00760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 _14837_ (.A(\design_top.core0.NXPC[31] ),
    .Y(_00762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o21a_2 _14838_ (.A1(_01320_),
    .A2(_06444_),
    .B1(_00865_),
    .X(_06653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14839_ (.A1_N(_01321_),
    .A2_N(_06653_),
    .B1(_01321_),
    .B2(_06653_),
    .X(_00764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__o22a_2 _14840_ (.A1(_00857_),
    .A2(_01267_),
    .B1(_06445_),
    .B2(_06449_),
    .X(_06654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14841_ (.A1_N(_06617_),
    .A2_N(_06654_),
    .B1(_06617_),
    .B2(_06654_),
    .X(_00765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or2_2 _14842_ (.A(_06114_),
    .B(_02132_),
    .X(_00771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__or3_2 _14843_ (.A(_00773_),
    .B(_06029_),
    .C(_06031_),
    .X(_00774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__nand2b_2 _14844_ (.A_N(\design_top.uart0.UART_RXDFF[1] ),
    .B(_05919_),
    .Y(_00784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__a2bb2o_2 _14845_ (.A1_N(_06892_),
    .A2_N(_06859_),
    .B1(\design_top.MEM[9][31] ),
    .B2(_06871_),
    .X(_05494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14846_ (.LO(io_oeb[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14847_ (.LO(io_oeb[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14848_ (.LO(io_oeb[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14849_ (.LO(io_oeb[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14850_ (.LO(io_oeb[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14851_ (.LO(io_oeb[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14852_ (.LO(io_oeb[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14853_ (.LO(io_oeb[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14854_ (.LO(io_oeb[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14855_ (.LO(io_oeb[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14856_ (.LO(io_oeb[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14857_ (.LO(io_oeb[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14858_ (.LO(io_oeb[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14859_ (.LO(io_oeb[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14860_ (.LO(io_oeb[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14861_ (.LO(io_oeb[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14862_ (.LO(io_oeb[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14863_ (.LO(io_oeb[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14864_ (.LO(io_oeb[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14865_ (.LO(io_oeb[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14866_ (.LO(io_oeb[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14867_ (.LO(io_oeb[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14868_ (.LO(io_oeb[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14869_ (.LO(io_oeb[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14870_ (.LO(io_oeb[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14871_ (.LO(io_oeb[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14872_ (.LO(io_oeb[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14873_ (.LO(io_oeb[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14874_ (.LO(io_oeb[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14875_ (.LO(io_oeb[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14876_ (.LO(io_oeb[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14877_ (.LO(io_oeb[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14878_ (.LO(io_oeb[32]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14879_ (.LO(io_oeb[33]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14880_ (.LO(io_oeb[34]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14881_ (.LO(io_oeb[35]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14882_ (.LO(io_oeb[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14883_ (.LO(io_oeb[37]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14884_ (.LO(io_out[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14885_ (.LO(io_out[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14886_ (.LO(io_out[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14887_ (.LO(io_out[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14888_ (.LO(io_out[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14889_ (.LO(io_out[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14890_ (.LO(io_out[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14891_ (.LO(io_out[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14892_ (.LO(io_out[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14893_ (.LO(io_out[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14894_ (.LO(io_out[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14895_ (.LO(io_out[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14896_ (.LO(io_out[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14897_ (.LO(io_out[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14898_ (.LO(io_out[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14899_ (.LO(io_out[32]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14900_ (.LO(io_out[33]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14901_ (.LO(io_out[34]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14902_ (.LO(io_out[35]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14903_ (.LO(io_out[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14904_ (.LO(io_out[37]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14905_ (.LO(la_data_out[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14906_ (.LO(la_data_out[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14907_ (.LO(la_data_out[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14908_ (.LO(la_data_out[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14909_ (.LO(la_data_out[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14910_ (.LO(la_data_out[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14911_ (.LO(la_data_out[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14912_ (.LO(la_data_out[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14913_ (.LO(la_data_out[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14914_ (.LO(la_data_out[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14915_ (.LO(la_data_out[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14916_ (.LO(la_data_out[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14917_ (.LO(la_data_out[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14918_ (.LO(la_data_out[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14919_ (.LO(la_data_out[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14920_ (.LO(la_data_out[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14921_ (.LO(la_data_out[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14922_ (.LO(la_data_out[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14923_ (.LO(la_data_out[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14924_ (.LO(la_data_out[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14925_ (.LO(la_data_out[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14926_ (.LO(la_data_out[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14927_ (.LO(la_data_out[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14928_ (.LO(la_data_out[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14929_ (.LO(la_data_out[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14930_ (.LO(la_data_out[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14931_ (.LO(la_data_out[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14932_ (.LO(la_data_out[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14933_ (.LO(la_data_out[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14934_ (.LO(la_data_out[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14935_ (.LO(la_data_out[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14936_ (.LO(la_data_out[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14937_ (.LO(la_data_out[32]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14938_ (.LO(la_data_out[33]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14939_ (.LO(la_data_out[34]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14940_ (.LO(la_data_out[35]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14941_ (.LO(la_data_out[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14942_ (.LO(la_data_out[37]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14943_ (.LO(la_data_out[38]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14944_ (.LO(la_data_out[39]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14945_ (.LO(la_data_out[40]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14946_ (.LO(la_data_out[41]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14947_ (.LO(la_data_out[42]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14948_ (.LO(la_data_out[43]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14949_ (.LO(la_data_out[44]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14950_ (.LO(la_data_out[45]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14951_ (.LO(la_data_out[46]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14952_ (.LO(la_data_out[47]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14953_ (.LO(la_data_out[48]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14954_ (.LO(la_data_out[49]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14955_ (.LO(la_data_out[50]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14956_ (.LO(la_data_out[51]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14957_ (.LO(la_data_out[52]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14958_ (.LO(la_data_out[53]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14959_ (.LO(la_data_out[54]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14960_ (.LO(la_data_out[55]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14961_ (.LO(la_data_out[56]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14962_ (.LO(la_data_out[57]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14963_ (.LO(la_data_out[58]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14964_ (.LO(la_data_out[59]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14965_ (.LO(la_data_out[60]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14966_ (.LO(la_data_out[61]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14967_ (.LO(la_data_out[62]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14968_ (.LO(la_data_out[63]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14969_ (.LO(la_data_out[64]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14970_ (.LO(la_data_out[65]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14971_ (.LO(la_data_out[66]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14972_ (.LO(la_data_out[67]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14973_ (.LO(la_data_out[68]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14974_ (.LO(la_data_out[69]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14975_ (.LO(la_data_out[70]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14976_ (.LO(la_data_out[71]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14977_ (.LO(la_data_out[72]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14978_ (.LO(la_data_out[73]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14979_ (.LO(la_data_out[74]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14980_ (.LO(la_data_out[75]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14981_ (.LO(la_data_out[76]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14982_ (.LO(la_data_out[77]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14983_ (.LO(la_data_out[78]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14984_ (.LO(la_data_out[79]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14985_ (.LO(la_data_out[80]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14986_ (.LO(la_data_out[81]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14987_ (.LO(la_data_out[82]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14988_ (.LO(la_data_out[83]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14989_ (.LO(la_data_out[84]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14990_ (.LO(la_data_out[85]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14991_ (.LO(la_data_out[86]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14992_ (.LO(la_data_out[87]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14993_ (.LO(la_data_out[88]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14994_ (.LO(la_data_out[89]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14995_ (.LO(la_data_out[90]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14996_ (.LO(la_data_out[91]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14997_ (.LO(la_data_out[92]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14998_ (.LO(la_data_out[93]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _14999_ (.LO(la_data_out[94]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15000_ (.LO(la_data_out[95]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15001_ (.LO(la_data_out[96]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15002_ (.LO(la_data_out[97]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15003_ (.LO(la_data_out[98]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15004_ (.LO(la_data_out[99]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15005_ (.LO(la_data_out[100]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15006_ (.LO(la_data_out[101]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15007_ (.LO(la_data_out[102]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15008_ (.LO(la_data_out[103]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15009_ (.LO(la_data_out[104]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15010_ (.LO(la_data_out[105]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15011_ (.LO(la_data_out[106]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15012_ (.LO(la_data_out[107]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15013_ (.LO(la_data_out[108]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15014_ (.LO(la_data_out[109]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15015_ (.LO(la_data_out[110]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15016_ (.LO(la_data_out[111]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15017_ (.LO(la_data_out[112]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15018_ (.LO(la_data_out[113]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15019_ (.LO(la_data_out[114]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15020_ (.LO(la_data_out[115]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15021_ (.LO(la_data_out[116]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15022_ (.LO(la_data_out[117]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15023_ (.LO(la_data_out[118]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15024_ (.LO(la_data_out[119]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15025_ (.LO(la_data_out[120]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15026_ (.LO(la_data_out[121]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15027_ (.LO(la_data_out[122]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15028_ (.LO(la_data_out[123]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15029_ (.LO(la_data_out[124]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15030_ (.LO(la_data_out[125]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15031_ (.LO(la_data_out[126]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15032_ (.LO(la_data_out[127]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15033_ (.LO(user_irq[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15034_ (.LO(user_irq[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15035_ (.LO(user_irq[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15036_ (.LO(wbs_ack_o),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15037_ (.LO(wbs_dat_o[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15038_ (.LO(wbs_dat_o[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15039_ (.LO(wbs_dat_o[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15040_ (.LO(wbs_dat_o[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15041_ (.LO(wbs_dat_o[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15042_ (.LO(wbs_dat_o[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15043_ (.LO(wbs_dat_o[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15044_ (.LO(wbs_dat_o[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15045_ (.LO(wbs_dat_o[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15046_ (.LO(wbs_dat_o[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15047_ (.LO(wbs_dat_o[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15048_ (.LO(wbs_dat_o[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15049_ (.LO(wbs_dat_o[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15050_ (.LO(wbs_dat_o[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15051_ (.LO(wbs_dat_o[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15052_ (.LO(wbs_dat_o[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15053_ (.LO(wbs_dat_o[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15054_ (.LO(wbs_dat_o[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15055_ (.LO(wbs_dat_o[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15056_ (.LO(wbs_dat_o[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15057_ (.LO(wbs_dat_o[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15058_ (.LO(wbs_dat_o[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15059_ (.LO(wbs_dat_o[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15060_ (.LO(wbs_dat_o[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15061_ (.LO(wbs_dat_o[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15062_ (.LO(wbs_dat_o[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15063_ (.LO(wbs_dat_o[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15064_ (.LO(wbs_dat_o[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15065_ (.LO(wbs_dat_o[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15066_ (.LO(wbs_dat_o[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15067_ (.LO(wbs_dat_o[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__conb_1 _15068_ (.LO(wbs_dat_o[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _15069_ (.A(io_out[15]),
    .X(\design_top.GPIOFF[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _15070_ (.A(io_out[8]),
    .X(\design_top.LEDFF[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _15071_ (.A(io_out[9]),
    .X(\design_top.LEDFF[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _15072_ (.A(io_out[10]),
    .X(\design_top.LEDFF[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _15073_ (.A(io_out[11]),
    .X(\design_top.LEDFF[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__buf_2 _15074_ (.A(io_out[14]),
    .X(\design_top.XTIMER ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15075_ (.A0(_01289_),
    .A1(_01366_),
    .S(io_out[12]),
    .X(_08561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15076_ (.A0(_01362_),
    .A1(_01525_),
    .S(_01323_),
    .X(_08562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15077_ (.A0(\design_top.ROMFF[0] ),
    .A1(\design_top.ROMFF2[0] ),
    .S(\design_top.HLT2 ),
    .X(io_out[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15078_ (.A0(\design_top.ROMFF[1] ),
    .A1(\design_top.ROMFF2[1] ),
    .S(\design_top.HLT2 ),
    .X(io_out[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15079_ (.A0(\design_top.ROMFF[2] ),
    .A1(\design_top.ROMFF2[2] ),
    .S(\design_top.HLT2 ),
    .X(io_out[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15080_ (.A0(\design_top.ROMFF[3] ),
    .A1(\design_top.ROMFF2[3] ),
    .S(\design_top.HLT2 ),
    .X(io_out[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15081_ (.A0(_01260_),
    .A1(_01425_),
    .S(_01362_),
    .X(_01426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15082_ (.A0(_01426_),
    .A1(_01424_),
    .S(_01323_),
    .X(\design_top.DATAO[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15083_ (.A0(_01253_),
    .A1(_01428_),
    .S(_01362_),
    .X(_01429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15084_ (.A0(_01429_),
    .A1(_01427_),
    .S(_01323_),
    .X(\design_top.DATAO[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15085_ (.A0(_01245_),
    .A1(_01431_),
    .S(_01362_),
    .X(_01432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15086_ (.A0(_01432_),
    .A1(_01430_),
    .S(_01323_),
    .X(\design_top.DATAO[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15087_ (.A0(_01237_),
    .A1(_01434_),
    .S(_01362_),
    .X(_01435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15088_ (.A0(_01435_),
    .A1(_01433_),
    .S(_01323_),
    .X(\design_top.DATAO[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15089_ (.A0(_01229_),
    .A1(_01437_),
    .S(_01362_),
    .X(_01438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15090_ (.A0(_01438_),
    .A1(_01436_),
    .S(_01323_),
    .X(\design_top.DATAO[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15091_ (.A0(_01215_),
    .A1(_01440_),
    .S(_01362_),
    .X(_01441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15092_ (.A0(_01441_),
    .A1(_01439_),
    .S(_01323_),
    .X(\design_top.DATAO[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15093_ (.A0(_01203_),
    .A1(_01443_),
    .S(_01362_),
    .X(_01444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15094_ (.A0(_01444_),
    .A1(_01442_),
    .S(_01323_),
    .X(\design_top.DATAO[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15095_ (.A0(_01189_),
    .A1(_01446_),
    .S(_01362_),
    .X(_01447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15096_ (.A0(_01447_),
    .A1(_01445_),
    .S(_01323_),
    .X(\design_top.DATAO[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15097_ (.A0(_01176_),
    .A1(_01449_),
    .S(_01362_),
    .X(_01450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15098_ (.A0(_01450_),
    .A1(_01448_),
    .S(_01323_),
    .X(\design_top.DATAO[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15099_ (.A0(_01161_),
    .A1(_01452_),
    .S(_01362_),
    .X(_01453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15100_ (.A0(_01453_),
    .A1(_01451_),
    .S(_01323_),
    .X(\design_top.DATAO[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15101_ (.A0(_01147_),
    .A1(_01455_),
    .S(_01362_),
    .X(_01456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15102_ (.A0(_01456_),
    .A1(_01454_),
    .S(_01323_),
    .X(\design_top.DATAO[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15103_ (.A0(_01133_),
    .A1(_01458_),
    .S(_01362_),
    .X(_01459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15104_ (.A0(_01459_),
    .A1(_01457_),
    .S(_01323_),
    .X(\design_top.DATAO[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15105_ (.A0(_01121_),
    .A1(_01461_),
    .S(_01362_),
    .X(_01462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15106_ (.A0(_01462_),
    .A1(_01460_),
    .S(_01323_),
    .X(\design_top.DATAO[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15107_ (.A0(_01107_),
    .A1(_01464_),
    .S(_01362_),
    .X(_01465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15108_ (.A0(_01465_),
    .A1(_01463_),
    .S(_01323_),
    .X(\design_top.DATAO[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15109_ (.A0(_01094_),
    .A1(_01467_),
    .S(_01362_),
    .X(_01468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15110_ (.A0(_01468_),
    .A1(_01466_),
    .S(_01323_),
    .X(\design_top.DATAO[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15111_ (.A0(_01080_),
    .A1(_01470_),
    .S(_01362_),
    .X(_01471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15112_ (.A0(_01471_),
    .A1(_01469_),
    .S(_01323_),
    .X(\design_top.DATAO[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15113_ (.A0(_01067_),
    .A1(_01473_),
    .S(_01362_),
    .X(_01474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15114_ (.A0(_01474_),
    .A1(_01472_),
    .S(_01323_),
    .X(\design_top.DATAO[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15115_ (.A0(_01053_),
    .A1(_01476_),
    .S(_01362_),
    .X(_01477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15116_ (.A0(_01477_),
    .A1(_01475_),
    .S(_01323_),
    .X(\design_top.DATAO[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15117_ (.A0(_01025_),
    .A1(_01479_),
    .S(_01362_),
    .X(_01480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15118_ (.A0(_01480_),
    .A1(_01478_),
    .S(_01323_),
    .X(\design_top.DATAO[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15119_ (.A0(_01011_),
    .A1(_01482_),
    .S(_01362_),
    .X(_01483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15120_ (.A0(_01483_),
    .A1(_01481_),
    .S(_01323_),
    .X(\design_top.DATAO[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15121_ (.A0(_00998_),
    .A1(_01485_),
    .S(_01362_),
    .X(_01486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15122_ (.A0(_01486_),
    .A1(_01484_),
    .S(_01323_),
    .X(\design_top.DATAO[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15123_ (.A0(_00984_),
    .A1(_01488_),
    .S(_01362_),
    .X(_01489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15124_ (.A0(_01489_),
    .A1(_01487_),
    .S(_01323_),
    .X(\design_top.DATAO[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15125_ (.A0(_00971_),
    .A1(_01491_),
    .S(_01362_),
    .X(_01492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15126_ (.A0(_01492_),
    .A1(_01490_),
    .S(_01323_),
    .X(\design_top.DATAO[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15127_ (.A0(_00957_),
    .A1(_01494_),
    .S(_01362_),
    .X(_01495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15128_ (.A0(_01495_),
    .A1(_01493_),
    .S(_01323_),
    .X(\design_top.DATAO[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15129_ (.A0(_00944_),
    .A1(_01497_),
    .S(_01362_),
    .X(_01498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15130_ (.A0(_01498_),
    .A1(_01496_),
    .S(_01323_),
    .X(\design_top.DATAO[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15131_ (.A0(_00930_),
    .A1(_01500_),
    .S(_01362_),
    .X(_01501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15132_ (.A0(_01501_),
    .A1(_01499_),
    .S(_01323_),
    .X(\design_top.DATAO[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15133_ (.A0(_00917_),
    .A1(_01503_),
    .S(_01362_),
    .X(_01504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15134_ (.A0(_01504_),
    .A1(_01502_),
    .S(_01323_),
    .X(\design_top.DATAO[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15135_ (.A0(_00903_),
    .A1(_01506_),
    .S(_01362_),
    .X(_01507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15136_ (.A0(_01507_),
    .A1(_01505_),
    .S(_01323_),
    .X(\design_top.DATAO[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15137_ (.A0(_00890_),
    .A1(_01509_),
    .S(_01362_),
    .X(_01510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15138_ (.A0(_01510_),
    .A1(_01508_),
    .S(_01323_),
    .X(\design_top.DATAO[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15139_ (.A0(_00876_),
    .A1(_01512_),
    .S(_01362_),
    .X(_01513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15140_ (.A0(_01513_),
    .A1(_01511_),
    .S(_01323_),
    .X(\design_top.DATAO[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15141_ (.A0(_00862_),
    .A1(_01515_),
    .S(_01362_),
    .X(_01516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15142_ (.A0(_01516_),
    .A1(_01514_),
    .S(_01323_),
    .X(\design_top.DATAO[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15143_ (.A0(_00848_),
    .A1(_01413_),
    .S(_01362_),
    .X(_01414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15144_ (.A0(_01414_),
    .A1(_01412_),
    .S(_01323_),
    .X(\design_top.DATAO[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15145_ (.A0(\design_top.ROMFF[7] ),
    .A1(\design_top.ROMFF2[7] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15146_ (.A0(\design_top.ROMFF[8] ),
    .A1(\design_top.ROMFF2[8] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15147_ (.A0(\design_top.ROMFF[9] ),
    .A1(\design_top.ROMFF2[9] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15148_ (.A0(\design_top.ROMFF[10] ),
    .A1(\design_top.ROMFF2[10] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15149_ (.A0(\design_top.ROMFF[12] ),
    .A1(\design_top.ROMFF2[12] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15150_ (.A0(\design_top.ROMFF[13] ),
    .A1(\design_top.ROMFF2[13] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15151_ (.A0(\design_top.ROMFF[14] ),
    .A1(\design_top.ROMFF2[14] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15152_ (.A0(\design_top.ROMFF[15] ),
    .A1(\design_top.ROMFF2[15] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15153_ (.A0(\design_top.ROMFF[16] ),
    .A1(\design_top.ROMFF2[16] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15154_ (.A0(\design_top.ROMFF[17] ),
    .A1(\design_top.ROMFF2[17] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15155_ (.A0(\design_top.ROMFF[18] ),
    .A1(\design_top.ROMFF2[18] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15156_ (.A0(\design_top.ROMFF[20] ),
    .A1(\design_top.ROMFF2[20] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15157_ (.A0(\design_top.ROMFF[21] ),
    .A1(\design_top.ROMFF2[21] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15158_ (.A0(\design_top.ROMFF[22] ),
    .A1(\design_top.ROMFF2[22] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15159_ (.A0(\design_top.ROMFF[23] ),
    .A1(\design_top.ROMFF2[23] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15160_ (.A0(\design_top.ROMFF[30] ),
    .A1(\design_top.ROMFF2[30] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15161_ (.A0(\design_top.ROMFF[31] ),
    .A1(\design_top.ROMFF2[31] ),
    .S(\design_top.HLT2 ),
    .X(\design_top.IDATA[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15162_ (.A0(_02588_),
    .A1(_02589_),
    .S(\design_top.uart0.UART_XSTATE[2] ),
    .X(_02590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15163_ (.A0(_02587_),
    .A1(_02590_),
    .S(\design_top.uart0.UART_XSTATE[3] ),
    .X(io_out[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15164_ (.A0(_02591_),
    .A1(_00784_),
    .S(_01370_),
    .X(_00785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15165_ (.A0(_00782_),
    .A1(_01572_),
    .S(_01417_),
    .X(_00783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15166_ (.A0(_00774_),
    .A1(_01321_),
    .S(_01263_),
    .X(_00775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15167_ (.A0(_00775_),
    .A1(_00850_),
    .S(_01287_),
    .X(_00776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15168_ (.A0(_02161_),
    .A1(_01943_),
    .S(_01363_),
    .X(_00777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15169_ (.A0(_00778_),
    .A1(_00763_),
    .S(_01593_),
    .X(_00779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15170_ (.A0(_00779_),
    .A1(_00762_),
    .S(_00822_),
    .X(_00780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15171_ (.A0(_00780_),
    .A1(_02584_),
    .S(_01596_),
    .X(_00781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15172_ (.A0(_00771_),
    .A1(_00843_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_00772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15173_ (.A0(_00843_),
    .A1(_00857_),
    .S(_01261_),
    .X(_00766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15174_ (.A0(_00766_),
    .A1(_02429_),
    .S(_01254_),
    .X(_00767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15175_ (.A0(_00767_),
    .A1(_02387_),
    .S(_01246_),
    .X(_00768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15176_ (.A0(_00768_),
    .A1(_02302_),
    .S(_01238_),
    .X(_00769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15177_ (.A0(_00769_),
    .A1(_02129_),
    .S(_01230_),
    .X(_00770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15178_ (.A0(_00760_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_00761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15179_ (.A0(_00758_),
    .A1(_00665_),
    .S(_00008_),
    .X(_00759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15180_ (.A0(_00756_),
    .A1(\design_top.IDATA[18] ),
    .S(_00008_),
    .X(_00757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15181_ (.A0(_00754_),
    .A1(\design_top.IDATA[17] ),
    .S(_00008_),
    .X(_00755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15182_ (.A0(_00752_),
    .A1(\design_top.IDATA[16] ),
    .S(_00008_),
    .X(_00753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15183_ (.A0(_00750_),
    .A1(\design_top.IDATA[15] ),
    .S(_00008_),
    .X(_00751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15184_ (.A0(_00748_),
    .A1(\design_top.IDATA[14] ),
    .S(_00008_),
    .X(_00749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15185_ (.A0(_00746_),
    .A1(\design_top.IDATA[13] ),
    .S(_00008_),
    .X(_00747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15186_ (.A0(_00743_),
    .A1(\design_top.IDATA[12] ),
    .S(_00008_),
    .X(_00744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15187_ (.A0(_00744_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15188_ (.A0(\design_top.ROMFF[11] ),
    .A1(\design_top.ROMFF2[11] ),
    .S(\design_top.HLT2 ),
    .X(_00718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15189_ (.A0(\design_top.ROMFF[29] ),
    .A1(\design_top.ROMFF2[29] ),
    .S(\design_top.HLT2 ),
    .X(_00701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15190_ (.A0(\design_top.ROMFF[28] ),
    .A1(\design_top.ROMFF2[28] ),
    .S(\design_top.HLT2 ),
    .X(_00697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15191_ (.A0(\design_top.ROMFF[27] ),
    .A1(\design_top.ROMFF2[27] ),
    .S(\design_top.HLT2 ),
    .X(_00693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15192_ (.A0(\design_top.ROMFF[26] ),
    .A1(\design_top.ROMFF2[26] ),
    .S(\design_top.HLT2 ),
    .X(_00689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15193_ (.A0(\design_top.ROMFF[25] ),
    .A1(\design_top.ROMFF2[25] ),
    .S(\design_top.HLT2 ),
    .X(_00685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15194_ (.A0(\design_top.ROMFF[24] ),
    .A1(\design_top.ROMFF2[24] ),
    .S(\design_top.HLT2 ),
    .X(_00681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15195_ (.A0(\design_top.ROMFF[19] ),
    .A1(\design_top.ROMFF2[19] ),
    .S(\design_top.HLT2 ),
    .X(_00665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15196_ (.A0(_01672_),
    .A1(_01364_),
    .S(_00821_),
    .X(_02469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15197_ (.A0(_01597_),
    .A1(_01367_),
    .S(_00821_),
    .X(_02468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15198_ (.A0(_02459_),
    .A1(_01320_),
    .S(_01263_),
    .X(_02460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15199_ (.A0(_02460_),
    .A1(_00864_),
    .S(_01287_),
    .X(_02461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15200_ (.A0(_02161_),
    .A1(_01900_),
    .S(_01363_),
    .X(_02462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15201_ (.A0(_02463_),
    .A1(_01338_),
    .S(_01593_),
    .X(_02464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15202_ (.A0(_02464_),
    .A1(_02447_),
    .S(_00822_),
    .X(_02465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15203_ (.A0(_02465_),
    .A1(_02466_),
    .S(_01596_),
    .X(_02467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15204_ (.A0(_02110_),
    .A1(_00843_),
    .S(_01230_),
    .X(_02456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15205_ (.A0(_02455_),
    .A1(_02456_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15206_ (.A0(_00857_),
    .A1(_00871_),
    .S(_01261_),
    .X(_02450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15207_ (.A0(_02450_),
    .A1(_02408_),
    .S(_01254_),
    .X(_02451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15208_ (.A0(_02451_),
    .A1(_02366_),
    .S(_01246_),
    .X(_02452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15209_ (.A0(_02452_),
    .A1(_02281_),
    .S(_01238_),
    .X(_02453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15210_ (.A0(_02453_),
    .A1(_02106_),
    .S(_01230_),
    .X(_02454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15211_ (.A0(_02438_),
    .A1(_01319_),
    .S(_01263_),
    .X(_02439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15212_ (.A0(_02439_),
    .A1(_00878_),
    .S(_01287_),
    .X(_02440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15213_ (.A0(_02161_),
    .A1(_01855_),
    .S(_01363_),
    .X(_02441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15214_ (.A0(_02442_),
    .A1(_01339_),
    .S(_01593_),
    .X(_02443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15215_ (.A0(_02443_),
    .A1(_02426_),
    .S(_00822_),
    .X(_02444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15216_ (.A0(_02444_),
    .A1(_02445_),
    .S(_01596_),
    .X(_02446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15217_ (.A0(_02084_),
    .A1(_00843_),
    .S(_01230_),
    .X(_02435_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15218_ (.A0(_02434_),
    .A1(_02435_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02436_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15219_ (.A0(_02429_),
    .A1(_02386_),
    .S(_01254_),
    .X(_02430_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15220_ (.A0(_02430_),
    .A1(_02344_),
    .S(_01246_),
    .X(_02431_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15221_ (.A0(_02431_),
    .A1(_02259_),
    .S(_01238_),
    .X(_02432_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15222_ (.A0(_02432_),
    .A1(_02080_),
    .S(_01230_),
    .X(_02433_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15223_ (.A0(_00871_),
    .A1(_00885_),
    .S(_01261_),
    .X(_02429_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15224_ (.A0(_02417_),
    .A1(_01318_),
    .S(_01263_),
    .X(_02418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15225_ (.A0(_02418_),
    .A1(_00892_),
    .S(_01287_),
    .X(_02419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15226_ (.A0(_02161_),
    .A1(_01811_),
    .S(_01363_),
    .X(_02420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15227_ (.A0(_02421_),
    .A1(_01340_),
    .S(_01593_),
    .X(_02422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15228_ (.A0(_02422_),
    .A1(_02404_),
    .S(_00822_),
    .X(_02423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15229_ (.A0(_02423_),
    .A1(_02424_),
    .S(_01596_),
    .X(_02425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15230_ (.A0(_02061_),
    .A1(_00843_),
    .S(_01230_),
    .X(_02414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15231_ (.A0(_02413_),
    .A1(_02414_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15232_ (.A0(_02408_),
    .A1(_02365_),
    .S(_01254_),
    .X(_02409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15233_ (.A0(_02409_),
    .A1(_02323_),
    .S(_01246_),
    .X(_02410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15234_ (.A0(_02410_),
    .A1(_02238_),
    .S(_01238_),
    .X(_02411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15235_ (.A0(_02411_),
    .A1(_02057_),
    .S(_01230_),
    .X(_02412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15236_ (.A0(_00885_),
    .A1(_00898_),
    .S(_01261_),
    .X(_02408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15237_ (.A0(_02395_),
    .A1(_01317_),
    .S(_01263_),
    .X(_02396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15238_ (.A0(_02396_),
    .A1(_00905_),
    .S(_01287_),
    .X(_02397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15239_ (.A0(_02161_),
    .A1(_01767_),
    .S(_01363_),
    .X(_02398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15240_ (.A0(_02399_),
    .A1(_01341_),
    .S(_01593_),
    .X(_02400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15241_ (.A0(_02400_),
    .A1(_02383_),
    .S(_00822_),
    .X(_02401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15242_ (.A0(_02401_),
    .A1(_02402_),
    .S(_01596_),
    .X(_02403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15243_ (.A0(_02037_),
    .A1(_00843_),
    .S(_01230_),
    .X(_02392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15244_ (.A0(_02391_),
    .A1(_02392_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15245_ (.A0(_02387_),
    .A1(_02301_),
    .S(_01246_),
    .X(_02388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15246_ (.A0(_02388_),
    .A1(_02216_),
    .S(_01238_),
    .X(_02389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15247_ (.A0(_02389_),
    .A1(_02033_),
    .S(_01230_),
    .X(_02390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15248_ (.A0(_02386_),
    .A1(_02343_),
    .S(_01254_),
    .X(_02387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15249_ (.A0(_00898_),
    .A1(_00912_),
    .S(_01261_),
    .X(_02386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15250_ (.A0(_02374_),
    .A1(_01316_),
    .S(_01263_),
    .X(_02375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15251_ (.A0(_02375_),
    .A1(_00919_),
    .S(_01287_),
    .X(_02376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15252_ (.A0(_02161_),
    .A1(_01716_),
    .S(_01363_),
    .X(_02377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15253_ (.A0(_02378_),
    .A1(_01342_),
    .S(_01593_),
    .X(_02379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15254_ (.A0(_02379_),
    .A1(_02361_),
    .S(_00822_),
    .X(_02380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15255_ (.A0(_02380_),
    .A1(_02381_),
    .S(_01596_),
    .X(_02382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15256_ (.A0(_02014_),
    .A1(_00843_),
    .S(_01230_),
    .X(_02371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15257_ (.A0(_02370_),
    .A1(_02371_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15258_ (.A0(_02366_),
    .A1(_02280_),
    .S(_01246_),
    .X(_02367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15259_ (.A0(_02367_),
    .A1(_02195_),
    .S(_01238_),
    .X(_02368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15260_ (.A0(_02368_),
    .A1(_02010_),
    .S(_01230_),
    .X(_02369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15261_ (.A0(_02365_),
    .A1(_02322_),
    .S(_01254_),
    .X(_02366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15262_ (.A0(_00912_),
    .A1(_00925_),
    .S(_01261_),
    .X(_02365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15263_ (.A0(_02352_),
    .A1(_01315_),
    .S(_01263_),
    .X(_02353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15264_ (.A0(_02353_),
    .A1(_00932_),
    .S(_01287_),
    .X(_02354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15265_ (.A0(_02161_),
    .A1(_01662_),
    .S(_01363_),
    .X(_02355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15266_ (.A0(_02356_),
    .A1(_01343_),
    .S(_01593_),
    .X(_02357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15267_ (.A0(_02357_),
    .A1(_02340_),
    .S(_00822_),
    .X(_02358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15268_ (.A0(_02358_),
    .A1(_02359_),
    .S(_01596_),
    .X(_02360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15269_ (.A0(_01990_),
    .A1(_00843_),
    .S(_01230_),
    .X(_02349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15270_ (.A0(_02348_),
    .A1(_02349_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15271_ (.A0(_02344_),
    .A1(_02258_),
    .S(_01246_),
    .X(_02345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15272_ (.A0(_02345_),
    .A1(_02173_),
    .S(_01238_),
    .X(_02346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15273_ (.A0(_02346_),
    .A1(_01986_),
    .S(_01230_),
    .X(_02347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15274_ (.A0(_02343_),
    .A1(_02300_),
    .S(_01254_),
    .X(_02344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15275_ (.A0(_00925_),
    .A1(_00939_),
    .S(_01261_),
    .X(_02343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15276_ (.A0(_02331_),
    .A1(_01314_),
    .S(_01263_),
    .X(_02332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15277_ (.A0(_02332_),
    .A1(_00946_),
    .S(_01287_),
    .X(_02333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15278_ (.A0(_02161_),
    .A1(_01585_),
    .S(_01363_),
    .X(_02334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15279_ (.A0(_02335_),
    .A1(_01344_),
    .S(_01593_),
    .X(_02336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15280_ (.A0(_02336_),
    .A1(_02318_),
    .S(_00822_),
    .X(_02337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15281_ (.A0(_02337_),
    .A1(_02338_),
    .S(_01596_),
    .X(_02339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15282_ (.A0(_01966_),
    .A1(_00843_),
    .S(_01230_),
    .X(_02328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15283_ (.A0(_02327_),
    .A1(_02328_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15284_ (.A0(_02323_),
    .A1(_02237_),
    .S(_01246_),
    .X(_02324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15285_ (.A0(_02324_),
    .A1(_02151_),
    .S(_01238_),
    .X(_02325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15286_ (.A0(_02325_),
    .A1(_01962_),
    .S(_01230_),
    .X(_02326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15287_ (.A0(_02322_),
    .A1(_02279_),
    .S(_01254_),
    .X(_02323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15288_ (.A0(_00939_),
    .A1(_00952_),
    .S(_01261_),
    .X(_02322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15289_ (.A0(_02309_),
    .A1(_01313_),
    .S(_01263_),
    .X(_02310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15290_ (.A0(_02310_),
    .A1(_00959_),
    .S(_01287_),
    .X(_02311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15291_ (.A0(_02161_),
    .A1(_01937_),
    .S(_01363_),
    .X(_02312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15292_ (.A0(_02313_),
    .A1(_01345_),
    .S(_01593_),
    .X(_02314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15293_ (.A0(_02314_),
    .A1(_02297_),
    .S(_00822_),
    .X(_02315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15294_ (.A0(_02315_),
    .A1(_02316_),
    .S(_01596_),
    .X(_02317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15295_ (.A0(_01926_),
    .A1(_00843_),
    .S(_01230_),
    .X(_02306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15296_ (.A0(_02305_),
    .A1(_02306_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15297_ (.A0(_02302_),
    .A1(_02128_),
    .S(_01238_),
    .X(_02303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15298_ (.A0(_02303_),
    .A1(_01918_),
    .S(_01230_),
    .X(_02304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15299_ (.A0(_02301_),
    .A1(_02215_),
    .S(_01246_),
    .X(_02302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15300_ (.A0(_02300_),
    .A1(_02257_),
    .S(_01254_),
    .X(_02301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15301_ (.A0(_00952_),
    .A1(_00966_),
    .S(_01261_),
    .X(_02300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15302_ (.A0(_02288_),
    .A1(_01312_),
    .S(_01263_),
    .X(_02289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15303_ (.A0(_02289_),
    .A1(_00973_),
    .S(_01287_),
    .X(_02290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15304_ (.A0(_02161_),
    .A1(_01895_),
    .S(_01363_),
    .X(_02291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15305_ (.A0(_02292_),
    .A1(_01346_),
    .S(_01593_),
    .X(_02293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15306_ (.A0(_02293_),
    .A1(_02275_),
    .S(_00822_),
    .X(_02294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15307_ (.A0(_02294_),
    .A1(_02295_),
    .S(_01596_),
    .X(_02296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15308_ (.A0(_01883_),
    .A1(_00843_),
    .S(_01230_),
    .X(_02285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15309_ (.A0(_02284_),
    .A1(_02285_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15310_ (.A0(_02281_),
    .A1(_02105_),
    .S(_01238_),
    .X(_02282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15311_ (.A0(_02282_),
    .A1(_01874_),
    .S(_01230_),
    .X(_02283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15312_ (.A0(_02280_),
    .A1(_02194_),
    .S(_01246_),
    .X(_02281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15313_ (.A0(_02279_),
    .A1(_02236_),
    .S(_01254_),
    .X(_02280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15314_ (.A0(_00966_),
    .A1(_00979_),
    .S(_01261_),
    .X(_02279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15315_ (.A0(_02266_),
    .A1(_01311_),
    .S(_01263_),
    .X(_02267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15316_ (.A0(_02267_),
    .A1(_00986_),
    .S(_01287_),
    .X(_02268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15317_ (.A0(_02161_),
    .A1(_01850_),
    .S(_01363_),
    .X(_02269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15318_ (.A0(_02270_),
    .A1(_01347_),
    .S(_01593_),
    .X(_02271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15319_ (.A0(_02271_),
    .A1(_02254_),
    .S(_00822_),
    .X(_02272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15320_ (.A0(_02272_),
    .A1(_02273_),
    .S(_01596_),
    .X(_02274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15321_ (.A0(_01838_),
    .A1(_00843_),
    .S(_01230_),
    .X(_02263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15322_ (.A0(_02262_),
    .A1(_02263_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15323_ (.A0(_02259_),
    .A1(_02079_),
    .S(_01238_),
    .X(_02260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15324_ (.A0(_02260_),
    .A1(_01829_),
    .S(_01230_),
    .X(_02261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15325_ (.A0(_02258_),
    .A1(_02172_),
    .S(_01246_),
    .X(_02259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15326_ (.A0(_02257_),
    .A1(_02214_),
    .S(_01254_),
    .X(_02258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15327_ (.A0(_00979_),
    .A1(_00993_),
    .S(_01261_),
    .X(_02257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15328_ (.A0(_02245_),
    .A1(_01310_),
    .S(_01263_),
    .X(_02246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15329_ (.A0(_02246_),
    .A1(_01000_),
    .S(_01287_),
    .X(_02247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15330_ (.A0(_02161_),
    .A1(_01806_),
    .S(_01363_),
    .X(_02248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15331_ (.A0(_02249_),
    .A1(_01348_),
    .S(_01593_),
    .X(_02250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15332_ (.A0(_02250_),
    .A1(_02232_),
    .S(_00822_),
    .X(_02251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15333_ (.A0(_02251_),
    .A1(_02252_),
    .S(_01596_),
    .X(_02253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15334_ (.A0(_01795_),
    .A1(_00843_),
    .S(_01230_),
    .X(_02242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15335_ (.A0(_02241_),
    .A1(_02242_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15336_ (.A0(_02238_),
    .A1(_02056_),
    .S(_01238_),
    .X(_02239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15337_ (.A0(_02239_),
    .A1(_01786_),
    .S(_01230_),
    .X(_02240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15338_ (.A0(_02237_),
    .A1(_02150_),
    .S(_01246_),
    .X(_02238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15339_ (.A0(_02236_),
    .A1(_02193_),
    .S(_01254_),
    .X(_02237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15340_ (.A0(_00993_),
    .A1(_01006_),
    .S(_01261_),
    .X(_02236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15341_ (.A0(_02223_),
    .A1(_01309_),
    .S(_01263_),
    .X(_02224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15342_ (.A0(_02224_),
    .A1(_01013_),
    .S(_01287_),
    .X(_02225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15343_ (.A0(_02161_),
    .A1(_01762_),
    .S(_01363_),
    .X(_02226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15344_ (.A0(_02227_),
    .A1(_01349_),
    .S(_01593_),
    .X(_02228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15345_ (.A0(_02228_),
    .A1(_02211_),
    .S(_00822_),
    .X(_02229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15346_ (.A0(_02229_),
    .A1(_02230_),
    .S(_01596_),
    .X(_02231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15347_ (.A0(_01751_),
    .A1(_00843_),
    .S(_01230_),
    .X(_02220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15348_ (.A0(_02219_),
    .A1(_02220_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15349_ (.A0(_02216_),
    .A1(_02032_),
    .S(_01238_),
    .X(_02217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15350_ (.A0(_02217_),
    .A1(_01734_),
    .S(_01230_),
    .X(_02218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15351_ (.A0(_02215_),
    .A1(_02127_),
    .S(_01246_),
    .X(_02216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15352_ (.A0(_02214_),
    .A1(_02171_),
    .S(_01254_),
    .X(_02215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15353_ (.A0(_01006_),
    .A1(_01020_),
    .S(_01261_),
    .X(_02214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15354_ (.A0(_02202_),
    .A1(_01308_),
    .S(_01263_),
    .X(_02203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15355_ (.A0(_02203_),
    .A1(_01027_),
    .S(_01287_),
    .X(_02204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15356_ (.A0(_02161_),
    .A1(_01711_),
    .S(_01363_),
    .X(_02205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15357_ (.A0(_02206_),
    .A1(_01350_),
    .S(_01593_),
    .X(_02207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15358_ (.A0(_02207_),
    .A1(_02189_),
    .S(_00822_),
    .X(_02208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15359_ (.A0(_02208_),
    .A1(_02209_),
    .S(_01596_),
    .X(_02210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15360_ (.A0(_01699_),
    .A1(_00843_),
    .S(_01230_),
    .X(_02199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15361_ (.A0(_02198_),
    .A1(_02199_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15362_ (.A0(_02195_),
    .A1(_02009_),
    .S(_01238_),
    .X(_02196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15363_ (.A0(_02196_),
    .A1(_01681_),
    .S(_01230_),
    .X(_02197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15364_ (.A0(_02194_),
    .A1(_02104_),
    .S(_01246_),
    .X(_02195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15365_ (.A0(_02193_),
    .A1(_02149_),
    .S(_01254_),
    .X(_02194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15366_ (.A0(_01020_),
    .A1(_01048_),
    .S(_01261_),
    .X(_02193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15367_ (.A0(_02180_),
    .A1(_01307_),
    .S(_01263_),
    .X(_02181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15368_ (.A0(_02181_),
    .A1(_01055_),
    .S(_01287_),
    .X(_02182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15369_ (.A0(_02161_),
    .A1(_01656_),
    .S(_01363_),
    .X(_02183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15370_ (.A0(_02184_),
    .A1(_01351_),
    .S(_01593_),
    .X(_02185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15371_ (.A0(_02185_),
    .A1(_02168_),
    .S(_00822_),
    .X(_02186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15372_ (.A0(_02186_),
    .A1(_02187_),
    .S(_01596_),
    .X(_02188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15373_ (.A0(_01645_),
    .A1(_00843_),
    .S(_01230_),
    .X(_02177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15374_ (.A0(_02176_),
    .A1(_02177_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15375_ (.A0(_02173_),
    .A1(_01985_),
    .S(_01238_),
    .X(_02174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15376_ (.A0(_02174_),
    .A1(_01611_),
    .S(_01230_),
    .X(_02175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15377_ (.A0(_02172_),
    .A1(_02078_),
    .S(_01246_),
    .X(_02173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15378_ (.A0(_02171_),
    .A1(_02126_),
    .S(_01254_),
    .X(_02172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15379_ (.A0(_01048_),
    .A1(_01062_),
    .S(_01261_),
    .X(_02171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15380_ (.A0(_02158_),
    .A1(_01306_),
    .S(_01263_),
    .X(_02159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15381_ (.A0(_02159_),
    .A1(_01069_),
    .S(_01287_),
    .X(_02160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15382_ (.A0(_02161_),
    .A1(_01578_),
    .S(_01363_),
    .X(_02162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15383_ (.A0(_02163_),
    .A1(_01352_),
    .S(_01593_),
    .X(_02164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15384_ (.A0(_02164_),
    .A1(_02145_),
    .S(_00822_),
    .X(_02165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15385_ (.A0(_02165_),
    .A1(_02166_),
    .S(_01596_),
    .X(_02167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15386_ (.A0(_01562_),
    .A1(_00843_),
    .S(_01230_),
    .X(_02155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15387_ (.A0(_02154_),
    .A1(_02155_),
    .S(\design_top.core0.FCT7[5] ),
    .X(_02156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15388_ (.A0(_02151_),
    .A1(_01961_),
    .S(_01238_),
    .X(_02152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15389_ (.A0(_02152_),
    .A1(_01529_),
    .S(_01230_),
    .X(_02153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15390_ (.A0(_02150_),
    .A1(_02055_),
    .S(_01246_),
    .X(_02151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15391_ (.A0(_02149_),
    .A1(_02103_),
    .S(_01254_),
    .X(_02150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15392_ (.A0(_01062_),
    .A1(_01075_),
    .S(_01261_),
    .X(_02149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15393_ (.A0(_02135_),
    .A1(_01305_),
    .S(_01263_),
    .X(_02136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15394_ (.A0(_02136_),
    .A1(_01082_),
    .S(_01287_),
    .X(_02137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15395_ (.A0(_02138_),
    .A1(_01946_),
    .S(_01363_),
    .X(_02139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15396_ (.A0(_02140_),
    .A1(_01353_),
    .S(_01593_),
    .X(_02141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15397_ (.A0(_02141_),
    .A1(_02123_),
    .S(_00822_),
    .X(_02142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15398_ (.A0(_02142_),
    .A1(_02143_),
    .S(_01596_),
    .X(_02144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15399_ (.A0(_01943_),
    .A1(_01946_),
    .S(_01364_),
    .X(_02138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15400_ (.A0(_01921_),
    .A1(_01923_),
    .S(_01238_),
    .X(_02131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15401_ (.A0(_02128_),
    .A1(_01917_),
    .S(_01238_),
    .X(_02129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15402_ (.A0(_02127_),
    .A1(_02031_),
    .S(_01246_),
    .X(_02128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15403_ (.A0(_02126_),
    .A1(_02077_),
    .S(_01254_),
    .X(_02127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15404_ (.A0(_01075_),
    .A1(_01089_),
    .S(_01261_),
    .X(_02126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15405_ (.A0(_02113_),
    .A1(_01304_),
    .S(_01263_),
    .X(_02114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15406_ (.A0(_02114_),
    .A1(_01096_),
    .S(_01287_),
    .X(_02115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15407_ (.A0(_01900_),
    .A1(_01903_),
    .S(_01364_),
    .X(_02116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15408_ (.A0(_02116_),
    .A1(_01903_),
    .S(_01363_),
    .X(_02117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15409_ (.A0(_02118_),
    .A1(_01354_),
    .S(_01593_),
    .X(_02119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15410_ (.A0(_02119_),
    .A1(_02099_),
    .S(_00822_),
    .X(_02120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15411_ (.A0(_02120_),
    .A1(_02121_),
    .S(_01596_),
    .X(_02122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15412_ (.A0(_01882_),
    .A1(_00843_),
    .S(_01238_),
    .X(_02110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15413_ (.A0(_01877_),
    .A1(_01879_),
    .S(_01238_),
    .X(_02108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15414_ (.A0(_02105_),
    .A1(_01873_),
    .S(_01238_),
    .X(_02106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15415_ (.A0(_02104_),
    .A1(_02008_),
    .S(_01246_),
    .X(_02105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15416_ (.A0(_02103_),
    .A1(_02054_),
    .S(_01254_),
    .X(_02104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15417_ (.A0(_01089_),
    .A1(_01102_),
    .S(_01261_),
    .X(_02103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15418_ (.A0(_02087_),
    .A1(_01303_),
    .S(_01263_),
    .X(_02088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15419_ (.A0(_02088_),
    .A1(_01109_),
    .S(_01287_),
    .X(_02089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15420_ (.A0(_01855_),
    .A1(_01858_),
    .S(_01364_),
    .X(_02090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15421_ (.A0(_02090_),
    .A1(_01858_),
    .S(_01363_),
    .X(_02091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15422_ (.A0(_02092_),
    .A1(_01355_),
    .S(_01593_),
    .X(_02093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15423_ (.A0(_02093_),
    .A1(_02074_),
    .S(_00822_),
    .X(_02094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15424_ (.A0(_02094_),
    .A1(_02095_),
    .S(_01596_),
    .X(_02096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15425_ (.A0(_01837_),
    .A1(_00843_),
    .S(_01238_),
    .X(_02084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15426_ (.A0(_01832_),
    .A1(_01834_),
    .S(_01238_),
    .X(_02082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15427_ (.A0(_02079_),
    .A1(_01828_),
    .S(_01238_),
    .X(_02080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15428_ (.A0(_02078_),
    .A1(_01984_),
    .S(_01246_),
    .X(_02079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15429_ (.A0(_02077_),
    .A1(_02030_),
    .S(_01254_),
    .X(_02078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15430_ (.A0(_01102_),
    .A1(_01116_),
    .S(_01261_),
    .X(_02077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15431_ (.A0(_02064_),
    .A1(_01302_),
    .S(_01263_),
    .X(_02065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15432_ (.A0(_02065_),
    .A1(_01123_),
    .S(_01287_),
    .X(_02066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15433_ (.A0(_01811_),
    .A1(_01814_),
    .S(_01364_),
    .X(_02067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15434_ (.A0(_02067_),
    .A1(_01814_),
    .S(_01363_),
    .X(_02068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15435_ (.A0(_02069_),
    .A1(_01356_),
    .S(_01593_),
    .X(_02070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15436_ (.A0(_02070_),
    .A1(_02050_),
    .S(_00822_),
    .X(_02071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15437_ (.A0(_02071_),
    .A1(_02072_),
    .S(_01596_),
    .X(_02073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15438_ (.A0(_01794_),
    .A1(_00843_),
    .S(_01238_),
    .X(_02061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15439_ (.A0(_01789_),
    .A1(_01791_),
    .S(_01238_),
    .X(_02059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15440_ (.A0(_02056_),
    .A1(_01785_),
    .S(_01238_),
    .X(_02057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15441_ (.A0(_02055_),
    .A1(_01960_),
    .S(_01246_),
    .X(_02056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15442_ (.A0(_02054_),
    .A1(_02007_),
    .S(_01254_),
    .X(_02055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15443_ (.A0(_01116_),
    .A1(_01540_),
    .S(_01261_),
    .X(_02054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15444_ (.A0(_02040_),
    .A1(_01301_),
    .S(_01263_),
    .X(_02041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15445_ (.A0(_02041_),
    .A1(_01135_),
    .S(_01287_),
    .X(_02042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15446_ (.A0(_01767_),
    .A1(_01770_),
    .S(_01364_),
    .X(_02043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15447_ (.A0(_02043_),
    .A1(_01770_),
    .S(_01363_),
    .X(_02044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15448_ (.A0(_02045_),
    .A1(_01357_),
    .S(_01593_),
    .X(_02046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15449_ (.A0(_02046_),
    .A1(_02027_),
    .S(_00822_),
    .X(_02047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15450_ (.A0(_02047_),
    .A1(_02048_),
    .S(_01596_),
    .X(_02049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15451_ (.A0(_01750_),
    .A1(_00843_),
    .S(_01238_),
    .X(_02037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15452_ (.A0(_01741_),
    .A1(_01745_),
    .S(_01238_),
    .X(_02035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15453_ (.A0(_02032_),
    .A1(_01733_),
    .S(_01238_),
    .X(_02033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15454_ (.A0(_02031_),
    .A1(_01916_),
    .S(_01246_),
    .X(_02032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15455_ (.A0(_02030_),
    .A1(_01983_),
    .S(_01254_),
    .X(_02031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15456_ (.A0(_01540_),
    .A1(_01142_),
    .S(_01261_),
    .X(_02030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15457_ (.A0(_02017_),
    .A1(_01300_),
    .S(_01263_),
    .X(_02018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15458_ (.A0(_02018_),
    .A1(_01149_),
    .S(_01287_),
    .X(_02019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15459_ (.A0(_01716_),
    .A1(_01719_),
    .S(_01364_),
    .X(_02020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15460_ (.A0(_02020_),
    .A1(_01719_),
    .S(_01363_),
    .X(_02021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15461_ (.A0(_02022_),
    .A1(_01358_),
    .S(_01593_),
    .X(_02023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15462_ (.A0(_02023_),
    .A1(_02003_),
    .S(_00822_),
    .X(_02024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15463_ (.A0(_02024_),
    .A1(_02025_),
    .S(_01596_),
    .X(_02026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15464_ (.A0(_01698_),
    .A1(_00843_),
    .S(_01238_),
    .X(_02014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15465_ (.A0(_01688_),
    .A1(_01692_),
    .S(_01238_),
    .X(_02012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15466_ (.A0(_02009_),
    .A1(_01680_),
    .S(_01238_),
    .X(_02010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15467_ (.A0(_02008_),
    .A1(_01872_),
    .S(_01246_),
    .X(_02009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15468_ (.A0(_02007_),
    .A1(_01959_),
    .S(_01254_),
    .X(_02008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15469_ (.A0(_01142_),
    .A1(_01156_),
    .S(_01261_),
    .X(_02007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15470_ (.A0(_01993_),
    .A1(_01299_),
    .S(_01263_),
    .X(_01994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15471_ (.A0(_01994_),
    .A1(_01163_),
    .S(_01287_),
    .X(_01995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15472_ (.A0(_01662_),
    .A1(_01665_),
    .S(_01364_),
    .X(_01996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15473_ (.A0(_01996_),
    .A1(_01665_),
    .S(_01363_),
    .X(_01997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15474_ (.A0(_01998_),
    .A1(_01359_),
    .S(_01593_),
    .X(_01999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15475_ (.A0(_01999_),
    .A1(_01980_),
    .S(_00822_),
    .X(_02000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15476_ (.A0(_02000_),
    .A1(_02001_),
    .S(_01596_),
    .X(_02002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15477_ (.A0(_01644_),
    .A1(_00843_),
    .S(_01238_),
    .X(_01990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15478_ (.A0(_01626_),
    .A1(_01634_),
    .S(_01238_),
    .X(_01988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15479_ (.A0(_01985_),
    .A1(_01610_),
    .S(_01238_),
    .X(_01986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15480_ (.A0(_01984_),
    .A1(_01827_),
    .S(_01246_),
    .X(_01985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15481_ (.A0(_01983_),
    .A1(_01915_),
    .S(_01254_),
    .X(_01984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15482_ (.A0(_01156_),
    .A1(_01171_),
    .S(_01261_),
    .X(_01983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15483_ (.A0(_01969_),
    .A1(_01298_),
    .S(_01263_),
    .X(_01970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15484_ (.A0(_01970_),
    .A1(_01178_),
    .S(_01287_),
    .X(_01971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15485_ (.A0(_01585_),
    .A1(_01588_),
    .S(_01364_),
    .X(_01972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15486_ (.A0(_01972_),
    .A1(_01588_),
    .S(_01363_),
    .X(_01973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15487_ (.A0(_01975_),
    .A1(_01360_),
    .S(_01593_),
    .X(_01976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15488_ (.A0(_01976_),
    .A1(_01955_),
    .S(_00822_),
    .X(_01977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15489_ (.A0(_01977_),
    .A1(_01978_),
    .S(_01596_),
    .X(_01979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15490_ (.A0(_01561_),
    .A1(_00843_),
    .S(_01238_),
    .X(_01966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15491_ (.A0(_01546_),
    .A1(_01554_),
    .S(_01238_),
    .X(_01964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15492_ (.A0(_01961_),
    .A1(_01528_),
    .S(_01238_),
    .X(_01962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15493_ (.A0(_01960_),
    .A1(_01784_),
    .S(_01246_),
    .X(_01961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15494_ (.A0(_01959_),
    .A1(_01871_),
    .S(_01254_),
    .X(_01960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15495_ (.A0(_01171_),
    .A1(_01184_),
    .S(_01261_),
    .X(_01959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15496_ (.A0(_01929_),
    .A1(_01297_),
    .S(_01263_),
    .X(_01930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15497_ (.A0(_01930_),
    .A1(_01191_),
    .S(_01287_),
    .X(_01931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15498_ (.A0(_01937_),
    .A1(_01934_),
    .S(_01364_),
    .X(_01938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15499_ (.A0(_01938_),
    .A1(_01934_),
    .S(_01363_),
    .X(_01939_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15500_ (.A0(_01950_),
    .A1(_01361_),
    .S(_01593_),
    .X(_01951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15501_ (.A0(_01951_),
    .A1(_01912_),
    .S(_00822_),
    .X(_01952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15502_ (.A0(_01952_),
    .A1(_01953_),
    .S(_01596_),
    .X(_01954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15503_ (.A0(_01934_),
    .A1(_01946_),
    .S(_01378_),
    .X(_01947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15504_ (.A0(_01947_),
    .A1(_01937_),
    .S(_01423_),
    .X(_01948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15505_ (.A0(_01948_),
    .A1(_01943_),
    .S(_01372_),
    .X(_01949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15506_ (.A0(_01944_),
    .A1(_01945_),
    .S(\design_top.XADDR[31] ),
    .X(_01946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15507_ (.A0(_01941_),
    .A1(_01376_),
    .S(_01573_),
    .X(_01942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15508_ (.A0(_01940_),
    .A1(_01942_),
    .S(\design_top.XADDR[31] ),
    .X(_01943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15509_ (.A0(_01935_),
    .A1(_01936_),
    .S(\design_top.XADDR[31] ),
    .X(_01937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15510_ (.A0(_01932_),
    .A1(_01933_),
    .S(\design_top.XADDR[31] ),
    .X(_01934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15511_ (.A0(_01923_),
    .A1(_00843_),
    .S(_01238_),
    .X(_01926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15512_ (.A0(_01923_),
    .A1(_01924_),
    .S(_01238_),
    .X(_01925_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15513_ (.A0(_01744_),
    .A1(_01746_),
    .S(_01246_),
    .X(_01923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15514_ (.A0(_01737_),
    .A1(_01739_),
    .S(_01246_),
    .X(_01920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15515_ (.A0(_01920_),
    .A1(_01921_),
    .S(_01238_),
    .X(_01922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15516_ (.A0(_01740_),
    .A1(_01743_),
    .S(_01246_),
    .X(_01921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15517_ (.A0(_01916_),
    .A1(_01732_),
    .S(_01246_),
    .X(_01917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15518_ (.A0(_01915_),
    .A1(_01826_),
    .S(_01254_),
    .X(_01916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15519_ (.A0(_01184_),
    .A1(_01198_),
    .S(_01261_),
    .X(_01915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15520_ (.A0(_01886_),
    .A1(_01296_),
    .S(_01263_),
    .X(_01887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15521_ (.A0(_01887_),
    .A1(_01205_),
    .S(_01287_),
    .X(_01888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15522_ (.A0(_01891_),
    .A1(_01903_),
    .S(_01378_),
    .X(_01904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15523_ (.A0(_01904_),
    .A1(_01895_),
    .S(_01423_),
    .X(_01905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15524_ (.A0(_01905_),
    .A1(_01900_),
    .S(_01372_),
    .X(_01906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15525_ (.A0(_01895_),
    .A1(_01891_),
    .S(_01364_),
    .X(_01896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15526_ (.A0(_01896_),
    .A1(_01891_),
    .S(_01363_),
    .X(_01897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15527_ (.A0(_01907_),
    .A1(_01336_),
    .S(_01593_),
    .X(_01908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15528_ (.A0(_01908_),
    .A1(_01867_),
    .S(_00822_),
    .X(_01909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15529_ (.A0(_01909_),
    .A1(_01910_),
    .S(_01596_),
    .X(_01911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15530_ (.A0(_01901_),
    .A1(_01902_),
    .S(\design_top.XADDR[31] ),
    .X(_01903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15531_ (.A0(_01898_),
    .A1(_01899_),
    .S(\design_top.XADDR[31] ),
    .X(_01900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15532_ (.A0(_01582_),
    .A1(_01893_),
    .S(\design_top.XADDR[3] ),
    .X(_01894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15533_ (.A0(_01892_),
    .A1(_01894_),
    .S(\design_top.XADDR[31] ),
    .X(_01895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15534_ (.A0(_01889_),
    .A1(_01890_),
    .S(\design_top.XADDR[31] ),
    .X(_01891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15535_ (.A0(_01879_),
    .A1(_01882_),
    .S(_01238_),
    .X(_01883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15536_ (.A0(_01697_),
    .A1(_00843_),
    .S(_01246_),
    .X(_01882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15537_ (.A0(_01879_),
    .A1(_01880_),
    .S(_01238_),
    .X(_01881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15538_ (.A0(_01691_),
    .A1(_01693_),
    .S(_01246_),
    .X(_01879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15539_ (.A0(_01684_),
    .A1(_01686_),
    .S(_01246_),
    .X(_01876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15540_ (.A0(_01876_),
    .A1(_01877_),
    .S(_01238_),
    .X(_01878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15541_ (.A0(_01687_),
    .A1(_01690_),
    .S(_01246_),
    .X(_01877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15542_ (.A0(_01872_),
    .A1(_01679_),
    .S(_01246_),
    .X(_01873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15543_ (.A0(_01871_),
    .A1(_01783_),
    .S(_01254_),
    .X(_01872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15544_ (.A0(_01198_),
    .A1(_01534_),
    .S(_01261_),
    .X(_01871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15545_ (.A0(_01841_),
    .A1(_01295_),
    .S(_01263_),
    .X(_01842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15546_ (.A0(_01842_),
    .A1(_01217_),
    .S(_01287_),
    .X(_01843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15547_ (.A0(_01846_),
    .A1(_01858_),
    .S(_01378_),
    .X(_01859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15548_ (.A0(_01859_),
    .A1(_01850_),
    .S(_01423_),
    .X(_01860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15549_ (.A0(_01860_),
    .A1(_01855_),
    .S(_01372_),
    .X(_01861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15550_ (.A0(_01850_),
    .A1(_01846_),
    .S(_01364_),
    .X(_01851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15551_ (.A0(_01851_),
    .A1(_01846_),
    .S(_01363_),
    .X(_01852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15552_ (.A0(_01862_),
    .A1(_01334_),
    .S(_01593_),
    .X(_01863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15553_ (.A0(_01863_),
    .A1(_01823_),
    .S(_00822_),
    .X(_01864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15554_ (.A0(_01864_),
    .A1(_01865_),
    .S(_01596_),
    .X(_01866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15555_ (.A0(_01856_),
    .A1(_01857_),
    .S(\design_top.XADDR[31] ),
    .X(_01858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15556_ (.A0(_01853_),
    .A1(_01854_),
    .S(\design_top.XADDR[31] ),
    .X(_01855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15557_ (.A0(_01582_),
    .A1(_01848_),
    .S(\design_top.XADDR[3] ),
    .X(_01849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15558_ (.A0(_01847_),
    .A1(_01849_),
    .S(\design_top.XADDR[31] ),
    .X(_01850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15559_ (.A0(_01844_),
    .A1(_01845_),
    .S(\design_top.XADDR[31] ),
    .X(_01846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15560_ (.A0(_01834_),
    .A1(_01837_),
    .S(_01238_),
    .X(_01838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15561_ (.A0(_01643_),
    .A1(_00843_),
    .S(_01246_),
    .X(_01837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15562_ (.A0(_01834_),
    .A1(_01835_),
    .S(_01238_),
    .X(_01836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15563_ (.A0(_01633_),
    .A1(_01637_),
    .S(_01246_),
    .X(_01834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15564_ (.A0(_01618_),
    .A1(_01622_),
    .S(_01246_),
    .X(_01831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15565_ (.A0(_01831_),
    .A1(_01832_),
    .S(_01238_),
    .X(_01833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15566_ (.A0(_01625_),
    .A1(_01630_),
    .S(_01246_),
    .X(_01832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15567_ (.A0(_01827_),
    .A1(_01609_),
    .S(_01246_),
    .X(_01828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15568_ (.A0(_01826_),
    .A1(_01731_),
    .S(_01254_),
    .X(_01827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15569_ (.A0(_01534_),
    .A1(_01224_),
    .S(_01261_),
    .X(_01826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15570_ (.A0(_01798_),
    .A1(_01294_),
    .S(_01263_),
    .X(_01799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15571_ (.A0(_01799_),
    .A1(_01231_),
    .S(_01287_),
    .X(_01800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15572_ (.A0(_01803_),
    .A1(_01814_),
    .S(_01378_),
    .X(_01815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15573_ (.A0(_01815_),
    .A1(_01806_),
    .S(_01423_),
    .X(_01816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15574_ (.A0(_01816_),
    .A1(_01811_),
    .S(_01372_),
    .X(_01817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15575_ (.A0(_01806_),
    .A1(_01803_),
    .S(_01364_),
    .X(_01807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15576_ (.A0(_01807_),
    .A1(_01803_),
    .S(_01363_),
    .X(_01808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15577_ (.A0(_01818_),
    .A1(_01332_),
    .S(_01593_),
    .X(_01819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15578_ (.A0(_01819_),
    .A1(_01779_),
    .S(_00822_),
    .X(_01820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15579_ (.A0(_01820_),
    .A1(_01821_),
    .S(_01596_),
    .X(_01822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15580_ (.A0(_01812_),
    .A1(_01813_),
    .S(\design_top.XADDR[31] ),
    .X(_01814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15581_ (.A0(_01809_),
    .A1(_01810_),
    .S(\design_top.XADDR[31] ),
    .X(_01811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15582_ (.A0(_01804_),
    .A1(_01805_),
    .S(\design_top.XADDR[31] ),
    .X(_01806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15583_ (.A0(_01801_),
    .A1(_01802_),
    .S(\design_top.XADDR[31] ),
    .X(_01803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15584_ (.A0(_01791_),
    .A1(_01794_),
    .S(_01238_),
    .X(_01795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15585_ (.A0(_01560_),
    .A1(_00843_),
    .S(_01246_),
    .X(_01794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15586_ (.A0(_01791_),
    .A1(_01792_),
    .S(_01238_),
    .X(_01793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15587_ (.A0(_01553_),
    .A1(_01557_),
    .S(_01246_),
    .X(_01791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15588_ (.A0(_01537_),
    .A1(_01542_),
    .S(_01246_),
    .X(_01788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15589_ (.A0(_01788_),
    .A1(_01789_),
    .S(_01238_),
    .X(_01790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15590_ (.A0(_01545_),
    .A1(_01550_),
    .S(_01246_),
    .X(_01789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15591_ (.A0(_01784_),
    .A1(_01527_),
    .S(_01246_),
    .X(_01785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15592_ (.A0(_01783_),
    .A1(_01678_),
    .S(_01254_),
    .X(_01784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15593_ (.A0(_01224_),
    .A1(_01232_),
    .S(_01261_),
    .X(_01783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15594_ (.A0(_01754_),
    .A1(_01293_),
    .S(_01263_),
    .X(_01755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15595_ (.A0(_01755_),
    .A1(_01239_),
    .S(_01287_),
    .X(_01756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15596_ (.A0(_01759_),
    .A1(_01770_),
    .S(_01378_),
    .X(_01771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15597_ (.A0(_01771_),
    .A1(_01762_),
    .S(_01423_),
    .X(_01772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15598_ (.A0(_01772_),
    .A1(_01767_),
    .S(_01372_),
    .X(_01773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15599_ (.A0(_01762_),
    .A1(_01759_),
    .S(_01364_),
    .X(_01763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15600_ (.A0(_01763_),
    .A1(_01759_),
    .S(_01363_),
    .X(_01764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15601_ (.A0(_01774_),
    .A1(_00811_),
    .S(_01593_),
    .X(_01775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15602_ (.A0(_01775_),
    .A1(_01728_),
    .S(_00822_),
    .X(_01776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15603_ (.A0(_01776_),
    .A1(_01777_),
    .S(_01596_),
    .X(_01778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15604_ (.A0(_01768_),
    .A1(_01769_),
    .S(\design_top.XADDR[31] ),
    .X(_01770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15605_ (.A0(_01765_),
    .A1(_01766_),
    .S(\design_top.XADDR[31] ),
    .X(_01767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15606_ (.A0(_01760_),
    .A1(_01761_),
    .S(\design_top.XADDR[31] ),
    .X(_01762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15607_ (.A0(_01757_),
    .A1(_01758_),
    .S(\design_top.XADDR[31] ),
    .X(_01759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15608_ (.A0(_01745_),
    .A1(_01750_),
    .S(_01238_),
    .X(_01751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15609_ (.A0(_01746_),
    .A1(_00843_),
    .S(_01246_),
    .X(_01750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15610_ (.A0(_01745_),
    .A1(_01748_),
    .S(_01238_),
    .X(_01749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15611_ (.A0(_01746_),
    .A1(_01747_),
    .S(_01246_),
    .X(_01748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15612_ (.A0(_01636_),
    .A1(_01638_),
    .S(_01254_),
    .X(_01746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15613_ (.A0(_01743_),
    .A1(_01744_),
    .S(_01246_),
    .X(_01745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15614_ (.A0(_01632_),
    .A1(_01635_),
    .S(_01254_),
    .X(_01744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15615_ (.A0(_01629_),
    .A1(_01631_),
    .S(_01254_),
    .X(_01743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15616_ (.A0(_01614_),
    .A1(_01616_),
    .S(_01254_),
    .X(_01736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15617_ (.A0(_01736_),
    .A1(_01737_),
    .S(_01246_),
    .X(_01738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15618_ (.A0(_01738_),
    .A1(_01741_),
    .S(_01238_),
    .X(_01742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15619_ (.A0(_01739_),
    .A1(_01740_),
    .S(_01246_),
    .X(_01741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15620_ (.A0(_01624_),
    .A1(_01628_),
    .S(_01254_),
    .X(_01740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15621_ (.A0(_01621_),
    .A1(_01623_),
    .S(_01254_),
    .X(_01739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15622_ (.A0(_01617_),
    .A1(_01620_),
    .S(_01254_),
    .X(_01737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15623_ (.A0(_01731_),
    .A1(_01608_),
    .S(_01254_),
    .X(_01732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15624_ (.A0(_01232_),
    .A1(_00793_),
    .S(_01261_),
    .X(_01731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15625_ (.A0(_01702_),
    .A1(_01292_),
    .S(_01263_),
    .X(_01703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15626_ (.A0(_01703_),
    .A1(_01247_),
    .S(_01287_),
    .X(_01704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15627_ (.A0(_01707_),
    .A1(_01719_),
    .S(_01378_),
    .X(_01720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15628_ (.A0(_01720_),
    .A1(_01711_),
    .S(_01423_),
    .X(_01721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15629_ (.A0(_01721_),
    .A1(_01716_),
    .S(_01372_),
    .X(_01722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15630_ (.A0(_01711_),
    .A1(_01707_),
    .S(_01364_),
    .X(_01712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15631_ (.A0(_01712_),
    .A1(_01707_),
    .S(_01363_),
    .X(_01713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15632_ (.A0(_01723_),
    .A1(_00819_),
    .S(_01593_),
    .X(_01724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15633_ (.A0(_01724_),
    .A1(_01674_),
    .S(_00822_),
    .X(_01725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15634_ (.A0(_01725_),
    .A1(_01726_),
    .S(_01596_),
    .X(_01727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15635_ (.A0(_01717_),
    .A1(_01718_),
    .S(\design_top.XADDR[31] ),
    .X(_01719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15636_ (.A0(_01714_),
    .A1(_01715_),
    .S(\design_top.XADDR[31] ),
    .X(_01716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15637_ (.A0(_01582_),
    .A1(_01709_),
    .S(\design_top.XADDR[3] ),
    .X(_01710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15638_ (.A0(_01708_),
    .A1(_01710_),
    .S(\design_top.XADDR[31] ),
    .X(_01711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15639_ (.A0(_01705_),
    .A1(_01706_),
    .S(\design_top.XADDR[31] ),
    .X(_01707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15640_ (.A0(_01692_),
    .A1(_01698_),
    .S(_01238_),
    .X(_01699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15641_ (.A0(_01693_),
    .A1(_01697_),
    .S(_01246_),
    .X(_01698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15642_ (.A0(_01559_),
    .A1(_00843_),
    .S(_01254_),
    .X(_01697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15643_ (.A0(_01692_),
    .A1(_01695_),
    .S(_01238_),
    .X(_01696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15644_ (.A0(_01693_),
    .A1(_01694_),
    .S(_01246_),
    .X(_01695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15645_ (.A0(_01556_),
    .A1(_01558_),
    .S(_01254_),
    .X(_01693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15646_ (.A0(_01690_),
    .A1(_01691_),
    .S(_01246_),
    .X(_01692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15647_ (.A0(_01552_),
    .A1(_01555_),
    .S(_01254_),
    .X(_01691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15648_ (.A0(_01549_),
    .A1(_01551_),
    .S(_01254_),
    .X(_01690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15649_ (.A0(_01532_),
    .A1(_01535_),
    .S(_01254_),
    .X(_01683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15650_ (.A0(_01683_),
    .A1(_01684_),
    .S(_01246_),
    .X(_01685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15651_ (.A0(_01685_),
    .A1(_01688_),
    .S(_01238_),
    .X(_01689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15652_ (.A0(_01686_),
    .A1(_01687_),
    .S(_01246_),
    .X(_01688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15653_ (.A0(_01544_),
    .A1(_01548_),
    .S(_01254_),
    .X(_01687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15654_ (.A0(_01541_),
    .A1(_01543_),
    .S(_01254_),
    .X(_01686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15655_ (.A0(_01536_),
    .A1(_01539_),
    .S(_01254_),
    .X(_01684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15656_ (.A0(_01678_),
    .A1(_01526_),
    .S(_01254_),
    .X(_01679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15657_ (.A0(_00793_),
    .A1(_01248_),
    .S(_01261_),
    .X(_01678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15658_ (.A0(_01648_),
    .A1(_01255_),
    .S(_01263_),
    .X(_01649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15659_ (.A0(_01649_),
    .A1(_01605_),
    .S(_01287_),
    .X(_01650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15660_ (.A0(_01653_),
    .A1(_01665_),
    .S(_01378_),
    .X(_01666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15661_ (.A0(_01666_),
    .A1(_01656_),
    .S(_01423_),
    .X(_01667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15662_ (.A0(_01667_),
    .A1(_01662_),
    .S(_01372_),
    .X(_01668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15663_ (.A0(_01656_),
    .A1(_01653_),
    .S(_01364_),
    .X(_01657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15664_ (.A0(_01657_),
    .A1(_01653_),
    .S(_01363_),
    .X(_01658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15665_ (.A0(_01669_),
    .A1(_00801_),
    .S(_01593_),
    .X(_01670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15666_ (.A0(_01670_),
    .A1(_01603_),
    .S(_00822_),
    .X(_01671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15667_ (.A0(_01671_),
    .A1(_01672_),
    .S(_01596_),
    .X(_01673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15668_ (.A0(_01663_),
    .A1(_01664_),
    .S(\design_top.XADDR[31] ),
    .X(_01665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15669_ (.A0(_01582_),
    .A1(_01660_),
    .S(\design_top.XADDR[3] ),
    .X(_01661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15670_ (.A0(_01659_),
    .A1(_01661_),
    .S(\design_top.XADDR[31] ),
    .X(_01662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15671_ (.A0(_01654_),
    .A1(_01655_),
    .S(\design_top.XADDR[31] ),
    .X(_01656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15672_ (.A0(_01651_),
    .A1(_01652_),
    .S(\design_top.XADDR[31] ),
    .X(_01653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15673_ (.A0(_01634_),
    .A1(_01644_),
    .S(_01238_),
    .X(_01645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15674_ (.A0(_01637_),
    .A1(_01643_),
    .S(_01246_),
    .X(_01644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15675_ (.A0(_01638_),
    .A1(_00843_),
    .S(_01254_),
    .X(_01643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15676_ (.A0(_01634_),
    .A1(_01641_),
    .S(_01238_),
    .X(_01642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15677_ (.A0(_01637_),
    .A1(_01640_),
    .S(_01246_),
    .X(_01641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15678_ (.A0(_01638_),
    .A1(_01639_),
    .S(_01254_),
    .X(_01640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15679_ (.A0(_00871_),
    .A1(_00857_),
    .S(_01261_),
    .X(_01638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15680_ (.A0(_01635_),
    .A1(_01636_),
    .S(_01254_),
    .X(_01637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15681_ (.A0(_00898_),
    .A1(_00885_),
    .S(_01261_),
    .X(_01636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15682_ (.A0(_00925_),
    .A1(_00912_),
    .S(_01261_),
    .X(_01635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15683_ (.A0(_01630_),
    .A1(_01633_),
    .S(_01246_),
    .X(_01634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15684_ (.A0(_01631_),
    .A1(_01632_),
    .S(_01254_),
    .X(_01633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15685_ (.A0(_00952_),
    .A1(_00939_),
    .S(_01261_),
    .X(_01632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15686_ (.A0(_00979_),
    .A1(_00966_),
    .S(_01261_),
    .X(_01631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15687_ (.A0(_01628_),
    .A1(_01629_),
    .S(_01254_),
    .X(_01630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15688_ (.A0(_01006_),
    .A1(_00993_),
    .S(_01261_),
    .X(_01629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15689_ (.A0(_01048_),
    .A1(_01020_),
    .S(_01261_),
    .X(_01628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15690_ (.A0(_01248_),
    .A1(_00793_),
    .S(_01261_),
    .X(_01613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15691_ (.A0(_01613_),
    .A1(_01614_),
    .S(_01254_),
    .X(_01615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15692_ (.A0(_01615_),
    .A1(_01618_),
    .S(_01246_),
    .X(_01619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15693_ (.A0(_01619_),
    .A1(_01626_),
    .S(_01238_),
    .X(_01627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15694_ (.A0(_01622_),
    .A1(_01625_),
    .S(_01246_),
    .X(_01626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15695_ (.A0(_01623_),
    .A1(_01624_),
    .S(_01254_),
    .X(_01625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15696_ (.A0(_01075_),
    .A1(_01062_),
    .S(_01261_),
    .X(_01624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15697_ (.A0(_01102_),
    .A1(_01089_),
    .S(_01261_),
    .X(_01623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15698_ (.A0(_01620_),
    .A1(_01621_),
    .S(_01254_),
    .X(_01622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15699_ (.A0(_01540_),
    .A1(_01116_),
    .S(_01261_),
    .X(_01621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15700_ (.A0(_01156_),
    .A1(_01142_),
    .S(_01261_),
    .X(_01620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15701_ (.A0(_01616_),
    .A1(_01617_),
    .S(_01254_),
    .X(_01618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15702_ (.A0(_01184_),
    .A1(_01171_),
    .S(_01261_),
    .X(_01617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15703_ (.A0(_01534_),
    .A1(_01198_),
    .S(_01261_),
    .X(_01616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15704_ (.A0(_01232_),
    .A1(_01224_),
    .S(_01261_),
    .X(_01614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15705_ (.A0(_01248_),
    .A1(_01290_),
    .S(_01261_),
    .X(_01608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15706_ (.A0(\design_top.core0.XIDATA[10] ),
    .A1(\design_top.core0.RESMODE[3] ),
    .S(\design_top.core0.XRES ),
    .X(_01602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15707_ (.A0(\design_top.core0.XIDATA[9] ),
    .A1(\design_top.core0.RESMODE[2] ),
    .S(\design_top.core0.XRES ),
    .X(_01601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15708_ (.A0(\design_top.core0.XIDATA[8] ),
    .A1(\design_top.core0.RESMODE[1] ),
    .S(\design_top.core0.XRES ),
    .X(_01600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15709_ (.A0(\design_top.core0.XIDATA[7] ),
    .A1(\design_top.core0.RESMODE[0] ),
    .S(\design_top.core0.XRES ),
    .X(_01599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15710_ (.A0(_01564_),
    .A1(_01530_),
    .S(_01362_),
    .X(_01565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15711_ (.A0(_01565_),
    .A1(_01291_),
    .S(_01323_),
    .X(_01566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15712_ (.A0(_01566_),
    .A1(_01262_),
    .S(_01524_),
    .X(_01567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15713_ (.A0(_01567_),
    .A1(_01286_),
    .S(_01523_),
    .X(_01568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15714_ (.A0(_01568_),
    .A1(_01291_),
    .S(_01263_),
    .X(_01569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15715_ (.A0(_01569_),
    .A1(_01522_),
    .S(_01287_),
    .X(_01570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15716_ (.A0(_01575_),
    .A1(_01588_),
    .S(_01378_),
    .X(_01589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15717_ (.A0(_01589_),
    .A1(_01578_),
    .S(_01423_),
    .X(_01590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15718_ (.A0(_01590_),
    .A1(_01585_),
    .S(_01372_),
    .X(_01591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15719_ (.A0(_01578_),
    .A1(_01575_),
    .S(_01364_),
    .X(_01579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15720_ (.A0(_01579_),
    .A1(_01575_),
    .S(_01363_),
    .X(_01580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15721_ (.A0(_01592_),
    .A1(_00802_),
    .S(_01593_),
    .X(_01594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15722_ (.A0(_01594_),
    .A1(_01520_),
    .S(_00822_),
    .X(_01595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15723_ (.A0(_01595_),
    .A1(_01597_),
    .S(_01596_),
    .X(_01598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15724_ (.A0(_01586_),
    .A1(_01587_),
    .S(\design_top.XADDR[31] ),
    .X(_01588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15725_ (.A0(_01582_),
    .A1(_01583_),
    .S(\design_top.XADDR[3] ),
    .X(_01584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15726_ (.A0(_01581_),
    .A1(_01584_),
    .S(\design_top.XADDR[31] ),
    .X(_01585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15727_ (.A0(_01576_),
    .A1(_01577_),
    .S(\design_top.XADDR[31] ),
    .X(_01578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15728_ (.A0(_01571_),
    .A1(_01574_),
    .S(\design_top.XADDR[31] ),
    .X(_01575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15729_ (.A0(_01290_),
    .A1(_01248_),
    .S(_01261_),
    .X(_01531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15730_ (.A0(_01531_),
    .A1(_01532_),
    .S(_01254_),
    .X(_01533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15731_ (.A0(_01533_),
    .A1(_01537_),
    .S(_01246_),
    .X(_01538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15732_ (.A0(_01538_),
    .A1(_01546_),
    .S(_01238_),
    .X(_01547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15733_ (.A0(_01547_),
    .A1(_01562_),
    .S(_01230_),
    .X(_01563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15734_ (.A0(_01554_),
    .A1(_01561_),
    .S(_01238_),
    .X(_01562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15735_ (.A0(_01557_),
    .A1(_01560_),
    .S(_01246_),
    .X(_01561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15736_ (.A0(_01558_),
    .A1(_01559_),
    .S(_01254_),
    .X(_01560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15737_ (.A0(_00857_),
    .A1(_00843_),
    .S(_01261_),
    .X(_01559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15738_ (.A0(_00885_),
    .A1(_00871_),
    .S(_01261_),
    .X(_01558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15739_ (.A0(_01555_),
    .A1(_01556_),
    .S(_01254_),
    .X(_01557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15740_ (.A0(_00912_),
    .A1(_00898_),
    .S(_01261_),
    .X(_01556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15741_ (.A0(_00939_),
    .A1(_00925_),
    .S(_01261_),
    .X(_01555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15742_ (.A0(_01550_),
    .A1(_01553_),
    .S(_01246_),
    .X(_01554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15743_ (.A0(_01551_),
    .A1(_01552_),
    .S(_01254_),
    .X(_01553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15744_ (.A0(_00966_),
    .A1(_00952_),
    .S(_01261_),
    .X(_01552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15745_ (.A0(_00993_),
    .A1(_00979_),
    .S(_01261_),
    .X(_01551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15746_ (.A0(_01548_),
    .A1(_01549_),
    .S(_01254_),
    .X(_01550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15747_ (.A0(_01020_),
    .A1(_01006_),
    .S(_01261_),
    .X(_01549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15748_ (.A0(_01062_),
    .A1(_01048_),
    .S(_01261_),
    .X(_01548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15749_ (.A0(_01542_),
    .A1(_01545_),
    .S(_01246_),
    .X(_01546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15750_ (.A0(_01543_),
    .A1(_01544_),
    .S(_01254_),
    .X(_01545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15751_ (.A0(_01089_),
    .A1(_01075_),
    .S(_01261_),
    .X(_01544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15752_ (.A0(_01116_),
    .A1(_01102_),
    .S(_01261_),
    .X(_01543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15753_ (.A0(_01539_),
    .A1(_01541_),
    .S(_01254_),
    .X(_01542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15754_ (.A0(_01142_),
    .A1(_01540_),
    .S(_01261_),
    .X(_01541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15755_ (.A0(_01171_),
    .A1(_01156_),
    .S(_01261_),
    .X(_01539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15756_ (.A0(_01535_),
    .A1(_01536_),
    .S(_01254_),
    .X(_01537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15757_ (.A0(_01198_),
    .A1(_01184_),
    .S(_01261_),
    .X(_01536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15758_ (.A0(_01224_),
    .A1(_01534_),
    .S(_01261_),
    .X(_01535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15759_ (.A0(_00793_),
    .A1(_01232_),
    .S(_01261_),
    .X(_01532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15760_ (.A0(\design_top.ROMFF[6] ),
    .A1(\design_top.ROMFF2[6] ),
    .S(\design_top.HLT2 ),
    .X(_01422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15761_ (.A0(\design_top.ROMFF[5] ),
    .A1(\design_top.ROMFF2[5] ),
    .S(\design_top.HLT2 ),
    .X(_01421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15762_ (.A0(\design_top.ROMFF[4] ),
    .A1(\design_top.ROMFF2[4] ),
    .S(\design_top.HLT2 ),
    .X(_01420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15763_ (.A0(_01381_),
    .A1(_01377_),
    .S(_01366_),
    .X(_01382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15764_ (.A0(_01379_),
    .A1(_01377_),
    .S(_01366_),
    .X(_01380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15765_ (.A0(_01373_),
    .A1(_01365_),
    .S(_01366_),
    .X(_01374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15766_ (.A0(_01368_),
    .A1(_01365_),
    .S(_01366_),
    .X(_01369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15767_ (.A0(_01291_),
    .A1(_01322_),
    .S(_01323_),
    .X(_01324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15768_ (.A0(_01324_),
    .A1(_01288_),
    .S(_01289_),
    .X(_01325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15769_ (.A0(_01325_),
    .A1(_01286_),
    .S(_01287_),
    .X(_01326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15770_ (.A0(_01326_),
    .A1(_01264_),
    .S(_01265_),
    .X(_01327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15771_ (.A0(_01327_),
    .A1(_01262_),
    .S(_01263_),
    .X(_01328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15772_ (.A0(_01121_),
    .A1(\design_top.core0.UIMM[12] ),
    .S(\design_top.core0.XMCC ),
    .X(_01285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15773_ (.A0(_01107_),
    .A1(\design_top.core0.UIMM[13] ),
    .S(\design_top.core0.XMCC ),
    .X(_01284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15774_ (.A0(_01094_),
    .A1(\design_top.core0.UIMM[14] ),
    .S(\design_top.core0.XMCC ),
    .X(_01283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15775_ (.A0(_01080_),
    .A1(\design_top.core0.UIMM[15] ),
    .S(\design_top.core0.XMCC ),
    .X(_01282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15776_ (.A0(_01067_),
    .A1(\design_top.core0.UIMM[16] ),
    .S(\design_top.core0.XMCC ),
    .X(_01281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15777_ (.A0(_01053_),
    .A1(\design_top.core0.UIMM[17] ),
    .S(\design_top.core0.XMCC ),
    .X(_01280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15778_ (.A0(_01025_),
    .A1(\design_top.core0.UIMM[18] ),
    .S(\design_top.core0.XMCC ),
    .X(_01279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15779_ (.A0(_01011_),
    .A1(\design_top.core0.UIMM[19] ),
    .S(\design_top.core0.XMCC ),
    .X(_01278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15780_ (.A0(_00998_),
    .A1(\design_top.core0.UIMM[20] ),
    .S(\design_top.core0.XMCC ),
    .X(_01277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15781_ (.A0(_00984_),
    .A1(\design_top.core0.UIMM[21] ),
    .S(\design_top.core0.XMCC ),
    .X(_01276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15782_ (.A0(_00971_),
    .A1(\design_top.core0.UIMM[22] ),
    .S(\design_top.core0.XMCC ),
    .X(_01275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15783_ (.A0(_00957_),
    .A1(\design_top.core0.UIMM[23] ),
    .S(\design_top.core0.XMCC ),
    .X(_01274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15784_ (.A0(_00944_),
    .A1(\design_top.core0.UIMM[24] ),
    .S(\design_top.core0.XMCC ),
    .X(_01273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15785_ (.A0(_00930_),
    .A1(\design_top.core0.UIMM[25] ),
    .S(\design_top.core0.XMCC ),
    .X(_01272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15786_ (.A0(_00917_),
    .A1(\design_top.core0.UIMM[26] ),
    .S(\design_top.core0.XMCC ),
    .X(_01271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15787_ (.A0(_00903_),
    .A1(\design_top.core0.UIMM[27] ),
    .S(\design_top.core0.XMCC ),
    .X(_01270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15788_ (.A0(_00890_),
    .A1(\design_top.core0.UIMM[28] ),
    .S(\design_top.core0.XMCC ),
    .X(_01269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15789_ (.A0(_00876_),
    .A1(\design_top.core0.UIMM[29] ),
    .S(\design_top.core0.XMCC ),
    .X(_01268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15790_ (.A0(_00862_),
    .A1(\design_top.core0.UIMM[30] ),
    .S(\design_top.core0.XMCC ),
    .X(_01267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15791_ (.A0(_00848_),
    .A1(\design_top.core0.UIMM[31] ),
    .S(\design_top.core0.XMCC ),
    .X(_01266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15792_ (.A0(_01260_),
    .A1(\design_top.core0.SIMM[0] ),
    .S(\design_top.core0.XMCC ),
    .X(_01261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15793_ (.A0(_01253_),
    .A1(\design_top.core0.SIMM[1] ),
    .S(\design_top.core0.XMCC ),
    .X(_01254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15794_ (.A0(_01245_),
    .A1(\design_top.core0.SIMM[2] ),
    .S(\design_top.core0.XMCC ),
    .X(_01246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15795_ (.A0(_01237_),
    .A1(\design_top.core0.SIMM[3] ),
    .S(\design_top.core0.XMCC ),
    .X(_01238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15796_ (.A0(_01229_),
    .A1(\design_top.core0.SIMM[4] ),
    .S(\design_top.core0.XMCC ),
    .X(_01230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15797_ (.A0(_01215_),
    .A1(\design_top.core0.SIMM[5] ),
    .S(\design_top.core0.XMCC ),
    .X(_01216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15798_ (.A0(_01203_),
    .A1(\design_top.core0.SIMM[6] ),
    .S(\design_top.core0.XMCC ),
    .X(_01204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15799_ (.A0(_01189_),
    .A1(\design_top.core0.SIMM[7] ),
    .S(\design_top.core0.XMCC ),
    .X(_01190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15800_ (.A0(_01176_),
    .A1(\design_top.core0.SIMM[8] ),
    .S(\design_top.core0.XMCC ),
    .X(_01177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15801_ (.A0(_01152_),
    .A1(_01155_),
    .S(_00432_),
    .X(_01164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15802_ (.A0(_01161_),
    .A1(\design_top.core0.SIMM[9] ),
    .S(\design_top.core0.XMCC ),
    .X(_01162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15803_ (.A0(_01153_),
    .A1(_01154_),
    .S(_00431_),
    .X(_01155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15804_ (.A0(_01150_),
    .A1(_01151_),
    .S(_00431_),
    .X(_01152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15805_ (.A0(_01147_),
    .A1(\design_top.core0.SIMM[10] ),
    .S(\design_top.core0.XMCC ),
    .X(_01148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15806_ (.A0(_01133_),
    .A1(\design_top.core0.SIMM[11] ),
    .S(\design_top.core0.XMCC ),
    .X(_01134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15807_ (.A0(_01121_),
    .A1(\design_top.core0.SIMM[12] ),
    .S(\design_top.core0.XMCC ),
    .X(_01122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15808_ (.A0(_01107_),
    .A1(\design_top.core0.SIMM[13] ),
    .S(\design_top.core0.XMCC ),
    .X(_01108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15809_ (.A0(_01094_),
    .A1(\design_top.core0.SIMM[14] ),
    .S(\design_top.core0.XMCC ),
    .X(_01095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15810_ (.A0(_01080_),
    .A1(\design_top.core0.SIMM[15] ),
    .S(\design_top.core0.XMCC ),
    .X(_01081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15811_ (.A0(_01067_),
    .A1(\design_top.core0.SIMM[16] ),
    .S(\design_top.core0.XMCC ),
    .X(_01068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15812_ (.A0(_01053_),
    .A1(\design_top.core0.SIMM[17] ),
    .S(\design_top.core0.XMCC ),
    .X(_01054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15813_ (.A0(_01025_),
    .A1(\design_top.core0.SIMM[18] ),
    .S(\design_top.core0.XMCC ),
    .X(_01026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15814_ (.A0(_01011_),
    .A1(\design_top.core0.SIMM[19] ),
    .S(\design_top.core0.XMCC ),
    .X(_01012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15815_ (.A0(_00998_),
    .A1(\design_top.core0.SIMM[20] ),
    .S(\design_top.core0.XMCC ),
    .X(_00999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15816_ (.A0(_00984_),
    .A1(\design_top.core0.SIMM[21] ),
    .S(\design_top.core0.XMCC ),
    .X(_00985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15817_ (.A0(_00971_),
    .A1(\design_top.core0.SIMM[22] ),
    .S(\design_top.core0.XMCC ),
    .X(_00972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15818_ (.A0(_00957_),
    .A1(\design_top.core0.SIMM[23] ),
    .S(\design_top.core0.XMCC ),
    .X(_00958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15819_ (.A0(_00944_),
    .A1(\design_top.core0.SIMM[24] ),
    .S(\design_top.core0.XMCC ),
    .X(_00945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15820_ (.A0(_00930_),
    .A1(\design_top.core0.SIMM[25] ),
    .S(\design_top.core0.XMCC ),
    .X(_00931_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15821_ (.A0(_00917_),
    .A1(\design_top.core0.SIMM[26] ),
    .S(\design_top.core0.XMCC ),
    .X(_00918_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15822_ (.A0(_00903_),
    .A1(\design_top.core0.SIMM[27] ),
    .S(\design_top.core0.XMCC ),
    .X(_00904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15823_ (.A0(_00890_),
    .A1(\design_top.core0.SIMM[28] ),
    .S(\design_top.core0.XMCC ),
    .X(_00891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15824_ (.A0(_00876_),
    .A1(\design_top.core0.SIMM[29] ),
    .S(\design_top.core0.XMCC ),
    .X(_00877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15825_ (.A0(_00862_),
    .A1(\design_top.core0.SIMM[30] ),
    .S(\design_top.core0.XMCC ),
    .X(_00863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15826_ (.A0(_00848_),
    .A1(\design_top.core0.SIMM[31] ),
    .S(\design_top.core0.XMCC ),
    .X(_00849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15827_ (.A0(_00814_),
    .A1(_00817_),
    .S(_00432_),
    .X(_00818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15828_ (.A0(_00815_),
    .A1(_00816_),
    .S(_00431_),
    .X(_00817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15829_ (.A0(_00812_),
    .A1(_00813_),
    .S(_00431_),
    .X(_00814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15830_ (.A0(_00805_),
    .A1(_00808_),
    .S(_00432_),
    .X(_00809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15831_ (.A0(_00806_),
    .A1(_00807_),
    .S(_00431_),
    .X(_00808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15832_ (.A0(_00803_),
    .A1(_00804_),
    .S(_00431_),
    .X(_00805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15833_ (.A0(_00796_),
    .A1(_00799_),
    .S(_00432_),
    .X(_00800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15834_ (.A0(_00797_),
    .A1(_00798_),
    .S(_00431_),
    .X(_00799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15835_ (.A0(_00794_),
    .A1(_00795_),
    .S(_00431_),
    .X(_00796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15836_ (.A0(_00790_),
    .A1(_00791_),
    .S(_00431_),
    .X(_00792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15837_ (.A0(_00787_),
    .A1(_00788_),
    .S(_00431_),
    .X(_00789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15838_ (.A0(\design_top.IDATA[15] ),
    .A1(\design_top.core0.S1PTR[0] ),
    .S(\design_top.HLT ),
    .X(_00000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15839_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_01396_),
    .X(_00412_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15840_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_01396_),
    .X(_00411_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15841_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_01396_),
    .X(_00410_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15842_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_01396_),
    .X(_00409_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15843_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_01396_),
    .X(_00408_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15844_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_01396_),
    .X(_00407_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15845_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_01396_),
    .X(_00406_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15846_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_01396_),
    .X(_00405_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15847_ (.A0(_00740_),
    .A1(\design_top.IDATA[20] ),
    .S(_00008_),
    .X(_00741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15848_ (.A0(_00741_),
    .A1(\design_top.IDATA[7] ),
    .S(_00009_),
    .X(_00742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15849_ (.A0(_00742_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15850_ (.A0(_00737_),
    .A1(\design_top.IDATA[30] ),
    .S(_00008_),
    .X(_00738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15851_ (.A0(_00738_),
    .A1(\design_top.IDATA[30] ),
    .S(_00009_),
    .X(_00739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15852_ (.A0(_00739_),
    .A1(\design_top.IDATA[30] ),
    .S(_00010_),
    .X(_00048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15853_ (.A0(_00734_),
    .A1(_00701_),
    .S(_00008_),
    .X(_00735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15854_ (.A0(_00735_),
    .A1(_00701_),
    .S(_00009_),
    .X(_00736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15855_ (.A0(_00736_),
    .A1(_00701_),
    .S(_00010_),
    .X(_00077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15856_ (.A0(_00731_),
    .A1(_00697_),
    .S(_00008_),
    .X(_00732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15857_ (.A0(_00732_),
    .A1(_00697_),
    .S(_00009_),
    .X(_00733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15858_ (.A0(_00733_),
    .A1(_00697_),
    .S(_00010_),
    .X(_00076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15859_ (.A0(_00728_),
    .A1(_00693_),
    .S(_00008_),
    .X(_00729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15860_ (.A0(_00729_),
    .A1(_00693_),
    .S(_00009_),
    .X(_00730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15861_ (.A0(_00730_),
    .A1(_00693_),
    .S(_00010_),
    .X(_00075_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15862_ (.A0(_00725_),
    .A1(_00689_),
    .S(_00008_),
    .X(_00726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15863_ (.A0(_00726_),
    .A1(_00689_),
    .S(_00009_),
    .X(_00727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15864_ (.A0(_00727_),
    .A1(_00689_),
    .S(_00010_),
    .X(_00074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15865_ (.A0(_00722_),
    .A1(_00685_),
    .S(_00008_),
    .X(_00723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15866_ (.A0(_00723_),
    .A1(_00685_),
    .S(_00009_),
    .X(_00724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15867_ (.A0(_00724_),
    .A1(_00685_),
    .S(_00010_),
    .X(_00073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15868_ (.A0(_00719_),
    .A1(_00681_),
    .S(_00008_),
    .X(_00720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15869_ (.A0(_00720_),
    .A1(_00718_),
    .S(_00009_),
    .X(_00721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15870_ (.A0(_00721_),
    .A1(_00718_),
    .S(_00010_),
    .X(_00072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15871_ (.A0(_00715_),
    .A1(\design_top.IDATA[23] ),
    .S(_00008_),
    .X(_00716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15872_ (.A0(_00716_),
    .A1(\design_top.IDATA[10] ),
    .S(_00009_),
    .X(_00717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15873_ (.A0(_00717_),
    .A1(\design_top.IDATA[10] ),
    .S(_00010_),
    .X(_00071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15874_ (.A0(_00712_),
    .A1(\design_top.IDATA[22] ),
    .S(_00008_),
    .X(_00713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15875_ (.A0(_00713_),
    .A1(\design_top.IDATA[9] ),
    .S(_00009_),
    .X(_00714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15876_ (.A0(_00714_),
    .A1(\design_top.IDATA[9] ),
    .S(_00010_),
    .X(_00069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15877_ (.A0(_00709_),
    .A1(\design_top.IDATA[21] ),
    .S(_00008_),
    .X(_00710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15878_ (.A0(_00710_),
    .A1(\design_top.IDATA[8] ),
    .S(_00009_),
    .X(_00711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15879_ (.A0(_00711_),
    .A1(\design_top.IDATA[8] ),
    .S(_00010_),
    .X(_00058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15880_ (.A0(_00708_),
    .A1(\design_top.IDATA[7] ),
    .S(_00010_),
    .X(_00047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15881_ (.A0(\design_top.IDATA[16] ),
    .A1(\design_top.core0.S1PTR[1] ),
    .S(\design_top.HLT ),
    .X(_00001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15882_ (.A0(\design_top.IDATA[30] ),
    .A1(\design_top.IDATA[31] ),
    .S(_00643_),
    .X(_00705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15883_ (.A0(_00705_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_00706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15884_ (.A0(_00706_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15885_ (.A0(_00707_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15886_ (.A0(_00701_),
    .A1(\design_top.IDATA[31] ),
    .S(_00643_),
    .X(_00702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15887_ (.A0(_00702_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_00703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15888_ (.A0(_00703_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15889_ (.A0(_00704_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00068_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15890_ (.A0(_00697_),
    .A1(\design_top.IDATA[31] ),
    .S(_00643_),
    .X(_00698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15891_ (.A0(_00698_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_00699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15892_ (.A0(_00699_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15893_ (.A0(_00700_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15894_ (.A0(_00693_),
    .A1(\design_top.IDATA[31] ),
    .S(_00643_),
    .X(_00694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15895_ (.A0(_00694_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_00695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15896_ (.A0(_00695_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15897_ (.A0(_00696_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15898_ (.A0(_00689_),
    .A1(\design_top.IDATA[31] ),
    .S(_00643_),
    .X(_00690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15899_ (.A0(_00690_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_00691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15900_ (.A0(_00691_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15901_ (.A0(_00692_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15902_ (.A0(_00685_),
    .A1(\design_top.IDATA[31] ),
    .S(_00643_),
    .X(_00686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15903_ (.A0(_00686_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_00687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15904_ (.A0(_00687_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15905_ (.A0(_00688_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15906_ (.A0(_00681_),
    .A1(\design_top.IDATA[31] ),
    .S(_00643_),
    .X(_00682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15907_ (.A0(_00682_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_00683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15908_ (.A0(_00683_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15909_ (.A0(_00684_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15910_ (.A0(\design_top.IDATA[23] ),
    .A1(\design_top.IDATA[31] ),
    .S(_00643_),
    .X(_00678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15911_ (.A0(_00678_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_00679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15912_ (.A0(_00679_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15913_ (.A0(_00680_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15914_ (.A0(\design_top.IDATA[22] ),
    .A1(\design_top.IDATA[31] ),
    .S(_00643_),
    .X(_00675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15915_ (.A0(_00675_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_00676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15916_ (.A0(_00676_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15917_ (.A0(_00677_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15918_ (.A0(\design_top.IDATA[21] ),
    .A1(\design_top.IDATA[31] ),
    .S(_00643_),
    .X(_00672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15919_ (.A0(_00672_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_00673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15920_ (.A0(_00673_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15921_ (.A0(_00674_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15922_ (.A0(\design_top.IDATA[20] ),
    .A1(\design_top.IDATA[31] ),
    .S(_00643_),
    .X(_00669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15923_ (.A0(_00669_),
    .A1(\design_top.IDATA[31] ),
    .S(_00008_),
    .X(_00670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15924_ (.A0(_00670_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15925_ (.A0(_00671_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15926_ (.A0(_00665_),
    .A1(\design_top.IDATA[31] ),
    .S(_00643_),
    .X(_00666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15927_ (.A0(_00666_),
    .A1(_00665_),
    .S(_00008_),
    .X(_00667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15928_ (.A0(_00667_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15929_ (.A0(_00668_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15930_ (.A0(\design_top.IDATA[18] ),
    .A1(\design_top.IDATA[31] ),
    .S(_00643_),
    .X(_00662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15931_ (.A0(_00662_),
    .A1(\design_top.IDATA[18] ),
    .S(_00008_),
    .X(_00663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15932_ (.A0(_00663_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15933_ (.A0(_00664_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15934_ (.A0(\design_top.IDATA[17] ),
    .A1(\design_top.IDATA[31] ),
    .S(_00643_),
    .X(_00659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15935_ (.A0(_00659_),
    .A1(\design_top.IDATA[17] ),
    .S(_00008_),
    .X(_00660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15936_ (.A0(_00660_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15937_ (.A0(_00661_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15938_ (.A0(\design_top.IDATA[16] ),
    .A1(\design_top.IDATA[31] ),
    .S(_00643_),
    .X(_00656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15939_ (.A0(_00656_),
    .A1(\design_top.IDATA[16] ),
    .S(_00008_),
    .X(_00657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15940_ (.A0(_00657_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15941_ (.A0(_00658_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15942_ (.A0(\design_top.IDATA[15] ),
    .A1(\design_top.IDATA[31] ),
    .S(_00643_),
    .X(_00653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15943_ (.A0(_00653_),
    .A1(\design_top.IDATA[15] ),
    .S(_00008_),
    .X(_00654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15944_ (.A0(_00654_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15945_ (.A0(_00655_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15946_ (.A0(\design_top.IDATA[14] ),
    .A1(\design_top.IDATA[31] ),
    .S(_00643_),
    .X(_00650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15947_ (.A0(_00650_),
    .A1(\design_top.IDATA[14] ),
    .S(_00008_),
    .X(_00651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15948_ (.A0(_00651_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15949_ (.A0(_00652_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15950_ (.A0(\design_top.IDATA[13] ),
    .A1(\design_top.IDATA[31] ),
    .S(_00643_),
    .X(_00647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15951_ (.A0(_00647_),
    .A1(\design_top.IDATA[13] ),
    .S(_00008_),
    .X(_00648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15952_ (.A0(_00648_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15953_ (.A0(_00649_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15954_ (.A0(\design_top.IDATA[12] ),
    .A1(\design_top.IDATA[31] ),
    .S(_00643_),
    .X(_00644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15955_ (.A0(_00644_),
    .A1(\design_top.IDATA[12] ),
    .S(_00008_),
    .X(_00645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15956_ (.A0(_00645_),
    .A1(\design_top.IDATA[31] ),
    .S(_00009_),
    .X(_00646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15957_ (.A0(_00646_),
    .A1(\design_top.IDATA[31] ),
    .S(_00010_),
    .X(_00050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15958_ (.A0(\design_top.IDATA[22] ),
    .A1(\design_top.core0.S2PTR[2] ),
    .S(\design_top.HLT ),
    .X(_00006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15959_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_01416_),
    .X(_00180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15960_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_01416_),
    .X(_00179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15961_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_01416_),
    .X(_00178_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15962_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_01416_),
    .X(_00177_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15963_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_01416_),
    .X(_00176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15964_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_01416_),
    .X(_00175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15965_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_01416_),
    .X(_00174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15966_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_01416_),
    .X(_00173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15967_ (.A0(\design_top.IDATA[23] ),
    .A1(\design_top.core0.S2PTR[3] ),
    .S(\design_top.HLT ),
    .X(_00007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15968_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_01397_),
    .X(_00268_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15969_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_01397_),
    .X(_00267_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15970_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_01397_),
    .X(_00266_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15971_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_01397_),
    .X(_00265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15972_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_01397_),
    .X(_00264_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15973_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_01397_),
    .X(_00263_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15974_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_01397_),
    .X(_00262_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15975_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_01397_),
    .X(_00261_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15976_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_01383_),
    .X(_00356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15977_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_01383_),
    .X(_00355_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15978_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_01383_),
    .X(_00354_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15979_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_01383_),
    .X(_00353_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15980_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_01383_),
    .X(_00352_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15981_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_01383_),
    .X(_00351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15982_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_01383_),
    .X(_00350_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15983_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_01383_),
    .X(_00349_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15984_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_01408_),
    .X(_00380_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15985_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_01408_),
    .X(_00379_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15986_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_01408_),
    .X(_00378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15987_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_01408_),
    .X(_00377_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15988_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_01408_),
    .X(_00376_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15989_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_01408_),
    .X(_00375_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15990_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_01408_),
    .X(_00374_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15991_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_01408_),
    .X(_00373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15992_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_01407_),
    .X(_00388_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15993_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_01407_),
    .X(_00387_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15994_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_01407_),
    .X(_00386_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15995_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_01407_),
    .X(_00385_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15996_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_01407_),
    .X(_00384_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15997_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_01407_),
    .X(_00383_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15998_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_01407_),
    .X(_00382_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _15999_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_01407_),
    .X(_00381_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16000_ (.A0(_00637_),
    .A1(_00642_),
    .S(\design_top.IADDR[6] ),
    .X(_00165_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16001_ (.A0(_00627_),
    .A1(_00632_),
    .S(\design_top.IADDR[6] ),
    .X(_00164_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16002_ (.A0(_00617_),
    .A1(_00622_),
    .S(\design_top.IADDR[6] ),
    .X(_00162_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16003_ (.A0(_00607_),
    .A1(_00612_),
    .S(\design_top.IADDR[6] ),
    .X(_00161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16004_ (.A0(_00597_),
    .A1(_00602_),
    .S(\design_top.IADDR[6] ),
    .X(_00160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16005_ (.A0(_00587_),
    .A1(_00592_),
    .S(\design_top.IADDR[6] ),
    .X(_00159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16006_ (.A0(_00577_),
    .A1(_00582_),
    .S(\design_top.IADDR[6] ),
    .X(_00158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16007_ (.A0(_00567_),
    .A1(_00572_),
    .S(\design_top.IADDR[6] ),
    .X(_00157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16008_ (.A0(_00557_),
    .A1(_00562_),
    .S(\design_top.IADDR[6] ),
    .X(_00156_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16009_ (.A0(_00547_),
    .A1(_00552_),
    .S(\design_top.IADDR[6] ),
    .X(_00155_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16010_ (.A0(_00537_),
    .A1(_00542_),
    .S(\design_top.IADDR[6] ),
    .X(_00154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16011_ (.A0(_00527_),
    .A1(_00532_),
    .S(\design_top.IADDR[6] ),
    .X(_00153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16012_ (.A0(_00517_),
    .A1(_00522_),
    .S(\design_top.IADDR[6] ),
    .X(_00151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16013_ (.A0(_00507_),
    .A1(_00512_),
    .S(\design_top.IADDR[6] ),
    .X(_00150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16014_ (.A0(_00497_),
    .A1(_00502_),
    .S(\design_top.IADDR[6] ),
    .X(_00149_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16015_ (.A0(_00487_),
    .A1(_00492_),
    .S(\design_top.IADDR[6] ),
    .X(_00148_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16016_ (.A0(_00477_),
    .A1(_00482_),
    .S(\design_top.IADDR[6] ),
    .X(_00147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16017_ (.A0(_00467_),
    .A1(_00472_),
    .S(\design_top.IADDR[6] ),
    .X(_00146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16018_ (.A0(_00457_),
    .A1(_00462_),
    .S(\design_top.IADDR[6] ),
    .X(_00145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16019_ (.A0(_00447_),
    .A1(_00452_),
    .S(\design_top.IADDR[6] ),
    .X(_00144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16020_ (.A0(_00437_),
    .A1(_00442_),
    .S(\design_top.IADDR[6] ),
    .X(_00143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16021_ (.A0(_03049_),
    .A1(_03054_),
    .S(\design_top.IADDR[6] ),
    .X(_00142_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16022_ (.A0(_03039_),
    .A1(_03044_),
    .S(\design_top.IADDR[6] ),
    .X(_00172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16023_ (.A0(_03029_),
    .A1(_03034_),
    .S(\design_top.IADDR[6] ),
    .X(_00171_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16024_ (.A0(_03019_),
    .A1(_03024_),
    .S(\design_top.IADDR[6] ),
    .X(_00170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16025_ (.A0(_03009_),
    .A1(_03014_),
    .S(\design_top.IADDR[6] ),
    .X(_00169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16026_ (.A0(_02999_),
    .A1(_03004_),
    .S(\design_top.IADDR[6] ),
    .X(_00168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16027_ (.A0(_02989_),
    .A1(_02994_),
    .S(\design_top.IADDR[6] ),
    .X(_00167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16028_ (.A0(_02979_),
    .A1(_02984_),
    .S(\design_top.IADDR[6] ),
    .X(_00166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16029_ (.A0(_02969_),
    .A1(_02974_),
    .S(\design_top.IADDR[6] ),
    .X(_00163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16030_ (.A0(_02959_),
    .A1(_02964_),
    .S(\design_top.IADDR[6] ),
    .X(_00152_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16031_ (.A0(_02949_),
    .A1(_02954_),
    .S(\design_top.IADDR[6] ),
    .X(_00141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16032_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_01406_),
    .X(_00396_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16033_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_01406_),
    .X(_00395_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16034_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_01406_),
    .X(_00394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16035_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_01406_),
    .X(_00393_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16036_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_01406_),
    .X(_00392_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16037_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_01406_),
    .X(_00391_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16038_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_01406_),
    .X(_00390_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16039_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_01406_),
    .X(_00389_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16040_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_01405_),
    .X(_00404_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16041_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_01405_),
    .X(_00403_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16042_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_01405_),
    .X(_00402_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16043_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_01405_),
    .X(_00401_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16044_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_01405_),
    .X(_00400_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16045_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_01405_),
    .X(_00399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16046_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_01405_),
    .X(_00398_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16047_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_01405_),
    .X(_00397_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16048_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_01384_),
    .X(_00348_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16049_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_01384_),
    .X(_00347_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16050_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_01384_),
    .X(_00346_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16051_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_01384_),
    .X(_00345_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16052_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_01384_),
    .X(_00344_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16053_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_01384_),
    .X(_00343_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16054_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_01384_),
    .X(_00342_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16055_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_01384_),
    .X(_00341_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16056_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_01410_),
    .X(_00364_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16057_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_01410_),
    .X(_00363_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16058_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_01410_),
    .X(_00362_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16059_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_01410_),
    .X(_00361_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16060_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_01410_),
    .X(_00360_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16061_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_01410_),
    .X(_00359_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16062_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_01410_),
    .X(_00358_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16063_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_01410_),
    .X(_00357_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16064_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_01409_),
    .X(_00372_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16065_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_01409_),
    .X(_00371_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16066_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_01409_),
    .X(_00370_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16067_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_01409_),
    .X(_00369_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16068_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_01409_),
    .X(_00368_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16069_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_01409_),
    .X(_00367_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16070_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_01409_),
    .X(_00366_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16071_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_01409_),
    .X(_00365_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16072_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_01391_),
    .X(_00420_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16073_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_01391_),
    .X(_00419_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16074_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_01391_),
    .X(_00418_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16075_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_01391_),
    .X(_00417_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16076_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_01391_),
    .X(_00416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16077_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_01391_),
    .X(_00415_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16078_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_01391_),
    .X(_00414_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16079_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_01391_),
    .X(_00413_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16080_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_01390_),
    .X(_00428_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16081_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_01390_),
    .X(_00427_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16082_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_01390_),
    .X(_00426_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16083_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_01390_),
    .X(_00425_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16084_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_01390_),
    .X(_00424_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16085_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_01390_),
    .X(_00423_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16086_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_01390_),
    .X(_00422_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16087_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_01390_),
    .X(_00421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16088_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_01415_),
    .X(_00188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16089_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_01415_),
    .X(_00187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16090_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_01415_),
    .X(_00186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16091_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_01415_),
    .X(_00185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16092_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_01415_),
    .X(_00184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16093_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_01415_),
    .X(_00183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16094_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_01415_),
    .X(_00182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16095_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_01415_),
    .X(_00181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16096_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_01411_),
    .X(_00196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16097_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_01411_),
    .X(_00195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16098_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_01411_),
    .X(_00194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16099_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_01411_),
    .X(_00193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16100_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_01411_),
    .X(_00192_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16101_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_01411_),
    .X(_00191_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16102_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_01411_),
    .X(_00190_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16103_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_01411_),
    .X(_00189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16104_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_01418_),
    .X(_00204_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16105_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_01418_),
    .X(_00203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16106_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_01418_),
    .X(_00202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16107_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_01418_),
    .X(_00201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16108_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_01418_),
    .X(_00200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16109_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_01418_),
    .X(_00199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16110_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_01418_),
    .X(_00198_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16111_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_01418_),
    .X(_00197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16112_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_01404_),
    .X(_00212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16113_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_01404_),
    .X(_00211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16114_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_01404_),
    .X(_00210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16115_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_01404_),
    .X(_00209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16116_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_01404_),
    .X(_00208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16117_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_01404_),
    .X(_00207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16118_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_01404_),
    .X(_00206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16119_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_01404_),
    .X(_00205_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16120_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_01403_),
    .X(_00220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16121_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_01403_),
    .X(_00219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16122_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_01403_),
    .X(_00218_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16123_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_01403_),
    .X(_00217_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16124_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_01403_),
    .X(_00216_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16125_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_01403_),
    .X(_00215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16126_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_01403_),
    .X(_00214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16127_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_01403_),
    .X(_00213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16128_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_01402_),
    .X(_00228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16129_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_01402_),
    .X(_00227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16130_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_01402_),
    .X(_00226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16131_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_01402_),
    .X(_00225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16132_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_01402_),
    .X(_00224_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16133_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_01402_),
    .X(_00223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16134_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_01402_),
    .X(_00222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16135_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_01402_),
    .X(_00221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16136_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_01401_),
    .X(_00236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16137_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_01401_),
    .X(_00235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16138_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_01401_),
    .X(_00234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16139_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_01401_),
    .X(_00233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16140_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_01401_),
    .X(_00232_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16141_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_01401_),
    .X(_00231_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16142_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_01401_),
    .X(_00230_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16143_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_01401_),
    .X(_00229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16144_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_01400_),
    .X(_00244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16145_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_01400_),
    .X(_00243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16146_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_01400_),
    .X(_00242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16147_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_01400_),
    .X(_00241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16148_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_01400_),
    .X(_00240_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16149_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_01400_),
    .X(_00239_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16150_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_01400_),
    .X(_00238_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16151_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_01400_),
    .X(_00237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16152_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_01399_),
    .X(_00252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16153_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_01399_),
    .X(_00251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16154_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_01399_),
    .X(_00250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16155_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_01399_),
    .X(_00249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16156_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_01399_),
    .X(_00248_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16157_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_01399_),
    .X(_00247_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16158_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_01399_),
    .X(_00246_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16159_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_01399_),
    .X(_00245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16160_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_01395_),
    .X(_00276_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16161_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_01395_),
    .X(_00275_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16162_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_01395_),
    .X(_00274_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16163_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_01395_),
    .X(_00273_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16164_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_01395_),
    .X(_00272_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16165_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_01395_),
    .X(_00271_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16166_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_01395_),
    .X(_00270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16167_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_01395_),
    .X(_00269_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16168_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_01394_),
    .X(_00284_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16169_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_01394_),
    .X(_00283_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16170_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_01394_),
    .X(_00282_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16171_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_01394_),
    .X(_00281_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16172_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_01394_),
    .X(_00280_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16173_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_01394_),
    .X(_00279_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16174_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_01394_),
    .X(_00278_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16175_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_01394_),
    .X(_00277_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16176_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_01393_),
    .X(_00292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16177_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_01393_),
    .X(_00291_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16178_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_01393_),
    .X(_00290_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16179_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_01393_),
    .X(_00289_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16180_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_01393_),
    .X(_00288_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16181_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_01393_),
    .X(_00287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16182_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_01393_),
    .X(_00286_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16183_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_01393_),
    .X(_00285_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16184_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_01392_),
    .X(_00300_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16185_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_01392_),
    .X(_00299_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16186_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_01392_),
    .X(_00298_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16187_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_01392_),
    .X(_00297_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16188_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_01392_),
    .X(_00296_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16189_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_01392_),
    .X(_00295_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16190_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_01392_),
    .X(_00294_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16191_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_01392_),
    .X(_00293_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16192_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_01398_),
    .X(_00260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16193_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_01398_),
    .X(_00259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16194_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_01398_),
    .X(_00258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16195_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_01398_),
    .X(_00257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16196_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_01398_),
    .X(_00256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16197_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_01398_),
    .X(_00255_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16198_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_01398_),
    .X(_00254_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16199_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_01398_),
    .X(_00253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16200_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_01389_),
    .X(_00308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16201_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_01389_),
    .X(_00307_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16202_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_01389_),
    .X(_00306_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16203_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_01389_),
    .X(_00305_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16204_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_01389_),
    .X(_00304_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16205_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_01389_),
    .X(_00303_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16206_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_01389_),
    .X(_00302_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16207_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_01389_),
    .X(_00301_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16208_ (.A0(wbs_dat_i[15]),
    .A1(\design_top.DATAO[7] ),
    .S(_01388_),
    .X(_00316_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16209_ (.A0(wbs_dat_i[14]),
    .A1(\design_top.DATAO[6] ),
    .S(_01388_),
    .X(_00315_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16210_ (.A0(wbs_dat_i[13]),
    .A1(\design_top.DATAO[5] ),
    .S(_01388_),
    .X(_00314_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16211_ (.A0(wbs_dat_i[12]),
    .A1(\design_top.DATAO[4] ),
    .S(_01388_),
    .X(_00313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16212_ (.A0(wbs_dat_i[11]),
    .A1(\design_top.DATAO[3] ),
    .S(_01388_),
    .X(_00312_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16213_ (.A0(wbs_dat_i[10]),
    .A1(\design_top.DATAO[2] ),
    .S(_01388_),
    .X(_00311_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16214_ (.A0(wbs_dat_i[9]),
    .A1(\design_top.DATAO[1] ),
    .S(_01388_),
    .X(_00310_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16215_ (.A0(wbs_dat_i[8]),
    .A1(\design_top.DATAO[0] ),
    .S(_01388_),
    .X(_00309_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16216_ (.A0(wbs_dat_i[23]),
    .A1(\design_top.DATAO[7] ),
    .S(_01387_),
    .X(_00324_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16217_ (.A0(wbs_dat_i[22]),
    .A1(\design_top.DATAO[6] ),
    .S(_01387_),
    .X(_00323_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16218_ (.A0(wbs_dat_i[21]),
    .A1(\design_top.DATAO[5] ),
    .S(_01387_),
    .X(_00322_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16219_ (.A0(wbs_dat_i[20]),
    .A1(\design_top.DATAO[4] ),
    .S(_01387_),
    .X(_00321_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16220_ (.A0(wbs_dat_i[19]),
    .A1(\design_top.DATAO[3] ),
    .S(_01387_),
    .X(_00320_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16221_ (.A0(wbs_dat_i[18]),
    .A1(\design_top.DATAO[2] ),
    .S(_01387_),
    .X(_00319_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16222_ (.A0(wbs_dat_i[17]),
    .A1(\design_top.DATAO[1] ),
    .S(_01387_),
    .X(_00318_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16223_ (.A0(wbs_dat_i[16]),
    .A1(\design_top.DATAO[0] ),
    .S(_01387_),
    .X(_00317_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16224_ (.A0(wbs_dat_i[31]),
    .A1(\design_top.DATAO[7] ),
    .S(_01386_),
    .X(_00332_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16225_ (.A0(wbs_dat_i[30]),
    .A1(\design_top.DATAO[6] ),
    .S(_01386_),
    .X(_00331_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16226_ (.A0(wbs_dat_i[29]),
    .A1(\design_top.DATAO[5] ),
    .S(_01386_),
    .X(_00330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16227_ (.A0(wbs_dat_i[28]),
    .A1(\design_top.DATAO[4] ),
    .S(_01386_),
    .X(_00329_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16228_ (.A0(wbs_dat_i[27]),
    .A1(\design_top.DATAO[3] ),
    .S(_01386_),
    .X(_00328_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16229_ (.A0(wbs_dat_i[26]),
    .A1(\design_top.DATAO[2] ),
    .S(_01386_),
    .X(_00327_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16230_ (.A0(wbs_dat_i[25]),
    .A1(\design_top.DATAO[1] ),
    .S(_01386_),
    .X(_00326_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16231_ (.A0(wbs_dat_i[24]),
    .A1(\design_top.DATAO[0] ),
    .S(_01386_),
    .X(_00325_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16232_ (.A0(wbs_dat_i[7]),
    .A1(\design_top.DATAO[7] ),
    .S(_01385_),
    .X(_00340_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16233_ (.A0(wbs_dat_i[6]),
    .A1(\design_top.DATAO[6] ),
    .S(_01385_),
    .X(_00339_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16234_ (.A0(wbs_dat_i[5]),
    .A1(\design_top.DATAO[5] ),
    .S(_01385_),
    .X(_00338_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16235_ (.A0(wbs_dat_i[4]),
    .A1(\design_top.DATAO[4] ),
    .S(_01385_),
    .X(_00337_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16236_ (.A0(wbs_dat_i[3]),
    .A1(\design_top.DATAO[3] ),
    .S(_01385_),
    .X(_00336_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16237_ (.A0(wbs_dat_i[2]),
    .A1(\design_top.DATAO[2] ),
    .S(_01385_),
    .X(_00335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16238_ (.A0(wbs_dat_i[1]),
    .A1(\design_top.DATAO[1] ),
    .S(_01385_),
    .X(_00334_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16239_ (.A0(wbs_dat_i[0]),
    .A1(\design_top.DATAO[0] ),
    .S(_01385_),
    .X(_00333_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16240_ (.A0(_02944_),
    .A1(io_out[12]),
    .S(_01419_),
    .X(_00012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16241_ (.A0(\design_top.IDATA[18] ),
    .A1(\design_top.core0.S1PTR[3] ),
    .S(\design_top.HLT ),
    .X(_00003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16242_ (.A0(\design_top.IDATA[21] ),
    .A1(\design_top.core0.S2PTR[1] ),
    .S(\design_top.HLT ),
    .X(_00005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16243_ (.A0(_02943_),
    .A1(\design_top.IOMUX[3][31] ),
    .S(_01375_),
    .X(_00037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16244_ (.A0(_02942_),
    .A1(\design_top.IOMUX[3][30] ),
    .S(_01375_),
    .X(_00036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16245_ (.A0(_02941_),
    .A1(\design_top.IOMUX[3][29] ),
    .S(_01375_),
    .X(_00034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16246_ (.A0(_02940_),
    .A1(\design_top.IOMUX[3][28] ),
    .S(_01375_),
    .X(_00033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16247_ (.A0(_02939_),
    .A1(\design_top.IOMUX[3][27] ),
    .S(_01375_),
    .X(_00032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16248_ (.A0(_02938_),
    .A1(\design_top.IOMUX[3][26] ),
    .S(_01375_),
    .X(_00031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16249_ (.A0(_02937_),
    .A1(\design_top.IOMUX[3][25] ),
    .S(_01375_),
    .X(_00030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16250_ (.A0(_02936_),
    .A1(\design_top.IOMUX[3][24] ),
    .S(_01375_),
    .X(_00029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16251_ (.A0(_02935_),
    .A1(\design_top.IOMUX[3][23] ),
    .S(_01375_),
    .X(_00028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16252_ (.A0(_02934_),
    .A1(\design_top.IOMUX[3][22] ),
    .S(_01375_),
    .X(_00027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16253_ (.A0(_02933_),
    .A1(\design_top.IOMUX[3][21] ),
    .S(_01375_),
    .X(_00026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16254_ (.A0(_02932_),
    .A1(\design_top.IOMUX[3][20] ),
    .S(_01375_),
    .X(_00025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16255_ (.A0(_02931_),
    .A1(\design_top.IOMUX[3][19] ),
    .S(_01375_),
    .X(_00023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16256_ (.A0(_02930_),
    .A1(\design_top.IOMUX[3][18] ),
    .S(_01375_),
    .X(_00022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16257_ (.A0(_02929_),
    .A1(\design_top.IOMUX[3][17] ),
    .S(_01375_),
    .X(_00021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16258_ (.A0(_02928_),
    .A1(\design_top.IOMUX[3][16] ),
    .S(_01375_),
    .X(_00020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16259_ (.A0(_02927_),
    .A1(\design_top.IOMUX[3][15] ),
    .S(_01375_),
    .X(_00019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16260_ (.A0(_02926_),
    .A1(\design_top.IOMUX[3][14] ),
    .S(_01375_),
    .X(_00018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16261_ (.A0(_02925_),
    .A1(\design_top.IOMUX[3][13] ),
    .S(_01375_),
    .X(_00017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16262_ (.A0(_02924_),
    .A1(\design_top.IOMUX[3][12] ),
    .S(_01375_),
    .X(_00016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16263_ (.A0(_02923_),
    .A1(\design_top.IOMUX[3][11] ),
    .S(_01375_),
    .X(_00015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16264_ (.A0(_02922_),
    .A1(\design_top.IOMUX[3][10] ),
    .S(_01375_),
    .X(_00014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16265_ (.A0(_02921_),
    .A1(\design_top.IOMUX[3][9] ),
    .S(_01375_),
    .X(_00044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16266_ (.A0(_02920_),
    .A1(\design_top.IOMUX[3][8] ),
    .S(_01375_),
    .X(_00043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16267_ (.A0(_02919_),
    .A1(\design_top.IOMUX[3][7] ),
    .S(_01375_),
    .X(_00042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16268_ (.A0(_02918_),
    .A1(\design_top.IOMUX[3][6] ),
    .S(_01375_),
    .X(_00041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16269_ (.A0(_02917_),
    .A1(\design_top.IOMUX[3][5] ),
    .S(_01375_),
    .X(_00040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16270_ (.A0(_02916_),
    .A1(\design_top.IOMUX[3][4] ),
    .S(_01375_),
    .X(_00039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16271_ (.A0(_02915_),
    .A1(\design_top.IOMUX[3][3] ),
    .S(_01375_),
    .X(_00038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16272_ (.A0(_02914_),
    .A1(\design_top.IOMUX[3][2] ),
    .S(_01375_),
    .X(_00035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16273_ (.A0(_02913_),
    .A1(\design_top.IOMUX[3][1] ),
    .S(_01375_),
    .X(_00024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16274_ (.A0(_02912_),
    .A1(\design_top.IOMUX[3][0] ),
    .S(_01375_),
    .X(_00013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16275_ (.A0(\design_top.IDATA[17] ),
    .A1(\design_top.core0.S1PTR[2] ),
    .S(\design_top.HLT ),
    .X(_00002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16276_ (.A0(\design_top.IDATA[20] ),
    .A1(\design_top.core0.S2PTR[0] ),
    .S(\design_top.HLT ),
    .X(_00004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16277_ (.A0(_02911_),
    .A1(_02906_),
    .S(_01337_),
    .X(_00133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16278_ (.A0(_02901_),
    .A1(_02896_),
    .S(_01337_),
    .X(_00132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16279_ (.A0(_02891_),
    .A1(_02886_),
    .S(_01337_),
    .X(_00130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16280_ (.A0(_02881_),
    .A1(_02876_),
    .S(_01337_),
    .X(_00129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16281_ (.A0(_02871_),
    .A1(_02866_),
    .S(_01337_),
    .X(_00128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16282_ (.A0(_02861_),
    .A1(_02856_),
    .S(_01337_),
    .X(_00127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16283_ (.A0(_02851_),
    .A1(_02846_),
    .S(_01337_),
    .X(_00126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16284_ (.A0(_02841_),
    .A1(_02836_),
    .S(_01337_),
    .X(_00125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16285_ (.A0(_02831_),
    .A1(_02826_),
    .S(_01337_),
    .X(_00124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16286_ (.A0(_02821_),
    .A1(_02816_),
    .S(_01337_),
    .X(_00123_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16287_ (.A0(_02811_),
    .A1(_02806_),
    .S(_01337_),
    .X(_00122_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16288_ (.A0(_02801_),
    .A1(_02796_),
    .S(_01337_),
    .X(_00121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16289_ (.A0(_02791_),
    .A1(_02786_),
    .S(_01337_),
    .X(_00119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16290_ (.A0(_02781_),
    .A1(_02776_),
    .S(_01337_),
    .X(_00118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16291_ (.A0(_02771_),
    .A1(_02766_),
    .S(_01337_),
    .X(_00117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16292_ (.A0(_02761_),
    .A1(_02756_),
    .S(_01337_),
    .X(_00116_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16293_ (.A0(_02751_),
    .A1(_02746_),
    .S(_01337_),
    .X(_00115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16294_ (.A0(_02741_),
    .A1(_02736_),
    .S(_01337_),
    .X(_00114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16295_ (.A0(_02731_),
    .A1(_02726_),
    .S(_01337_),
    .X(_00113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16296_ (.A0(_02721_),
    .A1(_02716_),
    .S(_01337_),
    .X(_00112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16297_ (.A0(_02711_),
    .A1(_02706_),
    .S(_01337_),
    .X(_00111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16298_ (.A0(_02701_),
    .A1(_02696_),
    .S(_01337_),
    .X(_00110_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16299_ (.A0(_02691_),
    .A1(_02686_),
    .S(_01337_),
    .X(_00140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16300_ (.A0(_02681_),
    .A1(_02676_),
    .S(_01337_),
    .X(_00139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16301_ (.A0(_02671_),
    .A1(_02666_),
    .S(_01337_),
    .X(_00138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16302_ (.A0(_02661_),
    .A1(_02656_),
    .S(_01337_),
    .X(_00137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16303_ (.A0(_02651_),
    .A1(_02646_),
    .S(_01337_),
    .X(_00136_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16304_ (.A0(_02641_),
    .A1(_02636_),
    .S(_01337_),
    .X(_00135_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16305_ (.A0(_02631_),
    .A1(_02626_),
    .S(_01337_),
    .X(_00134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16306_ (.A0(_02621_),
    .A1(_02616_),
    .S(_01337_),
    .X(_00131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16307_ (.A0(_02611_),
    .A1(_02606_),
    .S(_01337_),
    .X(_00120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16308_ (.A0(_02601_),
    .A1(_02596_),
    .S(_01337_),
    .X(_00109_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16309_ (.A0(_02585_),
    .A1(\design_top.DADDR[31] ),
    .S(_00821_),
    .X(_02586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16310_ (.A0(_02586_),
    .A1(_02583_),
    .S(_01329_),
    .X(_00101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16311_ (.A0(_02580_),
    .A1(_02581_),
    .S(_00821_),
    .X(_02582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16312_ (.A0(_02582_),
    .A1(_02579_),
    .S(_01329_),
    .X(_00100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16313_ (.A0(_02576_),
    .A1(_02577_),
    .S(_00821_),
    .X(_02578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16314_ (.A0(_02578_),
    .A1(_02575_),
    .S(_01329_),
    .X(_00098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16315_ (.A0(_02572_),
    .A1(_02573_),
    .S(_00821_),
    .X(_02574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16316_ (.A0(_02574_),
    .A1(_02571_),
    .S(_01329_),
    .X(_00097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16317_ (.A0(_02568_),
    .A1(_02569_),
    .S(_00821_),
    .X(_02570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16318_ (.A0(_02570_),
    .A1(_02567_),
    .S(_01329_),
    .X(_00096_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16319_ (.A0(_02564_),
    .A1(_02565_),
    .S(_00821_),
    .X(_02566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16320_ (.A0(_02566_),
    .A1(_02563_),
    .S(_01329_),
    .X(_00095_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16321_ (.A0(_02560_),
    .A1(_02561_),
    .S(_00821_),
    .X(_02562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16322_ (.A0(_02562_),
    .A1(_02559_),
    .S(_01329_),
    .X(_00094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16323_ (.A0(_02556_),
    .A1(_02557_),
    .S(_00821_),
    .X(_02558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16324_ (.A0(_02558_),
    .A1(_02555_),
    .S(_01329_),
    .X(_00093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16325_ (.A0(_02552_),
    .A1(_02553_),
    .S(_00821_),
    .X(_02554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16326_ (.A0(_02554_),
    .A1(_02551_),
    .S(_01329_),
    .X(_00092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16327_ (.A0(_02548_),
    .A1(_02549_),
    .S(_00821_),
    .X(_02550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16328_ (.A0(_02550_),
    .A1(_02547_),
    .S(_01329_),
    .X(_00091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16329_ (.A0(_02544_),
    .A1(_02545_),
    .S(_00821_),
    .X(_02546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16330_ (.A0(_02546_),
    .A1(_02543_),
    .S(_01329_),
    .X(_00090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16331_ (.A0(_02540_),
    .A1(_02541_),
    .S(_00821_),
    .X(_02542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16332_ (.A0(_02542_),
    .A1(_02539_),
    .S(_01329_),
    .X(_00089_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16333_ (.A0(_02536_),
    .A1(_02537_),
    .S(_00821_),
    .X(_02538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16334_ (.A0(_02538_),
    .A1(_02535_),
    .S(_01329_),
    .X(_00088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16335_ (.A0(_02532_),
    .A1(_02533_),
    .S(_00821_),
    .X(_02534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16336_ (.A0(_02534_),
    .A1(_02531_),
    .S(_01329_),
    .X(_00087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16337_ (.A0(_02528_),
    .A1(_02529_),
    .S(_00821_),
    .X(_02530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16338_ (.A0(_02530_),
    .A1(_02527_),
    .S(_01329_),
    .X(_00086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16339_ (.A0(_02524_),
    .A1(_02525_),
    .S(_00821_),
    .X(_02526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16340_ (.A0(_02526_),
    .A1(_02523_),
    .S(_01329_),
    .X(_00085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16341_ (.A0(_02520_),
    .A1(_02521_),
    .S(_00821_),
    .X(_02522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16342_ (.A0(_02522_),
    .A1(_02519_),
    .S(_01329_),
    .X(_00084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16343_ (.A0(_02516_),
    .A1(_02517_),
    .S(_00821_),
    .X(_02518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16344_ (.A0(_02518_),
    .A1(_02515_),
    .S(_01329_),
    .X(_00083_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16345_ (.A0(_02512_),
    .A1(_02513_),
    .S(_00821_),
    .X(_02514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16346_ (.A0(_02514_),
    .A1(_02511_),
    .S(_01329_),
    .X(_00082_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16347_ (.A0(_02508_),
    .A1(_02509_),
    .S(_00821_),
    .X(_02510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16348_ (.A0(_02510_),
    .A1(_02507_),
    .S(_01329_),
    .X(_00081_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16349_ (.A0(_02504_),
    .A1(_02505_),
    .S(_00821_),
    .X(_02506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16350_ (.A0(_02506_),
    .A1(_02503_),
    .S(_01329_),
    .X(_00080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16351_ (.A0(_02500_),
    .A1(_02501_),
    .S(_00821_),
    .X(_02502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16352_ (.A0(_02502_),
    .A1(_02499_),
    .S(_01329_),
    .X(_00079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16353_ (.A0(_02496_),
    .A1(_02497_),
    .S(_00821_),
    .X(_02498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16354_ (.A0(_02498_),
    .A1(_02495_),
    .S(_01329_),
    .X(_00108_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16355_ (.A0(_02492_),
    .A1(_02493_),
    .S(_00821_),
    .X(_02494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16356_ (.A0(_02494_),
    .A1(_02491_),
    .S(_01329_),
    .X(_00107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16357_ (.A0(_02488_),
    .A1(_02489_),
    .S(_00821_),
    .X(_02490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16358_ (.A0(_02490_),
    .A1(_02487_),
    .S(_01329_),
    .X(_00106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16359_ (.A0(_02485_),
    .A1(_02484_),
    .S(_00821_),
    .X(_02486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16360_ (.A0(_02486_),
    .A1(_02483_),
    .S(_01329_),
    .X(_00105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16361_ (.A0(_02481_),
    .A1(_02480_),
    .S(_00821_),
    .X(_02482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16362_ (.A0(_02482_),
    .A1(_02479_),
    .S(_01329_),
    .X(_00104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16363_ (.A0(_02477_),
    .A1(_01371_),
    .S(_00821_),
    .X(_02478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16364_ (.A0(_02478_),
    .A1(_02476_),
    .S(_01329_),
    .X(_00103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16365_ (.A0(_02474_),
    .A1(\design_top.DADDR[3] ),
    .S(_00821_),
    .X(_02475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16366_ (.A0(_02475_),
    .A1(_02473_),
    .S(_01329_),
    .X(_00102_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16367_ (.A0(_02471_),
    .A1(\design_top.DADDR[2] ),
    .S(_00821_),
    .X(_02472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16368_ (.A0(_02472_),
    .A1(_02470_),
    .S(_01329_),
    .X(_00099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16369_ (.A0(_02097_),
    .A1(_02098_),
    .S(\design_top.core0.XRES ),
    .X(_00045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16370_ (.A0(_01519_),
    .A1(_01518_),
    .S(_00786_),
    .X(_00011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_1 _16371_ (.A0(_01517_),
    .A1(_01331_),
    .S(_01330_),
    .X(_00078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16372_ (.A0(\design_top.uart0.UART_XFIFO[0] ),
    .A1(\design_top.uart0.UART_XFIFO[1] ),
    .A2(\design_top.uart0.UART_XFIFO[2] ),
    .A3(\design_top.uart0.UART_XFIFO[3] ),
    .S0(\design_top.uart0.UART_XSTATE[0] ),
    .S1(\design_top.uart0.UART_XSTATE[1] ),
    .X(_02588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16373_ (.A0(\design_top.uart0.UART_XFIFO[4] ),
    .A1(\design_top.uart0.UART_XFIFO[5] ),
    .A2(\design_top.uart0.UART_XFIFO[6] ),
    .A3(\design_top.uart0.UART_XFIFO[7] ),
    .S0(\design_top.uart0.UART_XSTATE[0] ),
    .S1(\design_top.uart0.UART_XSTATE[1] ),
    .X(_02589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16374_ (.A0(_00776_),
    .A1(_00851_),
    .A2(_01974_),
    .A3(_00777_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_00778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16375_ (.A0(_00772_),
    .A1(_00770_),
    .A2(_00764_),
    .A3(_00765_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_00773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16376_ (.A0(_02461_),
    .A1(_00865_),
    .A2(_01974_),
    .A3(_02462_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16377_ (.A0(_02457_),
    .A1(_02454_),
    .A2(_02448_),
    .A3(_02449_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16378_ (.A0(_02440_),
    .A1(_00879_),
    .A2(_01974_),
    .A3(_02441_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16379_ (.A0(_02436_),
    .A1(_02433_),
    .A2(_02427_),
    .A3(_02428_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16380_ (.A0(_02419_),
    .A1(_02405_),
    .A2(_01974_),
    .A3(_02420_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02421_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16381_ (.A0(_02415_),
    .A1(_02412_),
    .A2(_02406_),
    .A3(_02407_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02416_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16382_ (.A0(_02397_),
    .A1(_00906_),
    .A2(_01974_),
    .A3(_02398_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02399_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16383_ (.A0(_02393_),
    .A1(_02390_),
    .A2(_02384_),
    .A3(_02385_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02394_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16384_ (.A0(_02376_),
    .A1(_02362_),
    .A2(_01974_),
    .A3(_02377_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02378_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16385_ (.A0(_02372_),
    .A1(_02369_),
    .A2(_02363_),
    .A3(_02364_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02373_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16386_ (.A0(_02354_),
    .A1(_00933_),
    .A2(_01974_),
    .A3(_02355_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02356_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16387_ (.A0(_02350_),
    .A1(_02347_),
    .A2(_02341_),
    .A3(_02342_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02351_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16388_ (.A0(_02333_),
    .A1(_02319_),
    .A2(_01974_),
    .A3(_02334_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02335_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16389_ (.A0(_02329_),
    .A1(_02326_),
    .A2(_02320_),
    .A3(_02321_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02330_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16390_ (.A0(_02311_),
    .A1(_00960_),
    .A2(_01974_),
    .A3(_02312_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02313_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16391_ (.A0(_02307_),
    .A1(_02304_),
    .A2(_02298_),
    .A3(_02299_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02308_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16392_ (.A0(_02290_),
    .A1(_02276_),
    .A2(_01974_),
    .A3(_02291_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02292_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16393_ (.A0(_02286_),
    .A1(_02283_),
    .A2(_02277_),
    .A3(_02278_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02287_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16394_ (.A0(_02268_),
    .A1(_00987_),
    .A2(_01974_),
    .A3(_02269_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02270_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16395_ (.A0(_02264_),
    .A1(_02261_),
    .A2(_02255_),
    .A3(_02256_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02265_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16396_ (.A0(_02247_),
    .A1(_02233_),
    .A2(_01974_),
    .A3(_02248_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16397_ (.A0(_02243_),
    .A1(_02240_),
    .A2(_02234_),
    .A3(_02235_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16398_ (.A0(_02225_),
    .A1(_01014_),
    .A2(_01974_),
    .A3(_02226_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16399_ (.A0(_02221_),
    .A1(_02218_),
    .A2(_02212_),
    .A3(_02213_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16400_ (.A0(_02204_),
    .A1(_02190_),
    .A2(_01974_),
    .A3(_02205_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16401_ (.A0(_02200_),
    .A1(_02197_),
    .A2(_02191_),
    .A3(_02192_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16402_ (.A0(_02182_),
    .A1(_01056_),
    .A2(_01974_),
    .A3(_02183_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02184_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16403_ (.A0(_02178_),
    .A1(_02175_),
    .A2(_02169_),
    .A3(_02170_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16404_ (.A0(_02160_),
    .A1(_02146_),
    .A2(_01974_),
    .A3(_02162_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02163_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16405_ (.A0(_02156_),
    .A1(_02153_),
    .A2(_02147_),
    .A3(_02148_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16406_ (.A0(_02137_),
    .A1(_01083_),
    .A2(_01974_),
    .A3(_02139_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16407_ (.A0(_02131_),
    .A1(_02132_),
    .A2(_02131_),
    .A3(_00843_),
    .S0(_01230_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_02133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16408_ (.A0(_02133_),
    .A1(_02130_),
    .A2(_02124_),
    .A3(_02125_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02134_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16409_ (.A0(_02115_),
    .A1(_02100_),
    .A2(_01974_),
    .A3(_02117_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16410_ (.A0(_02108_),
    .A1(_02109_),
    .A2(_02108_),
    .A3(_02110_),
    .S0(_01230_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_02111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16411_ (.A0(_02111_),
    .A1(_02107_),
    .A2(_02101_),
    .A3(_02102_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16412_ (.A0(_02089_),
    .A1(_01110_),
    .A2(_01974_),
    .A3(_02091_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16413_ (.A0(_02082_),
    .A1(_02083_),
    .A2(_02082_),
    .A3(_02084_),
    .S0(_01230_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_02085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16414_ (.A0(_02085_),
    .A1(_02081_),
    .A2(_02075_),
    .A3(_02076_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16415_ (.A0(_02066_),
    .A1(_02051_),
    .A2(_01974_),
    .A3(_02068_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02069_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16416_ (.A0(_02059_),
    .A1(_02060_),
    .A2(_02059_),
    .A3(_02061_),
    .S0(_01230_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_02062_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16417_ (.A0(_02062_),
    .A1(_02058_),
    .A2(_02052_),
    .A3(_02053_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16418_ (.A0(_02042_),
    .A1(_01136_),
    .A2(_01974_),
    .A3(_02044_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16419_ (.A0(_02035_),
    .A1(_02036_),
    .A2(_02035_),
    .A3(_02037_),
    .S0(_01230_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_02038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16420_ (.A0(_02038_),
    .A1(_02034_),
    .A2(_02028_),
    .A3(_02029_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16421_ (.A0(_02019_),
    .A1(_02004_),
    .A2(_01974_),
    .A3(_02021_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_02022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16422_ (.A0(_02012_),
    .A1(_02013_),
    .A2(_02012_),
    .A3(_02014_),
    .S0(_01230_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_02015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16423_ (.A0(_02015_),
    .A1(_02011_),
    .A2(_02005_),
    .A3(_02006_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_02016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16424_ (.A0(_01995_),
    .A1(_01165_),
    .A2(_01974_),
    .A3(_01997_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_01998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16425_ (.A0(_01988_),
    .A1(_01989_),
    .A2(_01988_),
    .A3(_01990_),
    .S0(_01230_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16426_ (.A0(_01991_),
    .A1(_01987_),
    .A2(_01981_),
    .A3(_01982_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_01992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16427_ (.A0(_01971_),
    .A1(_01956_),
    .A2(_01974_),
    .A3(_01973_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_01975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16428_ (.A0(_01964_),
    .A1(_01965_),
    .A2(_01964_),
    .A3(_01966_),
    .S0(_01230_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16429_ (.A0(_01967_),
    .A1(_01963_),
    .A2(_01957_),
    .A3(_01958_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_01968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16430_ (.A0(_01931_),
    .A1(_01192_),
    .A2(_01949_),
    .A3(_01939_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_01950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16431_ (.A0(_01922_),
    .A1(_01925_),
    .A2(_01922_),
    .A3(_01926_),
    .S0(_01230_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16432_ (.A0(_01927_),
    .A1(_01919_),
    .A2(_01913_),
    .A3(_01914_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_01928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16433_ (.A0(_01888_),
    .A1(_01868_),
    .A2(_01906_),
    .A3(_01897_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_01907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16434_ (.A0(_01878_),
    .A1(_01881_),
    .A2(_01878_),
    .A3(_01883_),
    .S0(_01230_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16435_ (.A0(_01884_),
    .A1(_01875_),
    .A2(_01869_),
    .A3(_01870_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_01885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16436_ (.A0(_01843_),
    .A1(_01218_),
    .A2(_01861_),
    .A3(_01852_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_01862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16437_ (.A0(_01833_),
    .A1(_01836_),
    .A2(_01833_),
    .A3(_01838_),
    .S0(_01230_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16438_ (.A0(_01839_),
    .A1(_01830_),
    .A2(_01824_),
    .A3(_01825_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_01840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16439_ (.A0(_01800_),
    .A1(_01780_),
    .A2(_01817_),
    .A3(_01808_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_01818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16440_ (.A0(_01790_),
    .A1(_01793_),
    .A2(_01790_),
    .A3(_01795_),
    .S0(_01230_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16441_ (.A0(_01796_),
    .A1(_01787_),
    .A2(_01781_),
    .A3(_01782_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_01797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16442_ (.A0(_01756_),
    .A1(_01240_),
    .A2(_01773_),
    .A3(_01764_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_01774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16443_ (.A0(_01742_),
    .A1(_01749_),
    .A2(_01742_),
    .A3(_01751_),
    .S0(_01230_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16444_ (.A0(_01752_),
    .A1(_01735_),
    .A2(_01729_),
    .A3(_01730_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_01753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16445_ (.A0(_01704_),
    .A1(_01675_),
    .A2(_01722_),
    .A3(_01713_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_01723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16446_ (.A0(_01689_),
    .A1(_01696_),
    .A2(_01689_),
    .A3(_01699_),
    .S0(_01230_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16447_ (.A0(_01700_),
    .A1(_01682_),
    .A2(_01676_),
    .A3(_01677_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_01701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16448_ (.A0(_01650_),
    .A1(_01604_),
    .A2(_01668_),
    .A3(_01658_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_01669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16449_ (.A0(_01627_),
    .A1(_01642_),
    .A2(_01627_),
    .A3(_01645_),
    .S0(_01230_),
    .S1(\design_top.core0.FCT7[5] ),
    .X(_01646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16450_ (.A0(_01646_),
    .A1(_01612_),
    .A2(_01606_),
    .A3(_01607_),
    .S0(_08562_),
    .S1(_01323_),
    .X(_01647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16451_ (.A0(_01570_),
    .A1(_01521_),
    .A2(_01591_),
    .A3(_01580_),
    .S0(_08561_),
    .S1(io_out[12]),
    .X(_01592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16452_ (.A0(\design_top.core0.REG2[0][0] ),
    .A1(\design_top.core0.REG2[1][0] ),
    .A2(\design_top.core0.REG2[2][0] ),
    .A3(\design_top.core0.REG2[3][0] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01256_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16453_ (.A0(\design_top.core0.REG2[4][0] ),
    .A1(\design_top.core0.REG2[5][0] ),
    .A2(\design_top.core0.REG2[6][0] ),
    .A3(\design_top.core0.REG2[7][0] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01257_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16454_ (.A0(\design_top.core0.REG2[8][0] ),
    .A1(\design_top.core0.REG2[9][0] ),
    .A2(\design_top.core0.REG2[10][0] ),
    .A3(\design_top.core0.REG2[11][0] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01258_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16455_ (.A0(\design_top.core0.REG2[12][0] ),
    .A1(\design_top.core0.REG2[13][0] ),
    .A2(\design_top.core0.REG2[14][0] ),
    .A3(\design_top.core0.REG2[15][0] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01259_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16456_ (.A0(_01256_),
    .A1(_01257_),
    .A2(_01258_),
    .A3(_01259_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_01260_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16457_ (.A0(\design_top.core0.REG2[0][1] ),
    .A1(\design_top.core0.REG2[1][1] ),
    .A2(\design_top.core0.REG2[2][1] ),
    .A3(\design_top.core0.REG2[3][1] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01249_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16458_ (.A0(\design_top.core0.REG2[4][1] ),
    .A1(\design_top.core0.REG2[5][1] ),
    .A2(\design_top.core0.REG2[6][1] ),
    .A3(\design_top.core0.REG2[7][1] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01250_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16459_ (.A0(\design_top.core0.REG2[8][1] ),
    .A1(\design_top.core0.REG2[9][1] ),
    .A2(\design_top.core0.REG2[10][1] ),
    .A3(\design_top.core0.REG2[11][1] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01251_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16460_ (.A0(\design_top.core0.REG2[12][1] ),
    .A1(\design_top.core0.REG2[13][1] ),
    .A2(\design_top.core0.REG2[14][1] ),
    .A3(\design_top.core0.REG2[15][1] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01252_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16461_ (.A0(_01249_),
    .A1(_01250_),
    .A2(_01251_),
    .A3(_01252_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_01253_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16462_ (.A0(\design_top.core0.REG2[0][2] ),
    .A1(\design_top.core0.REG2[1][2] ),
    .A2(\design_top.core0.REG2[2][2] ),
    .A3(\design_top.core0.REG2[3][2] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01241_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16463_ (.A0(\design_top.core0.REG2[4][2] ),
    .A1(\design_top.core0.REG2[5][2] ),
    .A2(\design_top.core0.REG2[6][2] ),
    .A3(\design_top.core0.REG2[7][2] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01242_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16464_ (.A0(\design_top.core0.REG2[8][2] ),
    .A1(\design_top.core0.REG2[9][2] ),
    .A2(\design_top.core0.REG2[10][2] ),
    .A3(\design_top.core0.REG2[11][2] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01243_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16465_ (.A0(\design_top.core0.REG2[12][2] ),
    .A1(\design_top.core0.REG2[13][2] ),
    .A2(\design_top.core0.REG2[14][2] ),
    .A3(\design_top.core0.REG2[15][2] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01244_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16466_ (.A0(_01241_),
    .A1(_01242_),
    .A2(_01243_),
    .A3(_01244_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_01245_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16467_ (.A0(\design_top.core0.REG2[0][3] ),
    .A1(\design_top.core0.REG2[1][3] ),
    .A2(\design_top.core0.REG2[2][3] ),
    .A3(\design_top.core0.REG2[3][3] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01233_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16468_ (.A0(\design_top.core0.REG2[4][3] ),
    .A1(\design_top.core0.REG2[5][3] ),
    .A2(\design_top.core0.REG2[6][3] ),
    .A3(\design_top.core0.REG2[7][3] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01234_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16469_ (.A0(\design_top.core0.REG2[8][3] ),
    .A1(\design_top.core0.REG2[9][3] ),
    .A2(\design_top.core0.REG2[10][3] ),
    .A3(\design_top.core0.REG2[11][3] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01235_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16470_ (.A0(\design_top.core0.REG2[12][3] ),
    .A1(\design_top.core0.REG2[13][3] ),
    .A2(\design_top.core0.REG2[14][3] ),
    .A3(\design_top.core0.REG2[15][3] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01236_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16471_ (.A0(_01233_),
    .A1(_01234_),
    .A2(_01235_),
    .A3(_01236_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_01237_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16472_ (.A0(\design_top.core0.REG2[0][4] ),
    .A1(\design_top.core0.REG2[1][4] ),
    .A2(\design_top.core0.REG2[2][4] ),
    .A3(\design_top.core0.REG2[3][4] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01225_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16473_ (.A0(\design_top.core0.REG2[4][4] ),
    .A1(\design_top.core0.REG2[5][4] ),
    .A2(\design_top.core0.REG2[6][4] ),
    .A3(\design_top.core0.REG2[7][4] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01226_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16474_ (.A0(\design_top.core0.REG2[8][4] ),
    .A1(\design_top.core0.REG2[9][4] ),
    .A2(\design_top.core0.REG2[10][4] ),
    .A3(\design_top.core0.REG2[11][4] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01227_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16475_ (.A0(\design_top.core0.REG2[12][4] ),
    .A1(\design_top.core0.REG2[13][4] ),
    .A2(\design_top.core0.REG2[14][4] ),
    .A3(\design_top.core0.REG2[15][4] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01228_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16476_ (.A0(_01225_),
    .A1(_01226_),
    .A2(_01227_),
    .A3(_01228_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_01229_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16477_ (.A0(\design_top.core0.REG1[0][4] ),
    .A1(\design_top.core0.REG1[1][4] ),
    .A2(\design_top.core0.REG1[2][4] ),
    .A3(\design_top.core0.REG1[3][4] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01219_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16478_ (.A0(\design_top.core0.REG1[4][4] ),
    .A1(\design_top.core0.REG1[5][4] ),
    .A2(\design_top.core0.REG1[6][4] ),
    .A3(\design_top.core0.REG1[7][4] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01220_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16479_ (.A0(\design_top.core0.REG1[8][4] ),
    .A1(\design_top.core0.REG1[9][4] ),
    .A2(\design_top.core0.REG1[10][4] ),
    .A3(\design_top.core0.REG1[11][4] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01221_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16480_ (.A0(\design_top.core0.REG1[12][4] ),
    .A1(\design_top.core0.REG1[13][4] ),
    .A2(\design_top.core0.REG1[14][4] ),
    .A3(\design_top.core0.REG1[15][4] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01222_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16481_ (.A0(_01219_),
    .A1(_01220_),
    .A2(_01221_),
    .A3(_01222_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_01223_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16482_ (.A0(\design_top.core0.REG2[0][5] ),
    .A1(\design_top.core0.REG2[1][5] ),
    .A2(\design_top.core0.REG2[2][5] ),
    .A3(\design_top.core0.REG2[3][5] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01211_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16483_ (.A0(\design_top.core0.REG2[4][5] ),
    .A1(\design_top.core0.REG2[5][5] ),
    .A2(\design_top.core0.REG2[6][5] ),
    .A3(\design_top.core0.REG2[7][5] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01212_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16484_ (.A0(\design_top.core0.REG2[8][5] ),
    .A1(\design_top.core0.REG2[9][5] ),
    .A2(\design_top.core0.REG2[10][5] ),
    .A3(\design_top.core0.REG2[11][5] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01213_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16485_ (.A0(\design_top.core0.REG2[12][5] ),
    .A1(\design_top.core0.REG2[13][5] ),
    .A2(\design_top.core0.REG2[14][5] ),
    .A3(\design_top.core0.REG2[15][5] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01214_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16486_ (.A0(_01211_),
    .A1(_01212_),
    .A2(_01213_),
    .A3(_01214_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_01215_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16487_ (.A0(\design_top.core0.REG1[0][5] ),
    .A1(\design_top.core0.REG1[1][5] ),
    .A2(\design_top.core0.REG1[2][5] ),
    .A3(\design_top.core0.REG1[3][5] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01206_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16488_ (.A0(\design_top.core0.REG1[4][5] ),
    .A1(\design_top.core0.REG1[5][5] ),
    .A2(\design_top.core0.REG1[6][5] ),
    .A3(\design_top.core0.REG1[7][5] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01207_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16489_ (.A0(\design_top.core0.REG1[8][5] ),
    .A1(\design_top.core0.REG1[9][5] ),
    .A2(\design_top.core0.REG1[10][5] ),
    .A3(\design_top.core0.REG1[11][5] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01208_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16490_ (.A0(\design_top.core0.REG1[12][5] ),
    .A1(\design_top.core0.REG1[13][5] ),
    .A2(\design_top.core0.REG1[14][5] ),
    .A3(\design_top.core0.REG1[15][5] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01209_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16491_ (.A0(_01206_),
    .A1(_01207_),
    .A2(_01208_),
    .A3(_01209_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_01210_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16492_ (.A0(\design_top.core0.REG2[0][6] ),
    .A1(\design_top.core0.REG2[1][6] ),
    .A2(\design_top.core0.REG2[2][6] ),
    .A3(\design_top.core0.REG2[3][6] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01199_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16493_ (.A0(\design_top.core0.REG2[4][6] ),
    .A1(\design_top.core0.REG2[5][6] ),
    .A2(\design_top.core0.REG2[6][6] ),
    .A3(\design_top.core0.REG2[7][6] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01200_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16494_ (.A0(\design_top.core0.REG2[8][6] ),
    .A1(\design_top.core0.REG2[9][6] ),
    .A2(\design_top.core0.REG2[10][6] ),
    .A3(\design_top.core0.REG2[11][6] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01201_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16495_ (.A0(\design_top.core0.REG2[12][6] ),
    .A1(\design_top.core0.REG2[13][6] ),
    .A2(\design_top.core0.REG2[14][6] ),
    .A3(\design_top.core0.REG2[15][6] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01202_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16496_ (.A0(_01199_),
    .A1(_01200_),
    .A2(_01201_),
    .A3(_01202_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_01203_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16497_ (.A0(\design_top.core0.REG1[0][6] ),
    .A1(\design_top.core0.REG1[1][6] ),
    .A2(\design_top.core0.REG1[2][6] ),
    .A3(\design_top.core0.REG1[3][6] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01193_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16498_ (.A0(\design_top.core0.REG1[4][6] ),
    .A1(\design_top.core0.REG1[5][6] ),
    .A2(\design_top.core0.REG1[6][6] ),
    .A3(\design_top.core0.REG1[7][6] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01194_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16499_ (.A0(\design_top.core0.REG1[8][6] ),
    .A1(\design_top.core0.REG1[9][6] ),
    .A2(\design_top.core0.REG1[10][6] ),
    .A3(\design_top.core0.REG1[11][6] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01195_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16500_ (.A0(\design_top.core0.REG1[12][6] ),
    .A1(\design_top.core0.REG1[13][6] ),
    .A2(\design_top.core0.REG1[14][6] ),
    .A3(\design_top.core0.REG1[15][6] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01196_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16501_ (.A0(_01193_),
    .A1(_01194_),
    .A2(_01195_),
    .A3(_01196_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_01197_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16502_ (.A0(\design_top.core0.REG2[0][7] ),
    .A1(\design_top.core0.REG2[1][7] ),
    .A2(\design_top.core0.REG2[2][7] ),
    .A3(\design_top.core0.REG2[3][7] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01185_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16503_ (.A0(\design_top.core0.REG2[4][7] ),
    .A1(\design_top.core0.REG2[5][7] ),
    .A2(\design_top.core0.REG2[6][7] ),
    .A3(\design_top.core0.REG2[7][7] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01186_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16504_ (.A0(\design_top.core0.REG2[8][7] ),
    .A1(\design_top.core0.REG2[9][7] ),
    .A2(\design_top.core0.REG2[10][7] ),
    .A3(\design_top.core0.REG2[11][7] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01187_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16505_ (.A0(\design_top.core0.REG2[12][7] ),
    .A1(\design_top.core0.REG2[13][7] ),
    .A2(\design_top.core0.REG2[14][7] ),
    .A3(\design_top.core0.REG2[15][7] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01188_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16506_ (.A0(_01185_),
    .A1(_01186_),
    .A2(_01187_),
    .A3(_01188_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_01189_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16507_ (.A0(\design_top.core0.REG1[0][7] ),
    .A1(\design_top.core0.REG1[1][7] ),
    .A2(\design_top.core0.REG1[2][7] ),
    .A3(\design_top.core0.REG1[3][7] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01179_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16508_ (.A0(\design_top.core0.REG1[4][7] ),
    .A1(\design_top.core0.REG1[5][7] ),
    .A2(\design_top.core0.REG1[6][7] ),
    .A3(\design_top.core0.REG1[7][7] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01180_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16509_ (.A0(\design_top.core0.REG1[8][7] ),
    .A1(\design_top.core0.REG1[9][7] ),
    .A2(\design_top.core0.REG1[10][7] ),
    .A3(\design_top.core0.REG1[11][7] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01181_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16510_ (.A0(\design_top.core0.REG1[12][7] ),
    .A1(\design_top.core0.REG1[13][7] ),
    .A2(\design_top.core0.REG1[14][7] ),
    .A3(\design_top.core0.REG1[15][7] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01182_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16511_ (.A0(_01179_),
    .A1(_01180_),
    .A2(_01181_),
    .A3(_01182_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_01183_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16512_ (.A0(\design_top.core0.REG2[0][8] ),
    .A1(\design_top.core0.REG2[1][8] ),
    .A2(\design_top.core0.REG2[2][8] ),
    .A3(\design_top.core0.REG2[3][8] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01172_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16513_ (.A0(\design_top.core0.REG2[4][8] ),
    .A1(\design_top.core0.REG2[5][8] ),
    .A2(\design_top.core0.REG2[6][8] ),
    .A3(\design_top.core0.REG2[7][8] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01173_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16514_ (.A0(\design_top.core0.REG2[8][8] ),
    .A1(\design_top.core0.REG2[9][8] ),
    .A2(\design_top.core0.REG2[10][8] ),
    .A3(\design_top.core0.REG2[11][8] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01174_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16515_ (.A0(\design_top.core0.REG2[12][8] ),
    .A1(\design_top.core0.REG2[13][8] ),
    .A2(\design_top.core0.REG2[14][8] ),
    .A3(\design_top.core0.REG2[15][8] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01175_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16516_ (.A0(_01172_),
    .A1(_01173_),
    .A2(_01174_),
    .A3(_01175_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_01176_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16517_ (.A0(\design_top.core0.REG1[0][8] ),
    .A1(\design_top.core0.REG1[1][8] ),
    .A2(\design_top.core0.REG1[2][8] ),
    .A3(\design_top.core0.REG1[3][8] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01166_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16518_ (.A0(\design_top.core0.REG1[4][8] ),
    .A1(\design_top.core0.REG1[5][8] ),
    .A2(\design_top.core0.REG1[6][8] ),
    .A3(\design_top.core0.REG1[7][8] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01167_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16519_ (.A0(\design_top.core0.REG1[8][8] ),
    .A1(\design_top.core0.REG1[9][8] ),
    .A2(\design_top.core0.REG1[10][8] ),
    .A3(\design_top.core0.REG1[11][8] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01168_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16520_ (.A0(\design_top.core0.REG1[12][8] ),
    .A1(\design_top.core0.REG1[13][8] ),
    .A2(\design_top.core0.REG1[14][8] ),
    .A3(\design_top.core0.REG1[15][8] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01169_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16521_ (.A0(_01166_),
    .A1(_01167_),
    .A2(_01168_),
    .A3(_01169_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_01170_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16522_ (.A0(\design_top.core0.REG2[0][9] ),
    .A1(\design_top.core0.REG2[1][9] ),
    .A2(\design_top.core0.REG2[2][9] ),
    .A3(\design_top.core0.REG2[3][9] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01157_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16523_ (.A0(\design_top.core0.REG2[4][9] ),
    .A1(\design_top.core0.REG2[5][9] ),
    .A2(\design_top.core0.REG2[6][9] ),
    .A3(\design_top.core0.REG2[7][9] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01158_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16524_ (.A0(\design_top.core0.REG2[8][9] ),
    .A1(\design_top.core0.REG2[9][9] ),
    .A2(\design_top.core0.REG2[10][9] ),
    .A3(\design_top.core0.REG2[11][9] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01159_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16525_ (.A0(\design_top.core0.REG2[12][9] ),
    .A1(\design_top.core0.REG2[13][9] ),
    .A2(\design_top.core0.REG2[14][9] ),
    .A3(\design_top.core0.REG2[15][9] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01160_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16526_ (.A0(_01157_),
    .A1(_01158_),
    .A2(_01159_),
    .A3(_01160_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_01161_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16527_ (.A0(\design_top.core0.REG1[8][9] ),
    .A1(\design_top.core0.REG1[9][9] ),
    .A2(\design_top.core0.REG1[10][9] ),
    .A3(\design_top.core0.REG1[11][9] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01153_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16528_ (.A0(\design_top.core0.REG1[12][9] ),
    .A1(\design_top.core0.REG1[13][9] ),
    .A2(\design_top.core0.REG1[14][9] ),
    .A3(\design_top.core0.REG1[15][9] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01154_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16529_ (.A0(\design_top.core0.REG1[0][9] ),
    .A1(\design_top.core0.REG1[1][9] ),
    .A2(\design_top.core0.REG1[2][9] ),
    .A3(\design_top.core0.REG1[3][9] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01150_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16530_ (.A0(\design_top.core0.REG1[4][9] ),
    .A1(\design_top.core0.REG1[5][9] ),
    .A2(\design_top.core0.REG1[6][9] ),
    .A3(\design_top.core0.REG1[7][9] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01151_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16531_ (.A0(\design_top.core0.REG2[0][10] ),
    .A1(\design_top.core0.REG2[1][10] ),
    .A2(\design_top.core0.REG2[2][10] ),
    .A3(\design_top.core0.REG2[3][10] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01143_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16532_ (.A0(\design_top.core0.REG2[4][10] ),
    .A1(\design_top.core0.REG2[5][10] ),
    .A2(\design_top.core0.REG2[6][10] ),
    .A3(\design_top.core0.REG2[7][10] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01144_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16533_ (.A0(\design_top.core0.REG2[8][10] ),
    .A1(\design_top.core0.REG2[9][10] ),
    .A2(\design_top.core0.REG2[10][10] ),
    .A3(\design_top.core0.REG2[11][10] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01145_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16534_ (.A0(\design_top.core0.REG2[12][10] ),
    .A1(\design_top.core0.REG2[13][10] ),
    .A2(\design_top.core0.REG2[14][10] ),
    .A3(\design_top.core0.REG2[15][10] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01146_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16535_ (.A0(_01143_),
    .A1(_01144_),
    .A2(_01145_),
    .A3(_01146_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_01147_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16536_ (.A0(\design_top.core0.REG1[0][10] ),
    .A1(\design_top.core0.REG1[1][10] ),
    .A2(\design_top.core0.REG1[2][10] ),
    .A3(\design_top.core0.REG1[3][10] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01137_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16537_ (.A0(\design_top.core0.REG1[4][10] ),
    .A1(\design_top.core0.REG1[5][10] ),
    .A2(\design_top.core0.REG1[6][10] ),
    .A3(\design_top.core0.REG1[7][10] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01138_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16538_ (.A0(\design_top.core0.REG1[8][10] ),
    .A1(\design_top.core0.REG1[9][10] ),
    .A2(\design_top.core0.REG1[10][10] ),
    .A3(\design_top.core0.REG1[11][10] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01139_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16539_ (.A0(\design_top.core0.REG1[12][10] ),
    .A1(\design_top.core0.REG1[13][10] ),
    .A2(\design_top.core0.REG1[14][10] ),
    .A3(\design_top.core0.REG1[15][10] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01140_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16540_ (.A0(_01137_),
    .A1(_01138_),
    .A2(_01139_),
    .A3(_01140_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_01141_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16541_ (.A0(\design_top.core0.REG2[0][11] ),
    .A1(\design_top.core0.REG2[1][11] ),
    .A2(\design_top.core0.REG2[2][11] ),
    .A3(\design_top.core0.REG2[3][11] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01129_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16542_ (.A0(\design_top.core0.REG2[4][11] ),
    .A1(\design_top.core0.REG2[5][11] ),
    .A2(\design_top.core0.REG2[6][11] ),
    .A3(\design_top.core0.REG2[7][11] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01130_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16543_ (.A0(\design_top.core0.REG2[8][11] ),
    .A1(\design_top.core0.REG2[9][11] ),
    .A2(\design_top.core0.REG2[10][11] ),
    .A3(\design_top.core0.REG2[11][11] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01131_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16544_ (.A0(\design_top.core0.REG2[12][11] ),
    .A1(\design_top.core0.REG2[13][11] ),
    .A2(\design_top.core0.REG2[14][11] ),
    .A3(\design_top.core0.REG2[15][11] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01132_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16545_ (.A0(_01129_),
    .A1(_01130_),
    .A2(_01131_),
    .A3(_01132_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_01133_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16546_ (.A0(\design_top.core0.REG1[0][11] ),
    .A1(\design_top.core0.REG1[1][11] ),
    .A2(\design_top.core0.REG1[2][11] ),
    .A3(\design_top.core0.REG1[3][11] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01124_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16547_ (.A0(\design_top.core0.REG1[4][11] ),
    .A1(\design_top.core0.REG1[5][11] ),
    .A2(\design_top.core0.REG1[6][11] ),
    .A3(\design_top.core0.REG1[7][11] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01125_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16548_ (.A0(\design_top.core0.REG1[8][11] ),
    .A1(\design_top.core0.REG1[9][11] ),
    .A2(\design_top.core0.REG1[10][11] ),
    .A3(\design_top.core0.REG1[11][11] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01126_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16549_ (.A0(\design_top.core0.REG1[12][11] ),
    .A1(\design_top.core0.REG1[13][11] ),
    .A2(\design_top.core0.REG1[14][11] ),
    .A3(\design_top.core0.REG1[15][11] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01127_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16550_ (.A0(_01124_),
    .A1(_01125_),
    .A2(_01126_),
    .A3(_01127_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_01128_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16551_ (.A0(\design_top.core0.REG2[0][12] ),
    .A1(\design_top.core0.REG2[1][12] ),
    .A2(\design_top.core0.REG2[2][12] ),
    .A3(\design_top.core0.REG2[3][12] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01117_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16552_ (.A0(\design_top.core0.REG2[4][12] ),
    .A1(\design_top.core0.REG2[5][12] ),
    .A2(\design_top.core0.REG2[6][12] ),
    .A3(\design_top.core0.REG2[7][12] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01118_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16553_ (.A0(\design_top.core0.REG2[8][12] ),
    .A1(\design_top.core0.REG2[9][12] ),
    .A2(\design_top.core0.REG2[10][12] ),
    .A3(\design_top.core0.REG2[11][12] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01119_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16554_ (.A0(\design_top.core0.REG2[12][12] ),
    .A1(\design_top.core0.REG2[13][12] ),
    .A2(\design_top.core0.REG2[14][12] ),
    .A3(\design_top.core0.REG2[15][12] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01120_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16555_ (.A0(_01117_),
    .A1(_01118_),
    .A2(_01119_),
    .A3(_01120_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_01121_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16556_ (.A0(\design_top.core0.REG1[0][12] ),
    .A1(\design_top.core0.REG1[1][12] ),
    .A2(\design_top.core0.REG1[2][12] ),
    .A3(\design_top.core0.REG1[3][12] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01111_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16557_ (.A0(\design_top.core0.REG1[4][12] ),
    .A1(\design_top.core0.REG1[5][12] ),
    .A2(\design_top.core0.REG1[6][12] ),
    .A3(\design_top.core0.REG1[7][12] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01112_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16558_ (.A0(\design_top.core0.REG1[8][12] ),
    .A1(\design_top.core0.REG1[9][12] ),
    .A2(\design_top.core0.REG1[10][12] ),
    .A3(\design_top.core0.REG1[11][12] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01113_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16559_ (.A0(\design_top.core0.REG1[12][12] ),
    .A1(\design_top.core0.REG1[13][12] ),
    .A2(\design_top.core0.REG1[14][12] ),
    .A3(\design_top.core0.REG1[15][12] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01114_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16560_ (.A0(_01111_),
    .A1(_01112_),
    .A2(_01113_),
    .A3(_01114_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_01115_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16561_ (.A0(\design_top.core0.REG2[0][13] ),
    .A1(\design_top.core0.REG2[1][13] ),
    .A2(\design_top.core0.REG2[2][13] ),
    .A3(\design_top.core0.REG2[3][13] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01103_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16562_ (.A0(\design_top.core0.REG2[4][13] ),
    .A1(\design_top.core0.REG2[5][13] ),
    .A2(\design_top.core0.REG2[6][13] ),
    .A3(\design_top.core0.REG2[7][13] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01104_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16563_ (.A0(\design_top.core0.REG2[8][13] ),
    .A1(\design_top.core0.REG2[9][13] ),
    .A2(\design_top.core0.REG2[10][13] ),
    .A3(\design_top.core0.REG2[11][13] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01105_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16564_ (.A0(\design_top.core0.REG2[12][13] ),
    .A1(\design_top.core0.REG2[13][13] ),
    .A2(\design_top.core0.REG2[14][13] ),
    .A3(\design_top.core0.REG2[15][13] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01106_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16565_ (.A0(_01103_),
    .A1(_01104_),
    .A2(_01105_),
    .A3(_01106_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_01107_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16566_ (.A0(\design_top.core0.REG1[0][13] ),
    .A1(\design_top.core0.REG1[1][13] ),
    .A2(\design_top.core0.REG1[2][13] ),
    .A3(\design_top.core0.REG1[3][13] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01097_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16567_ (.A0(\design_top.core0.REG1[4][13] ),
    .A1(\design_top.core0.REG1[5][13] ),
    .A2(\design_top.core0.REG1[6][13] ),
    .A3(\design_top.core0.REG1[7][13] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01098_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16568_ (.A0(\design_top.core0.REG1[8][13] ),
    .A1(\design_top.core0.REG1[9][13] ),
    .A2(\design_top.core0.REG1[10][13] ),
    .A3(\design_top.core0.REG1[11][13] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01099_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16569_ (.A0(\design_top.core0.REG1[12][13] ),
    .A1(\design_top.core0.REG1[13][13] ),
    .A2(\design_top.core0.REG1[14][13] ),
    .A3(\design_top.core0.REG1[15][13] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01100_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16570_ (.A0(_01097_),
    .A1(_01098_),
    .A2(_01099_),
    .A3(_01100_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_01101_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16571_ (.A0(\design_top.core0.REG2[0][14] ),
    .A1(\design_top.core0.REG2[1][14] ),
    .A2(\design_top.core0.REG2[2][14] ),
    .A3(\design_top.core0.REG2[3][14] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01090_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16572_ (.A0(\design_top.core0.REG2[4][14] ),
    .A1(\design_top.core0.REG2[5][14] ),
    .A2(\design_top.core0.REG2[6][14] ),
    .A3(\design_top.core0.REG2[7][14] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01091_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16573_ (.A0(\design_top.core0.REG2[8][14] ),
    .A1(\design_top.core0.REG2[9][14] ),
    .A2(\design_top.core0.REG2[10][14] ),
    .A3(\design_top.core0.REG2[11][14] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01092_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16574_ (.A0(\design_top.core0.REG2[12][14] ),
    .A1(\design_top.core0.REG2[13][14] ),
    .A2(\design_top.core0.REG2[14][14] ),
    .A3(\design_top.core0.REG2[15][14] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01093_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16575_ (.A0(_01090_),
    .A1(_01091_),
    .A2(_01092_),
    .A3(_01093_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_01094_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16576_ (.A0(\design_top.core0.REG1[0][14] ),
    .A1(\design_top.core0.REG1[1][14] ),
    .A2(\design_top.core0.REG1[2][14] ),
    .A3(\design_top.core0.REG1[3][14] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01084_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16577_ (.A0(\design_top.core0.REG1[4][14] ),
    .A1(\design_top.core0.REG1[5][14] ),
    .A2(\design_top.core0.REG1[6][14] ),
    .A3(\design_top.core0.REG1[7][14] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01085_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16578_ (.A0(\design_top.core0.REG1[8][14] ),
    .A1(\design_top.core0.REG1[9][14] ),
    .A2(\design_top.core0.REG1[10][14] ),
    .A3(\design_top.core0.REG1[11][14] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01086_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16579_ (.A0(\design_top.core0.REG1[12][14] ),
    .A1(\design_top.core0.REG1[13][14] ),
    .A2(\design_top.core0.REG1[14][14] ),
    .A3(\design_top.core0.REG1[15][14] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01087_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16580_ (.A0(_01084_),
    .A1(_01085_),
    .A2(_01086_),
    .A3(_01087_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_01088_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16581_ (.A0(\design_top.core0.REG2[0][15] ),
    .A1(\design_top.core0.REG2[1][15] ),
    .A2(\design_top.core0.REG2[2][15] ),
    .A3(\design_top.core0.REG2[3][15] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01076_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16582_ (.A0(\design_top.core0.REG2[4][15] ),
    .A1(\design_top.core0.REG2[5][15] ),
    .A2(\design_top.core0.REG2[6][15] ),
    .A3(\design_top.core0.REG2[7][15] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01077_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16583_ (.A0(\design_top.core0.REG2[8][15] ),
    .A1(\design_top.core0.REG2[9][15] ),
    .A2(\design_top.core0.REG2[10][15] ),
    .A3(\design_top.core0.REG2[11][15] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01078_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16584_ (.A0(\design_top.core0.REG2[12][15] ),
    .A1(\design_top.core0.REG2[13][15] ),
    .A2(\design_top.core0.REG2[14][15] ),
    .A3(\design_top.core0.REG2[15][15] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01079_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16585_ (.A0(_01076_),
    .A1(_01077_),
    .A2(_01078_),
    .A3(_01079_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_01080_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16586_ (.A0(\design_top.core0.REG1[0][15] ),
    .A1(\design_top.core0.REG1[1][15] ),
    .A2(\design_top.core0.REG1[2][15] ),
    .A3(\design_top.core0.REG1[3][15] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01070_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16587_ (.A0(\design_top.core0.REG1[4][15] ),
    .A1(\design_top.core0.REG1[5][15] ),
    .A2(\design_top.core0.REG1[6][15] ),
    .A3(\design_top.core0.REG1[7][15] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01071_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16588_ (.A0(\design_top.core0.REG1[8][15] ),
    .A1(\design_top.core0.REG1[9][15] ),
    .A2(\design_top.core0.REG1[10][15] ),
    .A3(\design_top.core0.REG1[11][15] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01072_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16589_ (.A0(\design_top.core0.REG1[12][15] ),
    .A1(\design_top.core0.REG1[13][15] ),
    .A2(\design_top.core0.REG1[14][15] ),
    .A3(\design_top.core0.REG1[15][15] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01073_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16590_ (.A0(_01070_),
    .A1(_01071_),
    .A2(_01072_),
    .A3(_01073_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_01074_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16591_ (.A0(\design_top.core0.REG2[0][16] ),
    .A1(\design_top.core0.REG2[1][16] ),
    .A2(\design_top.core0.REG2[2][16] ),
    .A3(\design_top.core0.REG2[3][16] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01063_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16592_ (.A0(\design_top.core0.REG2[4][16] ),
    .A1(\design_top.core0.REG2[5][16] ),
    .A2(\design_top.core0.REG2[6][16] ),
    .A3(\design_top.core0.REG2[7][16] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16593_ (.A0(\design_top.core0.REG2[8][16] ),
    .A1(\design_top.core0.REG2[9][16] ),
    .A2(\design_top.core0.REG2[10][16] ),
    .A3(\design_top.core0.REG2[11][16] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01065_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16594_ (.A0(\design_top.core0.REG2[12][16] ),
    .A1(\design_top.core0.REG2[13][16] ),
    .A2(\design_top.core0.REG2[14][16] ),
    .A3(\design_top.core0.REG2[15][16] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16595_ (.A0(_01063_),
    .A1(_01064_),
    .A2(_01065_),
    .A3(_01066_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_01067_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16596_ (.A0(\design_top.core0.REG1[0][16] ),
    .A1(\design_top.core0.REG1[1][16] ),
    .A2(\design_top.core0.REG1[2][16] ),
    .A3(\design_top.core0.REG1[3][16] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16597_ (.A0(\design_top.core0.REG1[4][16] ),
    .A1(\design_top.core0.REG1[5][16] ),
    .A2(\design_top.core0.REG1[6][16] ),
    .A3(\design_top.core0.REG1[7][16] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16598_ (.A0(\design_top.core0.REG1[8][16] ),
    .A1(\design_top.core0.REG1[9][16] ),
    .A2(\design_top.core0.REG1[10][16] ),
    .A3(\design_top.core0.REG1[11][16] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16599_ (.A0(\design_top.core0.REG1[12][16] ),
    .A1(\design_top.core0.REG1[13][16] ),
    .A2(\design_top.core0.REG1[14][16] ),
    .A3(\design_top.core0.REG1[15][16] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16600_ (.A0(_01057_),
    .A1(_01058_),
    .A2(_01059_),
    .A3(_01060_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_01061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16601_ (.A0(\design_top.core0.REG2[0][17] ),
    .A1(\design_top.core0.REG2[1][17] ),
    .A2(\design_top.core0.REG2[2][17] ),
    .A3(\design_top.core0.REG2[3][17] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16602_ (.A0(\design_top.core0.REG2[4][17] ),
    .A1(\design_top.core0.REG2[5][17] ),
    .A2(\design_top.core0.REG2[6][17] ),
    .A3(\design_top.core0.REG2[7][17] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16603_ (.A0(\design_top.core0.REG2[8][17] ),
    .A1(\design_top.core0.REG2[9][17] ),
    .A2(\design_top.core0.REG2[10][17] ),
    .A3(\design_top.core0.REG2[11][17] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16604_ (.A0(\design_top.core0.REG2[12][17] ),
    .A1(\design_top.core0.REG2[13][17] ),
    .A2(\design_top.core0.REG2[14][17] ),
    .A3(\design_top.core0.REG2[15][17] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16605_ (.A0(_01049_),
    .A1(_01050_),
    .A2(_01051_),
    .A3(_01052_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_01053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16606_ (.A0(_01028_),
    .A1(_01029_),
    .A2(_01030_),
    .A3(_01031_),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16607_ (.A0(_01033_),
    .A1(_01034_),
    .A2(_01035_),
    .A3(_01036_),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16608_ (.A0(_01038_),
    .A1(_01039_),
    .A2(_01040_),
    .A3(_01041_),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16609_ (.A0(_01043_),
    .A1(_01044_),
    .A2(_01045_),
    .A3(_01046_),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16610_ (.A0(_01032_),
    .A1(_01037_),
    .A2(_01042_),
    .A3(_01047_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_01048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16611_ (.A0(\design_top.core0.REG2[0][18] ),
    .A1(\design_top.core0.REG2[1][18] ),
    .A2(\design_top.core0.REG2[2][18] ),
    .A3(\design_top.core0.REG2[3][18] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16612_ (.A0(\design_top.core0.REG2[4][18] ),
    .A1(\design_top.core0.REG2[5][18] ),
    .A2(\design_top.core0.REG2[6][18] ),
    .A3(\design_top.core0.REG2[7][18] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16613_ (.A0(\design_top.core0.REG2[8][18] ),
    .A1(\design_top.core0.REG2[9][18] ),
    .A2(\design_top.core0.REG2[10][18] ),
    .A3(\design_top.core0.REG2[11][18] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16614_ (.A0(\design_top.core0.REG2[12][18] ),
    .A1(\design_top.core0.REG2[13][18] ),
    .A2(\design_top.core0.REG2[14][18] ),
    .A3(\design_top.core0.REG2[15][18] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16615_ (.A0(_01021_),
    .A1(_01022_),
    .A2(_01023_),
    .A3(_01024_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_01025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16616_ (.A0(\design_top.core0.REG1[0][18] ),
    .A1(\design_top.core0.REG1[1][18] ),
    .A2(\design_top.core0.REG1[2][18] ),
    .A3(\design_top.core0.REG1[3][18] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16617_ (.A0(\design_top.core0.REG1[4][18] ),
    .A1(\design_top.core0.REG1[5][18] ),
    .A2(\design_top.core0.REG1[6][18] ),
    .A3(\design_top.core0.REG1[7][18] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16618_ (.A0(\design_top.core0.REG1[8][18] ),
    .A1(\design_top.core0.REG1[9][18] ),
    .A2(\design_top.core0.REG1[10][18] ),
    .A3(\design_top.core0.REG1[11][18] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16619_ (.A0(\design_top.core0.REG1[12][18] ),
    .A1(\design_top.core0.REG1[13][18] ),
    .A2(\design_top.core0.REG1[14][18] ),
    .A3(\design_top.core0.REG1[15][18] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16620_ (.A0(_01015_),
    .A1(_01016_),
    .A2(_01017_),
    .A3(_01018_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_01019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16621_ (.A0(\design_top.core0.REG2[0][19] ),
    .A1(\design_top.core0.REG2[1][19] ),
    .A2(\design_top.core0.REG2[2][19] ),
    .A3(\design_top.core0.REG2[3][19] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16622_ (.A0(\design_top.core0.REG2[4][19] ),
    .A1(\design_top.core0.REG2[5][19] ),
    .A2(\design_top.core0.REG2[6][19] ),
    .A3(\design_top.core0.REG2[7][19] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16623_ (.A0(\design_top.core0.REG2[8][19] ),
    .A1(\design_top.core0.REG2[9][19] ),
    .A2(\design_top.core0.REG2[10][19] ),
    .A3(\design_top.core0.REG2[11][19] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16624_ (.A0(\design_top.core0.REG2[12][19] ),
    .A1(\design_top.core0.REG2[13][19] ),
    .A2(\design_top.core0.REG2[14][19] ),
    .A3(\design_top.core0.REG2[15][19] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_01010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16625_ (.A0(_01007_),
    .A1(_01008_),
    .A2(_01009_),
    .A3(_01010_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_01011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16626_ (.A0(\design_top.core0.REG1[0][19] ),
    .A1(\design_top.core0.REG1[1][19] ),
    .A2(\design_top.core0.REG1[2][19] ),
    .A3(\design_top.core0.REG1[3][19] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16627_ (.A0(\design_top.core0.REG1[4][19] ),
    .A1(\design_top.core0.REG1[5][19] ),
    .A2(\design_top.core0.REG1[6][19] ),
    .A3(\design_top.core0.REG1[7][19] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16628_ (.A0(\design_top.core0.REG1[8][19] ),
    .A1(\design_top.core0.REG1[9][19] ),
    .A2(\design_top.core0.REG1[10][19] ),
    .A3(\design_top.core0.REG1[11][19] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16629_ (.A0(\design_top.core0.REG1[12][19] ),
    .A1(\design_top.core0.REG1[13][19] ),
    .A2(\design_top.core0.REG1[14][19] ),
    .A3(\design_top.core0.REG1[15][19] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_01004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16630_ (.A0(_01001_),
    .A1(_01002_),
    .A2(_01003_),
    .A3(_01004_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_01005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16631_ (.A0(\design_top.core0.REG2[0][20] ),
    .A1(\design_top.core0.REG2[1][20] ),
    .A2(\design_top.core0.REG2[2][20] ),
    .A3(\design_top.core0.REG2[3][20] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16632_ (.A0(\design_top.core0.REG2[4][20] ),
    .A1(\design_top.core0.REG2[5][20] ),
    .A2(\design_top.core0.REG2[6][20] ),
    .A3(\design_top.core0.REG2[7][20] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16633_ (.A0(\design_top.core0.REG2[8][20] ),
    .A1(\design_top.core0.REG2[9][20] ),
    .A2(\design_top.core0.REG2[10][20] ),
    .A3(\design_top.core0.REG2[11][20] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16634_ (.A0(\design_top.core0.REG2[12][20] ),
    .A1(\design_top.core0.REG2[13][20] ),
    .A2(\design_top.core0.REG2[14][20] ),
    .A3(\design_top.core0.REG2[15][20] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16635_ (.A0(_00994_),
    .A1(_00995_),
    .A2(_00996_),
    .A3(_00997_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_00998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16636_ (.A0(\design_top.core0.REG1[0][20] ),
    .A1(\design_top.core0.REG1[1][20] ),
    .A2(\design_top.core0.REG1[2][20] ),
    .A3(\design_top.core0.REG1[3][20] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16637_ (.A0(\design_top.core0.REG1[4][20] ),
    .A1(\design_top.core0.REG1[5][20] ),
    .A2(\design_top.core0.REG1[6][20] ),
    .A3(\design_top.core0.REG1[7][20] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16638_ (.A0(\design_top.core0.REG1[8][20] ),
    .A1(\design_top.core0.REG1[9][20] ),
    .A2(\design_top.core0.REG1[10][20] ),
    .A3(\design_top.core0.REG1[11][20] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16639_ (.A0(\design_top.core0.REG1[12][20] ),
    .A1(\design_top.core0.REG1[13][20] ),
    .A2(\design_top.core0.REG1[14][20] ),
    .A3(\design_top.core0.REG1[15][20] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16640_ (.A0(_00988_),
    .A1(_00989_),
    .A2(_00990_),
    .A3(_00991_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_00992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16641_ (.A0(\design_top.core0.REG2[0][21] ),
    .A1(\design_top.core0.REG2[1][21] ),
    .A2(\design_top.core0.REG2[2][21] ),
    .A3(\design_top.core0.REG2[3][21] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16642_ (.A0(\design_top.core0.REG2[4][21] ),
    .A1(\design_top.core0.REG2[5][21] ),
    .A2(\design_top.core0.REG2[6][21] ),
    .A3(\design_top.core0.REG2[7][21] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16643_ (.A0(\design_top.core0.REG2[8][21] ),
    .A1(\design_top.core0.REG2[9][21] ),
    .A2(\design_top.core0.REG2[10][21] ),
    .A3(\design_top.core0.REG2[11][21] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16644_ (.A0(\design_top.core0.REG2[12][21] ),
    .A1(\design_top.core0.REG2[13][21] ),
    .A2(\design_top.core0.REG2[14][21] ),
    .A3(\design_top.core0.REG2[15][21] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16645_ (.A0(_00980_),
    .A1(_00981_),
    .A2(_00982_),
    .A3(_00983_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_00984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16646_ (.A0(\design_top.core0.REG1[0][21] ),
    .A1(\design_top.core0.REG1[1][21] ),
    .A2(\design_top.core0.REG1[2][21] ),
    .A3(\design_top.core0.REG1[3][21] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16647_ (.A0(\design_top.core0.REG1[4][21] ),
    .A1(\design_top.core0.REG1[5][21] ),
    .A2(\design_top.core0.REG1[6][21] ),
    .A3(\design_top.core0.REG1[7][21] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16648_ (.A0(\design_top.core0.REG1[8][21] ),
    .A1(\design_top.core0.REG1[9][21] ),
    .A2(\design_top.core0.REG1[10][21] ),
    .A3(\design_top.core0.REG1[11][21] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16649_ (.A0(\design_top.core0.REG1[12][21] ),
    .A1(\design_top.core0.REG1[13][21] ),
    .A2(\design_top.core0.REG1[14][21] ),
    .A3(\design_top.core0.REG1[15][21] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16650_ (.A0(_00974_),
    .A1(_00975_),
    .A2(_00976_),
    .A3(_00977_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_00978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16651_ (.A0(\design_top.core0.REG2[0][22] ),
    .A1(\design_top.core0.REG2[1][22] ),
    .A2(\design_top.core0.REG2[2][22] ),
    .A3(\design_top.core0.REG2[3][22] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16652_ (.A0(\design_top.core0.REG2[4][22] ),
    .A1(\design_top.core0.REG2[5][22] ),
    .A2(\design_top.core0.REG2[6][22] ),
    .A3(\design_top.core0.REG2[7][22] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16653_ (.A0(\design_top.core0.REG2[8][22] ),
    .A1(\design_top.core0.REG2[9][22] ),
    .A2(\design_top.core0.REG2[10][22] ),
    .A3(\design_top.core0.REG2[11][22] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16654_ (.A0(\design_top.core0.REG2[12][22] ),
    .A1(\design_top.core0.REG2[13][22] ),
    .A2(\design_top.core0.REG2[14][22] ),
    .A3(\design_top.core0.REG2[15][22] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16655_ (.A0(_00967_),
    .A1(_00968_),
    .A2(_00969_),
    .A3(_00970_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_00971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16656_ (.A0(\design_top.core0.REG1[0][22] ),
    .A1(\design_top.core0.REG1[1][22] ),
    .A2(\design_top.core0.REG1[2][22] ),
    .A3(\design_top.core0.REG1[3][22] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16657_ (.A0(\design_top.core0.REG1[4][22] ),
    .A1(\design_top.core0.REG1[5][22] ),
    .A2(\design_top.core0.REG1[6][22] ),
    .A3(\design_top.core0.REG1[7][22] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16658_ (.A0(\design_top.core0.REG1[8][22] ),
    .A1(\design_top.core0.REG1[9][22] ),
    .A2(\design_top.core0.REG1[10][22] ),
    .A3(\design_top.core0.REG1[11][22] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16659_ (.A0(\design_top.core0.REG1[12][22] ),
    .A1(\design_top.core0.REG1[13][22] ),
    .A2(\design_top.core0.REG1[14][22] ),
    .A3(\design_top.core0.REG1[15][22] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16660_ (.A0(_00961_),
    .A1(_00962_),
    .A2(_00963_),
    .A3(_00964_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_00965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16661_ (.A0(\design_top.core0.REG2[0][23] ),
    .A1(\design_top.core0.REG2[1][23] ),
    .A2(\design_top.core0.REG2[2][23] ),
    .A3(\design_top.core0.REG2[3][23] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16662_ (.A0(\design_top.core0.REG2[4][23] ),
    .A1(\design_top.core0.REG2[5][23] ),
    .A2(\design_top.core0.REG2[6][23] ),
    .A3(\design_top.core0.REG2[7][23] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16663_ (.A0(\design_top.core0.REG2[8][23] ),
    .A1(\design_top.core0.REG2[9][23] ),
    .A2(\design_top.core0.REG2[10][23] ),
    .A3(\design_top.core0.REG2[11][23] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16664_ (.A0(\design_top.core0.REG2[12][23] ),
    .A1(\design_top.core0.REG2[13][23] ),
    .A2(\design_top.core0.REG2[14][23] ),
    .A3(\design_top.core0.REG2[15][23] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16665_ (.A0(_00953_),
    .A1(_00954_),
    .A2(_00955_),
    .A3(_00956_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_00957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16666_ (.A0(\design_top.core0.REG1[0][23] ),
    .A1(\design_top.core0.REG1[1][23] ),
    .A2(\design_top.core0.REG1[2][23] ),
    .A3(\design_top.core0.REG1[3][23] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16667_ (.A0(\design_top.core0.REG1[4][23] ),
    .A1(\design_top.core0.REG1[5][23] ),
    .A2(\design_top.core0.REG1[6][23] ),
    .A3(\design_top.core0.REG1[7][23] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16668_ (.A0(\design_top.core0.REG1[8][23] ),
    .A1(\design_top.core0.REG1[9][23] ),
    .A2(\design_top.core0.REG1[10][23] ),
    .A3(\design_top.core0.REG1[11][23] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16669_ (.A0(\design_top.core0.REG1[12][23] ),
    .A1(\design_top.core0.REG1[13][23] ),
    .A2(\design_top.core0.REG1[14][23] ),
    .A3(\design_top.core0.REG1[15][23] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16670_ (.A0(_00947_),
    .A1(_00948_),
    .A2(_00949_),
    .A3(_00950_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_00951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16671_ (.A0(\design_top.core0.REG2[0][24] ),
    .A1(\design_top.core0.REG2[1][24] ),
    .A2(\design_top.core0.REG2[2][24] ),
    .A3(\design_top.core0.REG2[3][24] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00940_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16672_ (.A0(\design_top.core0.REG2[4][24] ),
    .A1(\design_top.core0.REG2[5][24] ),
    .A2(\design_top.core0.REG2[6][24] ),
    .A3(\design_top.core0.REG2[7][24] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00941_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16673_ (.A0(\design_top.core0.REG2[8][24] ),
    .A1(\design_top.core0.REG2[9][24] ),
    .A2(\design_top.core0.REG2[10][24] ),
    .A3(\design_top.core0.REG2[11][24] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00942_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16674_ (.A0(\design_top.core0.REG2[12][24] ),
    .A1(\design_top.core0.REG2[13][24] ),
    .A2(\design_top.core0.REG2[14][24] ),
    .A3(\design_top.core0.REG2[15][24] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00943_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16675_ (.A0(_00940_),
    .A1(_00941_),
    .A2(_00942_),
    .A3(_00943_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_00944_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16676_ (.A0(\design_top.core0.REG1[0][24] ),
    .A1(\design_top.core0.REG1[1][24] ),
    .A2(\design_top.core0.REG1[2][24] ),
    .A3(\design_top.core0.REG1[3][24] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00934_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16677_ (.A0(\design_top.core0.REG1[4][24] ),
    .A1(\design_top.core0.REG1[5][24] ),
    .A2(\design_top.core0.REG1[6][24] ),
    .A3(\design_top.core0.REG1[7][24] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00935_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16678_ (.A0(\design_top.core0.REG1[8][24] ),
    .A1(\design_top.core0.REG1[9][24] ),
    .A2(\design_top.core0.REG1[10][24] ),
    .A3(\design_top.core0.REG1[11][24] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00936_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16679_ (.A0(\design_top.core0.REG1[12][24] ),
    .A1(\design_top.core0.REG1[13][24] ),
    .A2(\design_top.core0.REG1[14][24] ),
    .A3(\design_top.core0.REG1[15][24] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00937_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16680_ (.A0(_00934_),
    .A1(_00935_),
    .A2(_00936_),
    .A3(_00937_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_00938_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16681_ (.A0(\design_top.core0.REG2[0][25] ),
    .A1(\design_top.core0.REG2[1][25] ),
    .A2(\design_top.core0.REG2[2][25] ),
    .A3(\design_top.core0.REG2[3][25] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00926_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16682_ (.A0(\design_top.core0.REG2[4][25] ),
    .A1(\design_top.core0.REG2[5][25] ),
    .A2(\design_top.core0.REG2[6][25] ),
    .A3(\design_top.core0.REG2[7][25] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00927_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16683_ (.A0(\design_top.core0.REG2[8][25] ),
    .A1(\design_top.core0.REG2[9][25] ),
    .A2(\design_top.core0.REG2[10][25] ),
    .A3(\design_top.core0.REG2[11][25] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00928_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16684_ (.A0(\design_top.core0.REG2[12][25] ),
    .A1(\design_top.core0.REG2[13][25] ),
    .A2(\design_top.core0.REG2[14][25] ),
    .A3(\design_top.core0.REG2[15][25] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00929_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16685_ (.A0(_00926_),
    .A1(_00927_),
    .A2(_00928_),
    .A3(_00929_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_00930_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16686_ (.A0(\design_top.core0.REG1[0][25] ),
    .A1(\design_top.core0.REG1[1][25] ),
    .A2(\design_top.core0.REG1[2][25] ),
    .A3(\design_top.core0.REG1[3][25] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00920_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16687_ (.A0(\design_top.core0.REG1[4][25] ),
    .A1(\design_top.core0.REG1[5][25] ),
    .A2(\design_top.core0.REG1[6][25] ),
    .A3(\design_top.core0.REG1[7][25] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00921_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16688_ (.A0(\design_top.core0.REG1[8][25] ),
    .A1(\design_top.core0.REG1[9][25] ),
    .A2(\design_top.core0.REG1[10][25] ),
    .A3(\design_top.core0.REG1[11][25] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00922_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16689_ (.A0(\design_top.core0.REG1[12][25] ),
    .A1(\design_top.core0.REG1[13][25] ),
    .A2(\design_top.core0.REG1[14][25] ),
    .A3(\design_top.core0.REG1[15][25] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00923_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16690_ (.A0(_00920_),
    .A1(_00921_),
    .A2(_00922_),
    .A3(_00923_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_00924_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16691_ (.A0(\design_top.core0.REG2[0][26] ),
    .A1(\design_top.core0.REG2[1][26] ),
    .A2(\design_top.core0.REG2[2][26] ),
    .A3(\design_top.core0.REG2[3][26] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00913_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16692_ (.A0(\design_top.core0.REG2[4][26] ),
    .A1(\design_top.core0.REG2[5][26] ),
    .A2(\design_top.core0.REG2[6][26] ),
    .A3(\design_top.core0.REG2[7][26] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00914_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16693_ (.A0(\design_top.core0.REG2[8][26] ),
    .A1(\design_top.core0.REG2[9][26] ),
    .A2(\design_top.core0.REG2[10][26] ),
    .A3(\design_top.core0.REG2[11][26] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00915_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16694_ (.A0(\design_top.core0.REG2[12][26] ),
    .A1(\design_top.core0.REG2[13][26] ),
    .A2(\design_top.core0.REG2[14][26] ),
    .A3(\design_top.core0.REG2[15][26] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00916_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16695_ (.A0(_00913_),
    .A1(_00914_),
    .A2(_00915_),
    .A3(_00916_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_00917_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16696_ (.A0(\design_top.core0.REG1[0][26] ),
    .A1(\design_top.core0.REG1[1][26] ),
    .A2(\design_top.core0.REG1[2][26] ),
    .A3(\design_top.core0.REG1[3][26] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16697_ (.A0(\design_top.core0.REG1[4][26] ),
    .A1(\design_top.core0.REG1[5][26] ),
    .A2(\design_top.core0.REG1[6][26] ),
    .A3(\design_top.core0.REG1[7][26] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16698_ (.A0(\design_top.core0.REG1[8][26] ),
    .A1(\design_top.core0.REG1[9][26] ),
    .A2(\design_top.core0.REG1[10][26] ),
    .A3(\design_top.core0.REG1[11][26] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16699_ (.A0(\design_top.core0.REG1[12][26] ),
    .A1(\design_top.core0.REG1[13][26] ),
    .A2(\design_top.core0.REG1[14][26] ),
    .A3(\design_top.core0.REG1[15][26] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16700_ (.A0(_00907_),
    .A1(_00908_),
    .A2(_00909_),
    .A3(_00910_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_00911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16701_ (.A0(\design_top.core0.REG2[0][27] ),
    .A1(\design_top.core0.REG2[1][27] ),
    .A2(\design_top.core0.REG2[2][27] ),
    .A3(\design_top.core0.REG2[3][27] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16702_ (.A0(\design_top.core0.REG2[4][27] ),
    .A1(\design_top.core0.REG2[5][27] ),
    .A2(\design_top.core0.REG2[6][27] ),
    .A3(\design_top.core0.REG2[7][27] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16703_ (.A0(\design_top.core0.REG2[8][27] ),
    .A1(\design_top.core0.REG2[9][27] ),
    .A2(\design_top.core0.REG2[10][27] ),
    .A3(\design_top.core0.REG2[11][27] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16704_ (.A0(\design_top.core0.REG2[12][27] ),
    .A1(\design_top.core0.REG2[13][27] ),
    .A2(\design_top.core0.REG2[14][27] ),
    .A3(\design_top.core0.REG2[15][27] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16705_ (.A0(_00899_),
    .A1(_00900_),
    .A2(_00901_),
    .A3(_00902_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_00903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16706_ (.A0(\design_top.core0.REG1[0][27] ),
    .A1(\design_top.core0.REG1[1][27] ),
    .A2(\design_top.core0.REG1[2][27] ),
    .A3(\design_top.core0.REG1[3][27] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16707_ (.A0(\design_top.core0.REG1[4][27] ),
    .A1(\design_top.core0.REG1[5][27] ),
    .A2(\design_top.core0.REG1[6][27] ),
    .A3(\design_top.core0.REG1[7][27] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16708_ (.A0(\design_top.core0.REG1[8][27] ),
    .A1(\design_top.core0.REG1[9][27] ),
    .A2(\design_top.core0.REG1[10][27] ),
    .A3(\design_top.core0.REG1[11][27] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16709_ (.A0(\design_top.core0.REG1[12][27] ),
    .A1(\design_top.core0.REG1[13][27] ),
    .A2(\design_top.core0.REG1[14][27] ),
    .A3(\design_top.core0.REG1[15][27] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16710_ (.A0(_00893_),
    .A1(_00894_),
    .A2(_00895_),
    .A3(_00896_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_00897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16711_ (.A0(\design_top.core0.REG2[0][28] ),
    .A1(\design_top.core0.REG2[1][28] ),
    .A2(\design_top.core0.REG2[2][28] ),
    .A3(\design_top.core0.REG2[3][28] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16712_ (.A0(\design_top.core0.REG2[4][28] ),
    .A1(\design_top.core0.REG2[5][28] ),
    .A2(\design_top.core0.REG2[6][28] ),
    .A3(\design_top.core0.REG2[7][28] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16713_ (.A0(\design_top.core0.REG2[8][28] ),
    .A1(\design_top.core0.REG2[9][28] ),
    .A2(\design_top.core0.REG2[10][28] ),
    .A3(\design_top.core0.REG2[11][28] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16714_ (.A0(\design_top.core0.REG2[12][28] ),
    .A1(\design_top.core0.REG2[13][28] ),
    .A2(\design_top.core0.REG2[14][28] ),
    .A3(\design_top.core0.REG2[15][28] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16715_ (.A0(_00886_),
    .A1(_00887_),
    .A2(_00888_),
    .A3(_00889_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_00890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16716_ (.A0(\design_top.core0.REG1[0][28] ),
    .A1(\design_top.core0.REG1[1][28] ),
    .A2(\design_top.core0.REG1[2][28] ),
    .A3(\design_top.core0.REG1[3][28] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16717_ (.A0(\design_top.core0.REG1[4][28] ),
    .A1(\design_top.core0.REG1[5][28] ),
    .A2(\design_top.core0.REG1[6][28] ),
    .A3(\design_top.core0.REG1[7][28] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16718_ (.A0(\design_top.core0.REG1[8][28] ),
    .A1(\design_top.core0.REG1[9][28] ),
    .A2(\design_top.core0.REG1[10][28] ),
    .A3(\design_top.core0.REG1[11][28] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16719_ (.A0(\design_top.core0.REG1[12][28] ),
    .A1(\design_top.core0.REG1[13][28] ),
    .A2(\design_top.core0.REG1[14][28] ),
    .A3(\design_top.core0.REG1[15][28] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16720_ (.A0(_00880_),
    .A1(_00881_),
    .A2(_00882_),
    .A3(_00883_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_00884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16721_ (.A0(\design_top.core0.REG2[0][29] ),
    .A1(\design_top.core0.REG2[1][29] ),
    .A2(\design_top.core0.REG2[2][29] ),
    .A3(\design_top.core0.REG2[3][29] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16722_ (.A0(\design_top.core0.REG2[4][29] ),
    .A1(\design_top.core0.REG2[5][29] ),
    .A2(\design_top.core0.REG2[6][29] ),
    .A3(\design_top.core0.REG2[7][29] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16723_ (.A0(\design_top.core0.REG2[8][29] ),
    .A1(\design_top.core0.REG2[9][29] ),
    .A2(\design_top.core0.REG2[10][29] ),
    .A3(\design_top.core0.REG2[11][29] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16724_ (.A0(\design_top.core0.REG2[12][29] ),
    .A1(\design_top.core0.REG2[13][29] ),
    .A2(\design_top.core0.REG2[14][29] ),
    .A3(\design_top.core0.REG2[15][29] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16725_ (.A0(_00872_),
    .A1(_00873_),
    .A2(_00874_),
    .A3(_00875_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_00876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16726_ (.A0(\design_top.core0.REG1[0][29] ),
    .A1(\design_top.core0.REG1[1][29] ),
    .A2(\design_top.core0.REG1[2][29] ),
    .A3(\design_top.core0.REG1[3][29] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16727_ (.A0(\design_top.core0.REG1[4][29] ),
    .A1(\design_top.core0.REG1[5][29] ),
    .A2(\design_top.core0.REG1[6][29] ),
    .A3(\design_top.core0.REG1[7][29] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16728_ (.A0(\design_top.core0.REG1[8][29] ),
    .A1(\design_top.core0.REG1[9][29] ),
    .A2(\design_top.core0.REG1[10][29] ),
    .A3(\design_top.core0.REG1[11][29] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16729_ (.A0(\design_top.core0.REG1[12][29] ),
    .A1(\design_top.core0.REG1[13][29] ),
    .A2(\design_top.core0.REG1[14][29] ),
    .A3(\design_top.core0.REG1[15][29] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16730_ (.A0(_00866_),
    .A1(_00867_),
    .A2(_00868_),
    .A3(_00869_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_00870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16731_ (.A0(\design_top.core0.REG2[0][30] ),
    .A1(\design_top.core0.REG2[1][30] ),
    .A2(\design_top.core0.REG2[2][30] ),
    .A3(\design_top.core0.REG2[3][30] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16732_ (.A0(\design_top.core0.REG2[4][30] ),
    .A1(\design_top.core0.REG2[5][30] ),
    .A2(\design_top.core0.REG2[6][30] ),
    .A3(\design_top.core0.REG2[7][30] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16733_ (.A0(\design_top.core0.REG2[8][30] ),
    .A1(\design_top.core0.REG2[9][30] ),
    .A2(\design_top.core0.REG2[10][30] ),
    .A3(\design_top.core0.REG2[11][30] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16734_ (.A0(\design_top.core0.REG2[12][30] ),
    .A1(\design_top.core0.REG2[13][30] ),
    .A2(\design_top.core0.REG2[14][30] ),
    .A3(\design_top.core0.REG2[15][30] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16735_ (.A0(_00858_),
    .A1(_00859_),
    .A2(_00860_),
    .A3(_00861_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_00862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16736_ (.A0(\design_top.core0.REG1[0][30] ),
    .A1(\design_top.core0.REG1[1][30] ),
    .A2(\design_top.core0.REG1[2][30] ),
    .A3(\design_top.core0.REG1[3][30] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16737_ (.A0(\design_top.core0.REG1[4][30] ),
    .A1(\design_top.core0.REG1[5][30] ),
    .A2(\design_top.core0.REG1[6][30] ),
    .A3(\design_top.core0.REG1[7][30] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16738_ (.A0(\design_top.core0.REG1[8][30] ),
    .A1(\design_top.core0.REG1[9][30] ),
    .A2(\design_top.core0.REG1[10][30] ),
    .A3(\design_top.core0.REG1[11][30] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16739_ (.A0(\design_top.core0.REG1[12][30] ),
    .A1(\design_top.core0.REG1[13][30] ),
    .A2(\design_top.core0.REG1[14][30] ),
    .A3(\design_top.core0.REG1[15][30] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16740_ (.A0(_00852_),
    .A1(_00853_),
    .A2(_00854_),
    .A3(_00855_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_00856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16741_ (.A0(\design_top.core0.REG2[0][31] ),
    .A1(\design_top.core0.REG2[1][31] ),
    .A2(\design_top.core0.REG2[2][31] ),
    .A3(\design_top.core0.REG2[3][31] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16742_ (.A0(\design_top.core0.REG2[4][31] ),
    .A1(\design_top.core0.REG2[5][31] ),
    .A2(\design_top.core0.REG2[6][31] ),
    .A3(\design_top.core0.REG2[7][31] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16743_ (.A0(\design_top.core0.REG2[8][31] ),
    .A1(\design_top.core0.REG2[9][31] ),
    .A2(\design_top.core0.REG2[10][31] ),
    .A3(\design_top.core0.REG2[11][31] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16744_ (.A0(\design_top.core0.REG2[12][31] ),
    .A1(\design_top.core0.REG2[13][31] ),
    .A2(\design_top.core0.REG2[14][31] ),
    .A3(\design_top.core0.REG2[15][31] ),
    .S0(_00433_),
    .S1(_00434_),
    .X(_00847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16745_ (.A0(_00844_),
    .A1(_00845_),
    .A2(_00846_),
    .A3(_00847_),
    .S0(_00435_),
    .S1(_00436_),
    .X(_00848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16746_ (.A0(_00823_),
    .A1(_00824_),
    .A2(_00825_),
    .A3(_00826_),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16747_ (.A0(_00828_),
    .A1(_00829_),
    .A2(_00830_),
    .A3(_00831_),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16748_ (.A0(_00833_),
    .A1(_00834_),
    .A2(_00835_),
    .A3(_00836_),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16749_ (.A0(_00838_),
    .A1(_00839_),
    .A2(_00840_),
    .A3(_00841_),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16750_ (.A0(_00827_),
    .A1(_00832_),
    .A2(_00837_),
    .A3(_00842_),
    .S0(_00431_),
    .S1(_00432_),
    .X(_00843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16751_ (.A0(\design_top.core0.REG1[8][3] ),
    .A1(\design_top.core0.REG1[9][3] ),
    .A2(\design_top.core0.REG1[10][3] ),
    .A3(\design_top.core0.REG1[11][3] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16752_ (.A0(\design_top.core0.REG1[12][3] ),
    .A1(\design_top.core0.REG1[13][3] ),
    .A2(\design_top.core0.REG1[14][3] ),
    .A3(\design_top.core0.REG1[15][3] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16753_ (.A0(\design_top.core0.REG1[0][3] ),
    .A1(\design_top.core0.REG1[1][3] ),
    .A2(\design_top.core0.REG1[2][3] ),
    .A3(\design_top.core0.REG1[3][3] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16754_ (.A0(\design_top.core0.REG1[4][3] ),
    .A1(\design_top.core0.REG1[5][3] ),
    .A2(\design_top.core0.REG1[6][3] ),
    .A3(\design_top.core0.REG1[7][3] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16755_ (.A0(\design_top.core0.REG1[8][0] ),
    .A1(\design_top.core0.REG1[9][0] ),
    .A2(\design_top.core0.REG1[10][0] ),
    .A3(\design_top.core0.REG1[11][0] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16756_ (.A0(\design_top.core0.REG1[12][0] ),
    .A1(\design_top.core0.REG1[13][0] ),
    .A2(\design_top.core0.REG1[14][0] ),
    .A3(\design_top.core0.REG1[15][0] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16757_ (.A0(\design_top.core0.REG1[0][0] ),
    .A1(\design_top.core0.REG1[1][0] ),
    .A2(\design_top.core0.REG1[2][0] ),
    .A3(\design_top.core0.REG1[3][0] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16758_ (.A0(\design_top.core0.REG1[4][0] ),
    .A1(\design_top.core0.REG1[5][0] ),
    .A2(\design_top.core0.REG1[6][0] ),
    .A3(\design_top.core0.REG1[7][0] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16759_ (.A0(\design_top.core0.REG1[8][1] ),
    .A1(\design_top.core0.REG1[9][1] ),
    .A2(\design_top.core0.REG1[10][1] ),
    .A3(\design_top.core0.REG1[11][1] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16760_ (.A0(\design_top.core0.REG1[12][1] ),
    .A1(\design_top.core0.REG1[13][1] ),
    .A2(\design_top.core0.REG1[14][1] ),
    .A3(\design_top.core0.REG1[15][1] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16761_ (.A0(\design_top.core0.REG1[0][1] ),
    .A1(\design_top.core0.REG1[1][1] ),
    .A2(\design_top.core0.REG1[2][1] ),
    .A3(\design_top.core0.REG1[3][1] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16762_ (.A0(\design_top.core0.REG1[4][1] ),
    .A1(\design_top.core0.REG1[5][1] ),
    .A2(\design_top.core0.REG1[6][1] ),
    .A3(\design_top.core0.REG1[7][1] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16763_ (.A0(\design_top.core0.REG1[8][2] ),
    .A1(\design_top.core0.REG1[9][2] ),
    .A2(\design_top.core0.REG1[10][2] ),
    .A3(\design_top.core0.REG1[11][2] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16764_ (.A0(\design_top.core0.REG1[12][2] ),
    .A1(\design_top.core0.REG1[13][2] ),
    .A2(\design_top.core0.REG1[14][2] ),
    .A3(\design_top.core0.REG1[15][2] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16765_ (.A0(\design_top.core0.REG1[0][2] ),
    .A1(\design_top.core0.REG1[1][2] ),
    .A2(\design_top.core0.REG1[2][2] ),
    .A3(\design_top.core0.REG1[3][2] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16766_ (.A0(\design_top.core0.REG1[4][2] ),
    .A1(\design_top.core0.REG1[5][2] ),
    .A2(\design_top.core0.REG1[6][2] ),
    .A3(\design_top.core0.REG1[7][2] ),
    .S0(_00429_),
    .S1(_00430_),
    .X(_00788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16767_ (.A0(\design_top.MEM[0][31] ),
    .A1(\design_top.MEM[1][31] ),
    .A2(\design_top.MEM[2][31] ),
    .A3(\design_top.MEM[3][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16768_ (.A0(\design_top.MEM[4][31] ),
    .A1(\design_top.MEM[5][31] ),
    .A2(\design_top.MEM[6][31] ),
    .A3(\design_top.MEM[7][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16769_ (.A0(\design_top.MEM[8][31] ),
    .A1(\design_top.MEM[9][31] ),
    .A2(\design_top.MEM[10][31] ),
    .A3(\design_top.MEM[11][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16770_ (.A0(\design_top.MEM[12][31] ),
    .A1(\design_top.MEM[13][31] ),
    .A2(\design_top.MEM[14][31] ),
    .A3(\design_top.MEM[15][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16771_ (.A0(_00633_),
    .A1(_00634_),
    .A2(_00635_),
    .A3(_00636_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16772_ (.A0(\design_top.MEM[16][31] ),
    .A1(\design_top.MEM[17][31] ),
    .A2(\design_top.MEM[18][31] ),
    .A3(\design_top.MEM[19][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16773_ (.A0(\design_top.MEM[20][31] ),
    .A1(\design_top.MEM[21][31] ),
    .A2(\design_top.MEM[22][31] ),
    .A3(\design_top.MEM[23][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16774_ (.A0(\design_top.MEM[24][31] ),
    .A1(\design_top.MEM[25][31] ),
    .A2(\design_top.MEM[26][31] ),
    .A3(\design_top.MEM[27][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16775_ (.A0(\design_top.MEM[28][31] ),
    .A1(\design_top.MEM[29][31] ),
    .A2(\design_top.MEM[30][31] ),
    .A3(\design_top.MEM[31][31] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16776_ (.A0(_00638_),
    .A1(_00639_),
    .A2(_00640_),
    .A3(_00641_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16777_ (.A0(\design_top.MEM[0][30] ),
    .A1(\design_top.MEM[1][30] ),
    .A2(\design_top.MEM[2][30] ),
    .A3(\design_top.MEM[3][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16778_ (.A0(\design_top.MEM[4][30] ),
    .A1(\design_top.MEM[5][30] ),
    .A2(\design_top.MEM[6][30] ),
    .A3(\design_top.MEM[7][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16779_ (.A0(\design_top.MEM[8][30] ),
    .A1(\design_top.MEM[9][30] ),
    .A2(\design_top.MEM[10][30] ),
    .A3(\design_top.MEM[11][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16780_ (.A0(\design_top.MEM[12][30] ),
    .A1(\design_top.MEM[13][30] ),
    .A2(\design_top.MEM[14][30] ),
    .A3(\design_top.MEM[15][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16781_ (.A0(_00623_),
    .A1(_00624_),
    .A2(_00625_),
    .A3(_00626_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16782_ (.A0(\design_top.MEM[16][30] ),
    .A1(\design_top.MEM[17][30] ),
    .A2(\design_top.MEM[18][30] ),
    .A3(\design_top.MEM[19][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16783_ (.A0(\design_top.MEM[20][30] ),
    .A1(\design_top.MEM[21][30] ),
    .A2(\design_top.MEM[22][30] ),
    .A3(\design_top.MEM[23][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16784_ (.A0(\design_top.MEM[24][30] ),
    .A1(\design_top.MEM[25][30] ),
    .A2(\design_top.MEM[26][30] ),
    .A3(\design_top.MEM[27][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16785_ (.A0(\design_top.MEM[28][30] ),
    .A1(\design_top.MEM[29][30] ),
    .A2(\design_top.MEM[30][30] ),
    .A3(\design_top.MEM[31][30] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16786_ (.A0(_00628_),
    .A1(_00629_),
    .A2(_00630_),
    .A3(_00631_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16787_ (.A0(\design_top.MEM[0][29] ),
    .A1(\design_top.MEM[1][29] ),
    .A2(\design_top.MEM[2][29] ),
    .A3(\design_top.MEM[3][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16788_ (.A0(\design_top.MEM[4][29] ),
    .A1(\design_top.MEM[5][29] ),
    .A2(\design_top.MEM[6][29] ),
    .A3(\design_top.MEM[7][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16789_ (.A0(\design_top.MEM[8][29] ),
    .A1(\design_top.MEM[9][29] ),
    .A2(\design_top.MEM[10][29] ),
    .A3(\design_top.MEM[11][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16790_ (.A0(\design_top.MEM[12][29] ),
    .A1(\design_top.MEM[13][29] ),
    .A2(\design_top.MEM[14][29] ),
    .A3(\design_top.MEM[15][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16791_ (.A0(_00613_),
    .A1(_00614_),
    .A2(_00615_),
    .A3(_00616_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16792_ (.A0(\design_top.MEM[16][29] ),
    .A1(\design_top.MEM[17][29] ),
    .A2(\design_top.MEM[18][29] ),
    .A3(\design_top.MEM[19][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16793_ (.A0(\design_top.MEM[20][29] ),
    .A1(\design_top.MEM[21][29] ),
    .A2(\design_top.MEM[22][29] ),
    .A3(\design_top.MEM[23][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16794_ (.A0(\design_top.MEM[24][29] ),
    .A1(\design_top.MEM[25][29] ),
    .A2(\design_top.MEM[26][29] ),
    .A3(\design_top.MEM[27][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16795_ (.A0(\design_top.MEM[28][29] ),
    .A1(\design_top.MEM[29][29] ),
    .A2(\design_top.MEM[30][29] ),
    .A3(\design_top.MEM[31][29] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16796_ (.A0(_00618_),
    .A1(_00619_),
    .A2(_00620_),
    .A3(_00621_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16797_ (.A0(\design_top.MEM[0][28] ),
    .A1(\design_top.MEM[1][28] ),
    .A2(\design_top.MEM[2][28] ),
    .A3(\design_top.MEM[3][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16798_ (.A0(\design_top.MEM[4][28] ),
    .A1(\design_top.MEM[5][28] ),
    .A2(\design_top.MEM[6][28] ),
    .A3(\design_top.MEM[7][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16799_ (.A0(\design_top.MEM[8][28] ),
    .A1(\design_top.MEM[9][28] ),
    .A2(\design_top.MEM[10][28] ),
    .A3(\design_top.MEM[11][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16800_ (.A0(\design_top.MEM[12][28] ),
    .A1(\design_top.MEM[13][28] ),
    .A2(\design_top.MEM[14][28] ),
    .A3(\design_top.MEM[15][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16801_ (.A0(_00603_),
    .A1(_00604_),
    .A2(_00605_),
    .A3(_00606_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16802_ (.A0(\design_top.MEM[16][28] ),
    .A1(\design_top.MEM[17][28] ),
    .A2(\design_top.MEM[18][28] ),
    .A3(\design_top.MEM[19][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16803_ (.A0(\design_top.MEM[20][28] ),
    .A1(\design_top.MEM[21][28] ),
    .A2(\design_top.MEM[22][28] ),
    .A3(\design_top.MEM[23][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16804_ (.A0(\design_top.MEM[24][28] ),
    .A1(\design_top.MEM[25][28] ),
    .A2(\design_top.MEM[26][28] ),
    .A3(\design_top.MEM[27][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16805_ (.A0(\design_top.MEM[28][28] ),
    .A1(\design_top.MEM[29][28] ),
    .A2(\design_top.MEM[30][28] ),
    .A3(\design_top.MEM[31][28] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16806_ (.A0(_00608_),
    .A1(_00609_),
    .A2(_00610_),
    .A3(_00611_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16807_ (.A0(\design_top.MEM[0][27] ),
    .A1(\design_top.MEM[1][27] ),
    .A2(\design_top.MEM[2][27] ),
    .A3(\design_top.MEM[3][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16808_ (.A0(\design_top.MEM[4][27] ),
    .A1(\design_top.MEM[5][27] ),
    .A2(\design_top.MEM[6][27] ),
    .A3(\design_top.MEM[7][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16809_ (.A0(\design_top.MEM[8][27] ),
    .A1(\design_top.MEM[9][27] ),
    .A2(\design_top.MEM[10][27] ),
    .A3(\design_top.MEM[11][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16810_ (.A0(\design_top.MEM[12][27] ),
    .A1(\design_top.MEM[13][27] ),
    .A2(\design_top.MEM[14][27] ),
    .A3(\design_top.MEM[15][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16811_ (.A0(_00593_),
    .A1(_00594_),
    .A2(_00595_),
    .A3(_00596_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16812_ (.A0(\design_top.MEM[16][27] ),
    .A1(\design_top.MEM[17][27] ),
    .A2(\design_top.MEM[18][27] ),
    .A3(\design_top.MEM[19][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16813_ (.A0(\design_top.MEM[20][27] ),
    .A1(\design_top.MEM[21][27] ),
    .A2(\design_top.MEM[22][27] ),
    .A3(\design_top.MEM[23][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16814_ (.A0(\design_top.MEM[24][27] ),
    .A1(\design_top.MEM[25][27] ),
    .A2(\design_top.MEM[26][27] ),
    .A3(\design_top.MEM[27][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16815_ (.A0(\design_top.MEM[28][27] ),
    .A1(\design_top.MEM[29][27] ),
    .A2(\design_top.MEM[30][27] ),
    .A3(\design_top.MEM[31][27] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16816_ (.A0(_00598_),
    .A1(_00599_),
    .A2(_00600_),
    .A3(_00601_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16817_ (.A0(\design_top.MEM[0][26] ),
    .A1(\design_top.MEM[1][26] ),
    .A2(\design_top.MEM[2][26] ),
    .A3(\design_top.MEM[3][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00583_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16818_ (.A0(\design_top.MEM[4][26] ),
    .A1(\design_top.MEM[5][26] ),
    .A2(\design_top.MEM[6][26] ),
    .A3(\design_top.MEM[7][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00584_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16819_ (.A0(\design_top.MEM[8][26] ),
    .A1(\design_top.MEM[9][26] ),
    .A2(\design_top.MEM[10][26] ),
    .A3(\design_top.MEM[11][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00585_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16820_ (.A0(\design_top.MEM[12][26] ),
    .A1(\design_top.MEM[13][26] ),
    .A2(\design_top.MEM[14][26] ),
    .A3(\design_top.MEM[15][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00586_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16821_ (.A0(_00583_),
    .A1(_00584_),
    .A2(_00585_),
    .A3(_00586_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00587_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16822_ (.A0(\design_top.MEM[16][26] ),
    .A1(\design_top.MEM[17][26] ),
    .A2(\design_top.MEM[18][26] ),
    .A3(\design_top.MEM[19][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00588_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16823_ (.A0(\design_top.MEM[20][26] ),
    .A1(\design_top.MEM[21][26] ),
    .A2(\design_top.MEM[22][26] ),
    .A3(\design_top.MEM[23][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00589_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16824_ (.A0(\design_top.MEM[24][26] ),
    .A1(\design_top.MEM[25][26] ),
    .A2(\design_top.MEM[26][26] ),
    .A3(\design_top.MEM[27][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00590_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16825_ (.A0(\design_top.MEM[28][26] ),
    .A1(\design_top.MEM[29][26] ),
    .A2(\design_top.MEM[30][26] ),
    .A3(\design_top.MEM[31][26] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00591_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16826_ (.A0(_00588_),
    .A1(_00589_),
    .A2(_00590_),
    .A3(_00591_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16827_ (.A0(\design_top.MEM[0][25] ),
    .A1(\design_top.MEM[1][25] ),
    .A2(\design_top.MEM[2][25] ),
    .A3(\design_top.MEM[3][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00573_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16828_ (.A0(\design_top.MEM[4][25] ),
    .A1(\design_top.MEM[5][25] ),
    .A2(\design_top.MEM[6][25] ),
    .A3(\design_top.MEM[7][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00574_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16829_ (.A0(\design_top.MEM[8][25] ),
    .A1(\design_top.MEM[9][25] ),
    .A2(\design_top.MEM[10][25] ),
    .A3(\design_top.MEM[11][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00575_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16830_ (.A0(\design_top.MEM[12][25] ),
    .A1(\design_top.MEM[13][25] ),
    .A2(\design_top.MEM[14][25] ),
    .A3(\design_top.MEM[15][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00576_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16831_ (.A0(_00573_),
    .A1(_00574_),
    .A2(_00575_),
    .A3(_00576_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00577_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16832_ (.A0(\design_top.MEM[16][25] ),
    .A1(\design_top.MEM[17][25] ),
    .A2(\design_top.MEM[18][25] ),
    .A3(\design_top.MEM[19][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00578_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16833_ (.A0(\design_top.MEM[20][25] ),
    .A1(\design_top.MEM[21][25] ),
    .A2(\design_top.MEM[22][25] ),
    .A3(\design_top.MEM[23][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00579_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16834_ (.A0(\design_top.MEM[24][25] ),
    .A1(\design_top.MEM[25][25] ),
    .A2(\design_top.MEM[26][25] ),
    .A3(\design_top.MEM[27][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00580_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16835_ (.A0(\design_top.MEM[28][25] ),
    .A1(\design_top.MEM[29][25] ),
    .A2(\design_top.MEM[30][25] ),
    .A3(\design_top.MEM[31][25] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00581_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16836_ (.A0(_00578_),
    .A1(_00579_),
    .A2(_00580_),
    .A3(_00581_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00582_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16837_ (.A0(\design_top.MEM[0][24] ),
    .A1(\design_top.MEM[1][24] ),
    .A2(\design_top.MEM[2][24] ),
    .A3(\design_top.MEM[3][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00563_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16838_ (.A0(\design_top.MEM[4][24] ),
    .A1(\design_top.MEM[5][24] ),
    .A2(\design_top.MEM[6][24] ),
    .A3(\design_top.MEM[7][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00564_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16839_ (.A0(\design_top.MEM[8][24] ),
    .A1(\design_top.MEM[9][24] ),
    .A2(\design_top.MEM[10][24] ),
    .A3(\design_top.MEM[11][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00565_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16840_ (.A0(\design_top.MEM[12][24] ),
    .A1(\design_top.MEM[13][24] ),
    .A2(\design_top.MEM[14][24] ),
    .A3(\design_top.MEM[15][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00566_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16841_ (.A0(_00563_),
    .A1(_00564_),
    .A2(_00565_),
    .A3(_00566_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00567_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16842_ (.A0(\design_top.MEM[16][24] ),
    .A1(\design_top.MEM[17][24] ),
    .A2(\design_top.MEM[18][24] ),
    .A3(\design_top.MEM[19][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00568_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16843_ (.A0(\design_top.MEM[20][24] ),
    .A1(\design_top.MEM[21][24] ),
    .A2(\design_top.MEM[22][24] ),
    .A3(\design_top.MEM[23][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00569_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16844_ (.A0(\design_top.MEM[24][24] ),
    .A1(\design_top.MEM[25][24] ),
    .A2(\design_top.MEM[26][24] ),
    .A3(\design_top.MEM[27][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00570_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16845_ (.A0(\design_top.MEM[28][24] ),
    .A1(\design_top.MEM[29][24] ),
    .A2(\design_top.MEM[30][24] ),
    .A3(\design_top.MEM[31][24] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00571_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16846_ (.A0(_00568_),
    .A1(_00569_),
    .A2(_00570_),
    .A3(_00571_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00572_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16847_ (.A0(\design_top.MEM[0][23] ),
    .A1(\design_top.MEM[1][23] ),
    .A2(\design_top.MEM[2][23] ),
    .A3(\design_top.MEM[3][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00553_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16848_ (.A0(\design_top.MEM[4][23] ),
    .A1(\design_top.MEM[5][23] ),
    .A2(\design_top.MEM[6][23] ),
    .A3(\design_top.MEM[7][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00554_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16849_ (.A0(\design_top.MEM[8][23] ),
    .A1(\design_top.MEM[9][23] ),
    .A2(\design_top.MEM[10][23] ),
    .A3(\design_top.MEM[11][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00555_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16850_ (.A0(\design_top.MEM[12][23] ),
    .A1(\design_top.MEM[13][23] ),
    .A2(\design_top.MEM[14][23] ),
    .A3(\design_top.MEM[15][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00556_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16851_ (.A0(_00553_),
    .A1(_00554_),
    .A2(_00555_),
    .A3(_00556_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00557_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16852_ (.A0(\design_top.MEM[16][23] ),
    .A1(\design_top.MEM[17][23] ),
    .A2(\design_top.MEM[18][23] ),
    .A3(\design_top.MEM[19][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00558_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16853_ (.A0(\design_top.MEM[20][23] ),
    .A1(\design_top.MEM[21][23] ),
    .A2(\design_top.MEM[22][23] ),
    .A3(\design_top.MEM[23][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00559_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16854_ (.A0(\design_top.MEM[24][23] ),
    .A1(\design_top.MEM[25][23] ),
    .A2(\design_top.MEM[26][23] ),
    .A3(\design_top.MEM[27][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00560_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16855_ (.A0(\design_top.MEM[28][23] ),
    .A1(\design_top.MEM[29][23] ),
    .A2(\design_top.MEM[30][23] ),
    .A3(\design_top.MEM[31][23] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00561_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16856_ (.A0(_00558_),
    .A1(_00559_),
    .A2(_00560_),
    .A3(_00561_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00562_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16857_ (.A0(\design_top.MEM[0][22] ),
    .A1(\design_top.MEM[1][22] ),
    .A2(\design_top.MEM[2][22] ),
    .A3(\design_top.MEM[3][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00543_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16858_ (.A0(\design_top.MEM[4][22] ),
    .A1(\design_top.MEM[5][22] ),
    .A2(\design_top.MEM[6][22] ),
    .A3(\design_top.MEM[7][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00544_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16859_ (.A0(\design_top.MEM[8][22] ),
    .A1(\design_top.MEM[9][22] ),
    .A2(\design_top.MEM[10][22] ),
    .A3(\design_top.MEM[11][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00545_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16860_ (.A0(\design_top.MEM[12][22] ),
    .A1(\design_top.MEM[13][22] ),
    .A2(\design_top.MEM[14][22] ),
    .A3(\design_top.MEM[15][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00546_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16861_ (.A0(_00543_),
    .A1(_00544_),
    .A2(_00545_),
    .A3(_00546_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00547_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16862_ (.A0(\design_top.MEM[16][22] ),
    .A1(\design_top.MEM[17][22] ),
    .A2(\design_top.MEM[18][22] ),
    .A3(\design_top.MEM[19][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00548_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16863_ (.A0(\design_top.MEM[20][22] ),
    .A1(\design_top.MEM[21][22] ),
    .A2(\design_top.MEM[22][22] ),
    .A3(\design_top.MEM[23][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00549_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16864_ (.A0(\design_top.MEM[24][22] ),
    .A1(\design_top.MEM[25][22] ),
    .A2(\design_top.MEM[26][22] ),
    .A3(\design_top.MEM[27][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00550_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16865_ (.A0(\design_top.MEM[28][22] ),
    .A1(\design_top.MEM[29][22] ),
    .A2(\design_top.MEM[30][22] ),
    .A3(\design_top.MEM[31][22] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00551_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16866_ (.A0(_00548_),
    .A1(_00549_),
    .A2(_00550_),
    .A3(_00551_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00552_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16867_ (.A0(\design_top.MEM[0][21] ),
    .A1(\design_top.MEM[1][21] ),
    .A2(\design_top.MEM[2][21] ),
    .A3(\design_top.MEM[3][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00533_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16868_ (.A0(\design_top.MEM[4][21] ),
    .A1(\design_top.MEM[5][21] ),
    .A2(\design_top.MEM[6][21] ),
    .A3(\design_top.MEM[7][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00534_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16869_ (.A0(\design_top.MEM[8][21] ),
    .A1(\design_top.MEM[9][21] ),
    .A2(\design_top.MEM[10][21] ),
    .A3(\design_top.MEM[11][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00535_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16870_ (.A0(\design_top.MEM[12][21] ),
    .A1(\design_top.MEM[13][21] ),
    .A2(\design_top.MEM[14][21] ),
    .A3(\design_top.MEM[15][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00536_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16871_ (.A0(_00533_),
    .A1(_00534_),
    .A2(_00535_),
    .A3(_00536_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00537_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16872_ (.A0(\design_top.MEM[16][21] ),
    .A1(\design_top.MEM[17][21] ),
    .A2(\design_top.MEM[18][21] ),
    .A3(\design_top.MEM[19][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00538_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16873_ (.A0(\design_top.MEM[20][21] ),
    .A1(\design_top.MEM[21][21] ),
    .A2(\design_top.MEM[22][21] ),
    .A3(\design_top.MEM[23][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00539_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16874_ (.A0(\design_top.MEM[24][21] ),
    .A1(\design_top.MEM[25][21] ),
    .A2(\design_top.MEM[26][21] ),
    .A3(\design_top.MEM[27][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00540_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16875_ (.A0(\design_top.MEM[28][21] ),
    .A1(\design_top.MEM[29][21] ),
    .A2(\design_top.MEM[30][21] ),
    .A3(\design_top.MEM[31][21] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00541_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16876_ (.A0(_00538_),
    .A1(_00539_),
    .A2(_00540_),
    .A3(_00541_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00542_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16877_ (.A0(\design_top.MEM[0][20] ),
    .A1(\design_top.MEM[1][20] ),
    .A2(\design_top.MEM[2][20] ),
    .A3(\design_top.MEM[3][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00523_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16878_ (.A0(\design_top.MEM[4][20] ),
    .A1(\design_top.MEM[5][20] ),
    .A2(\design_top.MEM[6][20] ),
    .A3(\design_top.MEM[7][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00524_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16879_ (.A0(\design_top.MEM[8][20] ),
    .A1(\design_top.MEM[9][20] ),
    .A2(\design_top.MEM[10][20] ),
    .A3(\design_top.MEM[11][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00525_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16880_ (.A0(\design_top.MEM[12][20] ),
    .A1(\design_top.MEM[13][20] ),
    .A2(\design_top.MEM[14][20] ),
    .A3(\design_top.MEM[15][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00526_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16881_ (.A0(_00523_),
    .A1(_00524_),
    .A2(_00525_),
    .A3(_00526_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00527_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16882_ (.A0(\design_top.MEM[16][20] ),
    .A1(\design_top.MEM[17][20] ),
    .A2(\design_top.MEM[18][20] ),
    .A3(\design_top.MEM[19][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00528_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16883_ (.A0(\design_top.MEM[20][20] ),
    .A1(\design_top.MEM[21][20] ),
    .A2(\design_top.MEM[22][20] ),
    .A3(\design_top.MEM[23][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00529_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16884_ (.A0(\design_top.MEM[24][20] ),
    .A1(\design_top.MEM[25][20] ),
    .A2(\design_top.MEM[26][20] ),
    .A3(\design_top.MEM[27][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00530_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16885_ (.A0(\design_top.MEM[28][20] ),
    .A1(\design_top.MEM[29][20] ),
    .A2(\design_top.MEM[30][20] ),
    .A3(\design_top.MEM[31][20] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00531_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16886_ (.A0(_00528_),
    .A1(_00529_),
    .A2(_00530_),
    .A3(_00531_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00532_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16887_ (.A0(\design_top.MEM[0][19] ),
    .A1(\design_top.MEM[1][19] ),
    .A2(\design_top.MEM[2][19] ),
    .A3(\design_top.MEM[3][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00513_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16888_ (.A0(\design_top.MEM[4][19] ),
    .A1(\design_top.MEM[5][19] ),
    .A2(\design_top.MEM[6][19] ),
    .A3(\design_top.MEM[7][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00514_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16889_ (.A0(\design_top.MEM[8][19] ),
    .A1(\design_top.MEM[9][19] ),
    .A2(\design_top.MEM[10][19] ),
    .A3(\design_top.MEM[11][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00515_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16890_ (.A0(\design_top.MEM[12][19] ),
    .A1(\design_top.MEM[13][19] ),
    .A2(\design_top.MEM[14][19] ),
    .A3(\design_top.MEM[15][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00516_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16891_ (.A0(_00513_),
    .A1(_00514_),
    .A2(_00515_),
    .A3(_00516_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00517_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16892_ (.A0(\design_top.MEM[16][19] ),
    .A1(\design_top.MEM[17][19] ),
    .A2(\design_top.MEM[18][19] ),
    .A3(\design_top.MEM[19][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00518_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16893_ (.A0(\design_top.MEM[20][19] ),
    .A1(\design_top.MEM[21][19] ),
    .A2(\design_top.MEM[22][19] ),
    .A3(\design_top.MEM[23][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00519_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16894_ (.A0(\design_top.MEM[24][19] ),
    .A1(\design_top.MEM[25][19] ),
    .A2(\design_top.MEM[26][19] ),
    .A3(\design_top.MEM[27][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00520_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16895_ (.A0(\design_top.MEM[28][19] ),
    .A1(\design_top.MEM[29][19] ),
    .A2(\design_top.MEM[30][19] ),
    .A3(\design_top.MEM[31][19] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00521_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16896_ (.A0(_00518_),
    .A1(_00519_),
    .A2(_00520_),
    .A3(_00521_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00522_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16897_ (.A0(\design_top.MEM[0][18] ),
    .A1(\design_top.MEM[1][18] ),
    .A2(\design_top.MEM[2][18] ),
    .A3(\design_top.MEM[3][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00503_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16898_ (.A0(\design_top.MEM[4][18] ),
    .A1(\design_top.MEM[5][18] ),
    .A2(\design_top.MEM[6][18] ),
    .A3(\design_top.MEM[7][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00504_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16899_ (.A0(\design_top.MEM[8][18] ),
    .A1(\design_top.MEM[9][18] ),
    .A2(\design_top.MEM[10][18] ),
    .A3(\design_top.MEM[11][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00505_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16900_ (.A0(\design_top.MEM[12][18] ),
    .A1(\design_top.MEM[13][18] ),
    .A2(\design_top.MEM[14][18] ),
    .A3(\design_top.MEM[15][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00506_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16901_ (.A0(_00503_),
    .A1(_00504_),
    .A2(_00505_),
    .A3(_00506_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00507_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16902_ (.A0(\design_top.MEM[16][18] ),
    .A1(\design_top.MEM[17][18] ),
    .A2(\design_top.MEM[18][18] ),
    .A3(\design_top.MEM[19][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00508_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16903_ (.A0(\design_top.MEM[20][18] ),
    .A1(\design_top.MEM[21][18] ),
    .A2(\design_top.MEM[22][18] ),
    .A3(\design_top.MEM[23][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00509_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16904_ (.A0(\design_top.MEM[24][18] ),
    .A1(\design_top.MEM[25][18] ),
    .A2(\design_top.MEM[26][18] ),
    .A3(\design_top.MEM[27][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00510_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16905_ (.A0(\design_top.MEM[28][18] ),
    .A1(\design_top.MEM[29][18] ),
    .A2(\design_top.MEM[30][18] ),
    .A3(\design_top.MEM[31][18] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00511_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16906_ (.A0(_00508_),
    .A1(_00509_),
    .A2(_00510_),
    .A3(_00511_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00512_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16907_ (.A0(\design_top.MEM[0][17] ),
    .A1(\design_top.MEM[1][17] ),
    .A2(\design_top.MEM[2][17] ),
    .A3(\design_top.MEM[3][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00493_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16908_ (.A0(\design_top.MEM[4][17] ),
    .A1(\design_top.MEM[5][17] ),
    .A2(\design_top.MEM[6][17] ),
    .A3(\design_top.MEM[7][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00494_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16909_ (.A0(\design_top.MEM[8][17] ),
    .A1(\design_top.MEM[9][17] ),
    .A2(\design_top.MEM[10][17] ),
    .A3(\design_top.MEM[11][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00495_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16910_ (.A0(\design_top.MEM[12][17] ),
    .A1(\design_top.MEM[13][17] ),
    .A2(\design_top.MEM[14][17] ),
    .A3(\design_top.MEM[15][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00496_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16911_ (.A0(_00493_),
    .A1(_00494_),
    .A2(_00495_),
    .A3(_00496_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00497_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16912_ (.A0(\design_top.MEM[16][17] ),
    .A1(\design_top.MEM[17][17] ),
    .A2(\design_top.MEM[18][17] ),
    .A3(\design_top.MEM[19][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00498_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16913_ (.A0(\design_top.MEM[20][17] ),
    .A1(\design_top.MEM[21][17] ),
    .A2(\design_top.MEM[22][17] ),
    .A3(\design_top.MEM[23][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00499_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16914_ (.A0(\design_top.MEM[24][17] ),
    .A1(\design_top.MEM[25][17] ),
    .A2(\design_top.MEM[26][17] ),
    .A3(\design_top.MEM[27][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00500_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16915_ (.A0(\design_top.MEM[28][17] ),
    .A1(\design_top.MEM[29][17] ),
    .A2(\design_top.MEM[30][17] ),
    .A3(\design_top.MEM[31][17] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00501_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16916_ (.A0(_00498_),
    .A1(_00499_),
    .A2(_00500_),
    .A3(_00501_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00502_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16917_ (.A0(\design_top.MEM[0][16] ),
    .A1(\design_top.MEM[1][16] ),
    .A2(\design_top.MEM[2][16] ),
    .A3(\design_top.MEM[3][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00483_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16918_ (.A0(\design_top.MEM[4][16] ),
    .A1(\design_top.MEM[5][16] ),
    .A2(\design_top.MEM[6][16] ),
    .A3(\design_top.MEM[7][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00484_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16919_ (.A0(\design_top.MEM[8][16] ),
    .A1(\design_top.MEM[9][16] ),
    .A2(\design_top.MEM[10][16] ),
    .A3(\design_top.MEM[11][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00485_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16920_ (.A0(\design_top.MEM[12][16] ),
    .A1(\design_top.MEM[13][16] ),
    .A2(\design_top.MEM[14][16] ),
    .A3(\design_top.MEM[15][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00486_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16921_ (.A0(_00483_),
    .A1(_00484_),
    .A2(_00485_),
    .A3(_00486_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00487_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16922_ (.A0(\design_top.MEM[16][16] ),
    .A1(\design_top.MEM[17][16] ),
    .A2(\design_top.MEM[18][16] ),
    .A3(\design_top.MEM[19][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00488_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16923_ (.A0(\design_top.MEM[20][16] ),
    .A1(\design_top.MEM[21][16] ),
    .A2(\design_top.MEM[22][16] ),
    .A3(\design_top.MEM[23][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00489_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16924_ (.A0(\design_top.MEM[24][16] ),
    .A1(\design_top.MEM[25][16] ),
    .A2(\design_top.MEM[26][16] ),
    .A3(\design_top.MEM[27][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00490_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16925_ (.A0(\design_top.MEM[28][16] ),
    .A1(\design_top.MEM[29][16] ),
    .A2(\design_top.MEM[30][16] ),
    .A3(\design_top.MEM[31][16] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00491_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16926_ (.A0(_00488_),
    .A1(_00489_),
    .A2(_00490_),
    .A3(_00491_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00492_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16927_ (.A0(\design_top.MEM[0][15] ),
    .A1(\design_top.MEM[1][15] ),
    .A2(\design_top.MEM[2][15] ),
    .A3(\design_top.MEM[3][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00473_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16928_ (.A0(\design_top.MEM[4][15] ),
    .A1(\design_top.MEM[5][15] ),
    .A2(\design_top.MEM[6][15] ),
    .A3(\design_top.MEM[7][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00474_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16929_ (.A0(\design_top.MEM[8][15] ),
    .A1(\design_top.MEM[9][15] ),
    .A2(\design_top.MEM[10][15] ),
    .A3(\design_top.MEM[11][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00475_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16930_ (.A0(\design_top.MEM[12][15] ),
    .A1(\design_top.MEM[13][15] ),
    .A2(\design_top.MEM[14][15] ),
    .A3(\design_top.MEM[15][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00476_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16931_ (.A0(_00473_),
    .A1(_00474_),
    .A2(_00475_),
    .A3(_00476_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00477_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16932_ (.A0(\design_top.MEM[16][15] ),
    .A1(\design_top.MEM[17][15] ),
    .A2(\design_top.MEM[18][15] ),
    .A3(\design_top.MEM[19][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00478_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16933_ (.A0(\design_top.MEM[20][15] ),
    .A1(\design_top.MEM[21][15] ),
    .A2(\design_top.MEM[22][15] ),
    .A3(\design_top.MEM[23][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00479_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16934_ (.A0(\design_top.MEM[24][15] ),
    .A1(\design_top.MEM[25][15] ),
    .A2(\design_top.MEM[26][15] ),
    .A3(\design_top.MEM[27][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00480_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16935_ (.A0(\design_top.MEM[28][15] ),
    .A1(\design_top.MEM[29][15] ),
    .A2(\design_top.MEM[30][15] ),
    .A3(\design_top.MEM[31][15] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00481_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16936_ (.A0(_00478_),
    .A1(_00479_),
    .A2(_00480_),
    .A3(_00481_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00482_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16937_ (.A0(\design_top.MEM[0][14] ),
    .A1(\design_top.MEM[1][14] ),
    .A2(\design_top.MEM[2][14] ),
    .A3(\design_top.MEM[3][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00463_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16938_ (.A0(\design_top.MEM[4][14] ),
    .A1(\design_top.MEM[5][14] ),
    .A2(\design_top.MEM[6][14] ),
    .A3(\design_top.MEM[7][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00464_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16939_ (.A0(\design_top.MEM[8][14] ),
    .A1(\design_top.MEM[9][14] ),
    .A2(\design_top.MEM[10][14] ),
    .A3(\design_top.MEM[11][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00465_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16940_ (.A0(\design_top.MEM[12][14] ),
    .A1(\design_top.MEM[13][14] ),
    .A2(\design_top.MEM[14][14] ),
    .A3(\design_top.MEM[15][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00466_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16941_ (.A0(_00463_),
    .A1(_00464_),
    .A2(_00465_),
    .A3(_00466_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00467_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16942_ (.A0(\design_top.MEM[16][14] ),
    .A1(\design_top.MEM[17][14] ),
    .A2(\design_top.MEM[18][14] ),
    .A3(\design_top.MEM[19][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00468_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16943_ (.A0(\design_top.MEM[20][14] ),
    .A1(\design_top.MEM[21][14] ),
    .A2(\design_top.MEM[22][14] ),
    .A3(\design_top.MEM[23][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00469_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16944_ (.A0(\design_top.MEM[24][14] ),
    .A1(\design_top.MEM[25][14] ),
    .A2(\design_top.MEM[26][14] ),
    .A3(\design_top.MEM[27][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00470_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16945_ (.A0(\design_top.MEM[28][14] ),
    .A1(\design_top.MEM[29][14] ),
    .A2(\design_top.MEM[30][14] ),
    .A3(\design_top.MEM[31][14] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00471_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16946_ (.A0(_00468_),
    .A1(_00469_),
    .A2(_00470_),
    .A3(_00471_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00472_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16947_ (.A0(\design_top.MEM[0][13] ),
    .A1(\design_top.MEM[1][13] ),
    .A2(\design_top.MEM[2][13] ),
    .A3(\design_top.MEM[3][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00453_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16948_ (.A0(\design_top.MEM[4][13] ),
    .A1(\design_top.MEM[5][13] ),
    .A2(\design_top.MEM[6][13] ),
    .A3(\design_top.MEM[7][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00454_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16949_ (.A0(\design_top.MEM[8][13] ),
    .A1(\design_top.MEM[9][13] ),
    .A2(\design_top.MEM[10][13] ),
    .A3(\design_top.MEM[11][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00455_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16950_ (.A0(\design_top.MEM[12][13] ),
    .A1(\design_top.MEM[13][13] ),
    .A2(\design_top.MEM[14][13] ),
    .A3(\design_top.MEM[15][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00456_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16951_ (.A0(_00453_),
    .A1(_00454_),
    .A2(_00455_),
    .A3(_00456_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00457_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16952_ (.A0(\design_top.MEM[16][13] ),
    .A1(\design_top.MEM[17][13] ),
    .A2(\design_top.MEM[18][13] ),
    .A3(\design_top.MEM[19][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00458_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16953_ (.A0(\design_top.MEM[20][13] ),
    .A1(\design_top.MEM[21][13] ),
    .A2(\design_top.MEM[22][13] ),
    .A3(\design_top.MEM[23][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00459_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16954_ (.A0(\design_top.MEM[24][13] ),
    .A1(\design_top.MEM[25][13] ),
    .A2(\design_top.MEM[26][13] ),
    .A3(\design_top.MEM[27][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00460_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16955_ (.A0(\design_top.MEM[28][13] ),
    .A1(\design_top.MEM[29][13] ),
    .A2(\design_top.MEM[30][13] ),
    .A3(\design_top.MEM[31][13] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00461_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16956_ (.A0(_00458_),
    .A1(_00459_),
    .A2(_00460_),
    .A3(_00461_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00462_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16957_ (.A0(\design_top.MEM[0][12] ),
    .A1(\design_top.MEM[1][12] ),
    .A2(\design_top.MEM[2][12] ),
    .A3(\design_top.MEM[3][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00443_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16958_ (.A0(\design_top.MEM[4][12] ),
    .A1(\design_top.MEM[5][12] ),
    .A2(\design_top.MEM[6][12] ),
    .A3(\design_top.MEM[7][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00444_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16959_ (.A0(\design_top.MEM[8][12] ),
    .A1(\design_top.MEM[9][12] ),
    .A2(\design_top.MEM[10][12] ),
    .A3(\design_top.MEM[11][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00445_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16960_ (.A0(\design_top.MEM[12][12] ),
    .A1(\design_top.MEM[13][12] ),
    .A2(\design_top.MEM[14][12] ),
    .A3(\design_top.MEM[15][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00446_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16961_ (.A0(_00443_),
    .A1(_00444_),
    .A2(_00445_),
    .A3(_00446_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00447_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16962_ (.A0(\design_top.MEM[16][12] ),
    .A1(\design_top.MEM[17][12] ),
    .A2(\design_top.MEM[18][12] ),
    .A3(\design_top.MEM[19][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00448_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16963_ (.A0(\design_top.MEM[20][12] ),
    .A1(\design_top.MEM[21][12] ),
    .A2(\design_top.MEM[22][12] ),
    .A3(\design_top.MEM[23][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00449_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16964_ (.A0(\design_top.MEM[24][12] ),
    .A1(\design_top.MEM[25][12] ),
    .A2(\design_top.MEM[26][12] ),
    .A3(\design_top.MEM[27][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00450_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16965_ (.A0(\design_top.MEM[28][12] ),
    .A1(\design_top.MEM[29][12] ),
    .A2(\design_top.MEM[30][12] ),
    .A3(\design_top.MEM[31][12] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00451_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16966_ (.A0(_00448_),
    .A1(_00449_),
    .A2(_00450_),
    .A3(_00451_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00452_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16967_ (.A0(\design_top.MEM[0][11] ),
    .A1(\design_top.MEM[1][11] ),
    .A2(\design_top.MEM[2][11] ),
    .A3(\design_top.MEM[3][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03055_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16968_ (.A0(\design_top.MEM[4][11] ),
    .A1(\design_top.MEM[5][11] ),
    .A2(\design_top.MEM[6][11] ),
    .A3(\design_top.MEM[7][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03056_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16969_ (.A0(\design_top.MEM[8][11] ),
    .A1(\design_top.MEM[9][11] ),
    .A2(\design_top.MEM[10][11] ),
    .A3(\design_top.MEM[11][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16970_ (.A0(\design_top.MEM[12][11] ),
    .A1(\design_top.MEM[13][11] ),
    .A2(\design_top.MEM[14][11] ),
    .A3(\design_top.MEM[15][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03058_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16971_ (.A0(_03055_),
    .A1(_03056_),
    .A2(_03057_),
    .A3(_03058_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00437_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16972_ (.A0(\design_top.MEM[16][11] ),
    .A1(\design_top.MEM[17][11] ),
    .A2(\design_top.MEM[18][11] ),
    .A3(\design_top.MEM[19][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00438_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16973_ (.A0(\design_top.MEM[20][11] ),
    .A1(\design_top.MEM[21][11] ),
    .A2(\design_top.MEM[22][11] ),
    .A3(\design_top.MEM[23][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00439_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16974_ (.A0(\design_top.MEM[24][11] ),
    .A1(\design_top.MEM[25][11] ),
    .A2(\design_top.MEM[26][11] ),
    .A3(\design_top.MEM[27][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00440_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16975_ (.A0(\design_top.MEM[28][11] ),
    .A1(\design_top.MEM[29][11] ),
    .A2(\design_top.MEM[30][11] ),
    .A3(\design_top.MEM[31][11] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_00441_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16976_ (.A0(_00438_),
    .A1(_00439_),
    .A2(_00440_),
    .A3(_00441_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_00442_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16977_ (.A0(\design_top.MEM[0][10] ),
    .A1(\design_top.MEM[1][10] ),
    .A2(\design_top.MEM[2][10] ),
    .A3(\design_top.MEM[3][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16978_ (.A0(\design_top.MEM[4][10] ),
    .A1(\design_top.MEM[5][10] ),
    .A2(\design_top.MEM[6][10] ),
    .A3(\design_top.MEM[7][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16979_ (.A0(\design_top.MEM[8][10] ),
    .A1(\design_top.MEM[9][10] ),
    .A2(\design_top.MEM[10][10] ),
    .A3(\design_top.MEM[11][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16980_ (.A0(\design_top.MEM[12][10] ),
    .A1(\design_top.MEM[13][10] ),
    .A2(\design_top.MEM[14][10] ),
    .A3(\design_top.MEM[15][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16981_ (.A0(_03045_),
    .A1(_03046_),
    .A2(_03047_),
    .A3(_03048_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03049_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16982_ (.A0(\design_top.MEM[16][10] ),
    .A1(\design_top.MEM[17][10] ),
    .A2(\design_top.MEM[18][10] ),
    .A3(\design_top.MEM[19][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03050_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16983_ (.A0(\design_top.MEM[20][10] ),
    .A1(\design_top.MEM[21][10] ),
    .A2(\design_top.MEM[22][10] ),
    .A3(\design_top.MEM[23][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16984_ (.A0(\design_top.MEM[24][10] ),
    .A1(\design_top.MEM[25][10] ),
    .A2(\design_top.MEM[26][10] ),
    .A3(\design_top.MEM[27][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16985_ (.A0(\design_top.MEM[28][10] ),
    .A1(\design_top.MEM[29][10] ),
    .A2(\design_top.MEM[30][10] ),
    .A3(\design_top.MEM[31][10] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03053_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16986_ (.A0(_03050_),
    .A1(_03051_),
    .A2(_03052_),
    .A3(_03053_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16987_ (.A0(\design_top.MEM[0][9] ),
    .A1(\design_top.MEM[1][9] ),
    .A2(\design_top.MEM[2][9] ),
    .A3(\design_top.MEM[3][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03035_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16988_ (.A0(\design_top.MEM[4][9] ),
    .A1(\design_top.MEM[5][9] ),
    .A2(\design_top.MEM[6][9] ),
    .A3(\design_top.MEM[7][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16989_ (.A0(\design_top.MEM[8][9] ),
    .A1(\design_top.MEM[9][9] ),
    .A2(\design_top.MEM[10][9] ),
    .A3(\design_top.MEM[11][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16990_ (.A0(\design_top.MEM[12][9] ),
    .A1(\design_top.MEM[13][9] ),
    .A2(\design_top.MEM[14][9] ),
    .A3(\design_top.MEM[15][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16991_ (.A0(_03035_),
    .A1(_03036_),
    .A2(_03037_),
    .A3(_03038_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03039_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16992_ (.A0(\design_top.MEM[16][9] ),
    .A1(\design_top.MEM[17][9] ),
    .A2(\design_top.MEM[18][9] ),
    .A3(\design_top.MEM[19][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16993_ (.A0(\design_top.MEM[20][9] ),
    .A1(\design_top.MEM[21][9] ),
    .A2(\design_top.MEM[22][9] ),
    .A3(\design_top.MEM[23][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16994_ (.A0(\design_top.MEM[24][9] ),
    .A1(\design_top.MEM[25][9] ),
    .A2(\design_top.MEM[26][9] ),
    .A3(\design_top.MEM[27][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16995_ (.A0(\design_top.MEM[28][9] ),
    .A1(\design_top.MEM[29][9] ),
    .A2(\design_top.MEM[30][9] ),
    .A3(\design_top.MEM[31][9] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16996_ (.A0(_03040_),
    .A1(_03041_),
    .A2(_03042_),
    .A3(_03043_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16997_ (.A0(\design_top.MEM[0][8] ),
    .A1(\design_top.MEM[1][8] ),
    .A2(\design_top.MEM[2][8] ),
    .A3(\design_top.MEM[3][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16998_ (.A0(\design_top.MEM[4][8] ),
    .A1(\design_top.MEM[5][8] ),
    .A2(\design_top.MEM[6][8] ),
    .A3(\design_top.MEM[7][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03026_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _16999_ (.A0(\design_top.MEM[8][8] ),
    .A1(\design_top.MEM[9][8] ),
    .A2(\design_top.MEM[10][8] ),
    .A3(\design_top.MEM[11][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17000_ (.A0(\design_top.MEM[12][8] ),
    .A1(\design_top.MEM[13][8] ),
    .A2(\design_top.MEM[14][8] ),
    .A3(\design_top.MEM[15][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17001_ (.A0(_03025_),
    .A1(_03026_),
    .A2(_03027_),
    .A3(_03028_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03029_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17002_ (.A0(\design_top.MEM[16][8] ),
    .A1(\design_top.MEM[17][8] ),
    .A2(\design_top.MEM[18][8] ),
    .A3(\design_top.MEM[19][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03030_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17003_ (.A0(\design_top.MEM[20][8] ),
    .A1(\design_top.MEM[21][8] ),
    .A2(\design_top.MEM[22][8] ),
    .A3(\design_top.MEM[23][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17004_ (.A0(\design_top.MEM[24][8] ),
    .A1(\design_top.MEM[25][8] ),
    .A2(\design_top.MEM[26][8] ),
    .A3(\design_top.MEM[27][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03032_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17005_ (.A0(\design_top.MEM[28][8] ),
    .A1(\design_top.MEM[29][8] ),
    .A2(\design_top.MEM[30][8] ),
    .A3(\design_top.MEM[31][8] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03033_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17006_ (.A0(_03030_),
    .A1(_03031_),
    .A2(_03032_),
    .A3(_03033_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17007_ (.A0(\design_top.MEM[0][7] ),
    .A1(\design_top.MEM[1][7] ),
    .A2(\design_top.MEM[2][7] ),
    .A3(\design_top.MEM[3][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03015_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17008_ (.A0(\design_top.MEM[4][7] ),
    .A1(\design_top.MEM[5][7] ),
    .A2(\design_top.MEM[6][7] ),
    .A3(\design_top.MEM[7][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17009_ (.A0(\design_top.MEM[8][7] ),
    .A1(\design_top.MEM[9][7] ),
    .A2(\design_top.MEM[10][7] ),
    .A3(\design_top.MEM[11][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03017_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17010_ (.A0(\design_top.MEM[12][7] ),
    .A1(\design_top.MEM[13][7] ),
    .A2(\design_top.MEM[14][7] ),
    .A3(\design_top.MEM[15][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17011_ (.A0(_03015_),
    .A1(_03016_),
    .A2(_03017_),
    .A3(_03018_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17012_ (.A0(\design_top.MEM[16][7] ),
    .A1(\design_top.MEM[17][7] ),
    .A2(\design_top.MEM[18][7] ),
    .A3(\design_top.MEM[19][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17013_ (.A0(\design_top.MEM[20][7] ),
    .A1(\design_top.MEM[21][7] ),
    .A2(\design_top.MEM[22][7] ),
    .A3(\design_top.MEM[23][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03021_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17014_ (.A0(\design_top.MEM[24][7] ),
    .A1(\design_top.MEM[25][7] ),
    .A2(\design_top.MEM[26][7] ),
    .A3(\design_top.MEM[27][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17015_ (.A0(\design_top.MEM[28][7] ),
    .A1(\design_top.MEM[29][7] ),
    .A2(\design_top.MEM[30][7] ),
    .A3(\design_top.MEM[31][7] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17016_ (.A0(_03020_),
    .A1(_03021_),
    .A2(_03022_),
    .A3(_03023_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03024_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17017_ (.A0(\design_top.MEM[0][6] ),
    .A1(\design_top.MEM[1][6] ),
    .A2(\design_top.MEM[2][6] ),
    .A3(\design_top.MEM[3][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03005_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17018_ (.A0(\design_top.MEM[4][6] ),
    .A1(\design_top.MEM[5][6] ),
    .A2(\design_top.MEM[6][6] ),
    .A3(\design_top.MEM[7][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03006_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17019_ (.A0(\design_top.MEM[8][6] ),
    .A1(\design_top.MEM[9][6] ),
    .A2(\design_top.MEM[10][6] ),
    .A3(\design_top.MEM[11][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17020_ (.A0(\design_top.MEM[12][6] ),
    .A1(\design_top.MEM[13][6] ),
    .A2(\design_top.MEM[14][6] ),
    .A3(\design_top.MEM[15][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17021_ (.A0(_03005_),
    .A1(_03006_),
    .A2(_03007_),
    .A3(_03008_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17022_ (.A0(\design_top.MEM[16][6] ),
    .A1(\design_top.MEM[17][6] ),
    .A2(\design_top.MEM[18][6] ),
    .A3(\design_top.MEM[19][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17023_ (.A0(\design_top.MEM[20][6] ),
    .A1(\design_top.MEM[21][6] ),
    .A2(\design_top.MEM[22][6] ),
    .A3(\design_top.MEM[23][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17024_ (.A0(\design_top.MEM[24][6] ),
    .A1(\design_top.MEM[25][6] ),
    .A2(\design_top.MEM[26][6] ),
    .A3(\design_top.MEM[27][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17025_ (.A0(\design_top.MEM[28][6] ),
    .A1(\design_top.MEM[29][6] ),
    .A2(\design_top.MEM[30][6] ),
    .A3(\design_top.MEM[31][6] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17026_ (.A0(_03010_),
    .A1(_03011_),
    .A2(_03012_),
    .A3(_03013_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17027_ (.A0(\design_top.MEM[0][5] ),
    .A1(\design_top.MEM[1][5] ),
    .A2(\design_top.MEM[2][5] ),
    .A3(\design_top.MEM[3][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02995_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17028_ (.A0(\design_top.MEM[4][5] ),
    .A1(\design_top.MEM[5][5] ),
    .A2(\design_top.MEM[6][5] ),
    .A3(\design_top.MEM[7][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02996_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17029_ (.A0(\design_top.MEM[8][5] ),
    .A1(\design_top.MEM[9][5] ),
    .A2(\design_top.MEM[10][5] ),
    .A3(\design_top.MEM[11][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02997_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17030_ (.A0(\design_top.MEM[12][5] ),
    .A1(\design_top.MEM[13][5] ),
    .A2(\design_top.MEM[14][5] ),
    .A3(\design_top.MEM[15][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02998_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17031_ (.A0(_02995_),
    .A1(_02996_),
    .A2(_02997_),
    .A3(_02998_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_02999_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17032_ (.A0(\design_top.MEM[16][5] ),
    .A1(\design_top.MEM[17][5] ),
    .A2(\design_top.MEM[18][5] ),
    .A3(\design_top.MEM[19][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17033_ (.A0(\design_top.MEM[20][5] ),
    .A1(\design_top.MEM[21][5] ),
    .A2(\design_top.MEM[22][5] ),
    .A3(\design_top.MEM[23][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17034_ (.A0(\design_top.MEM[24][5] ),
    .A1(\design_top.MEM[25][5] ),
    .A2(\design_top.MEM[26][5] ),
    .A3(\design_top.MEM[27][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17035_ (.A0(\design_top.MEM[28][5] ),
    .A1(\design_top.MEM[29][5] ),
    .A2(\design_top.MEM[30][5] ),
    .A3(\design_top.MEM[31][5] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_03003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17036_ (.A0(_03000_),
    .A1(_03001_),
    .A2(_03002_),
    .A3(_03003_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_03004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17037_ (.A0(\design_top.MEM[0][4] ),
    .A1(\design_top.MEM[1][4] ),
    .A2(\design_top.MEM[2][4] ),
    .A3(\design_top.MEM[3][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02985_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17038_ (.A0(\design_top.MEM[4][4] ),
    .A1(\design_top.MEM[5][4] ),
    .A2(\design_top.MEM[6][4] ),
    .A3(\design_top.MEM[7][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02986_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17039_ (.A0(\design_top.MEM[8][4] ),
    .A1(\design_top.MEM[9][4] ),
    .A2(\design_top.MEM[10][4] ),
    .A3(\design_top.MEM[11][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02987_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17040_ (.A0(\design_top.MEM[12][4] ),
    .A1(\design_top.MEM[13][4] ),
    .A2(\design_top.MEM[14][4] ),
    .A3(\design_top.MEM[15][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02988_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17041_ (.A0(_02985_),
    .A1(_02986_),
    .A2(_02987_),
    .A3(_02988_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_02989_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17042_ (.A0(\design_top.MEM[16][4] ),
    .A1(\design_top.MEM[17][4] ),
    .A2(\design_top.MEM[18][4] ),
    .A3(\design_top.MEM[19][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02990_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17043_ (.A0(\design_top.MEM[20][4] ),
    .A1(\design_top.MEM[21][4] ),
    .A2(\design_top.MEM[22][4] ),
    .A3(\design_top.MEM[23][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02991_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17044_ (.A0(\design_top.MEM[24][4] ),
    .A1(\design_top.MEM[25][4] ),
    .A2(\design_top.MEM[26][4] ),
    .A3(\design_top.MEM[27][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02992_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17045_ (.A0(\design_top.MEM[28][4] ),
    .A1(\design_top.MEM[29][4] ),
    .A2(\design_top.MEM[30][4] ),
    .A3(\design_top.MEM[31][4] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02993_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17046_ (.A0(_02990_),
    .A1(_02991_),
    .A2(_02992_),
    .A3(_02993_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_02994_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17047_ (.A0(\design_top.MEM[0][3] ),
    .A1(\design_top.MEM[1][3] ),
    .A2(\design_top.MEM[2][3] ),
    .A3(\design_top.MEM[3][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02975_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17048_ (.A0(\design_top.MEM[4][3] ),
    .A1(\design_top.MEM[5][3] ),
    .A2(\design_top.MEM[6][3] ),
    .A3(\design_top.MEM[7][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02976_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17049_ (.A0(\design_top.MEM[8][3] ),
    .A1(\design_top.MEM[9][3] ),
    .A2(\design_top.MEM[10][3] ),
    .A3(\design_top.MEM[11][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02977_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17050_ (.A0(\design_top.MEM[12][3] ),
    .A1(\design_top.MEM[13][3] ),
    .A2(\design_top.MEM[14][3] ),
    .A3(\design_top.MEM[15][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02978_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17051_ (.A0(_02975_),
    .A1(_02976_),
    .A2(_02977_),
    .A3(_02978_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_02979_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17052_ (.A0(\design_top.MEM[16][3] ),
    .A1(\design_top.MEM[17][3] ),
    .A2(\design_top.MEM[18][3] ),
    .A3(\design_top.MEM[19][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02980_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17053_ (.A0(\design_top.MEM[20][3] ),
    .A1(\design_top.MEM[21][3] ),
    .A2(\design_top.MEM[22][3] ),
    .A3(\design_top.MEM[23][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02981_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17054_ (.A0(\design_top.MEM[24][3] ),
    .A1(\design_top.MEM[25][3] ),
    .A2(\design_top.MEM[26][3] ),
    .A3(\design_top.MEM[27][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02982_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17055_ (.A0(\design_top.MEM[28][3] ),
    .A1(\design_top.MEM[29][3] ),
    .A2(\design_top.MEM[30][3] ),
    .A3(\design_top.MEM[31][3] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02983_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17056_ (.A0(_02980_),
    .A1(_02981_),
    .A2(_02982_),
    .A3(_02983_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_02984_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17057_ (.A0(\design_top.MEM[0][2] ),
    .A1(\design_top.MEM[1][2] ),
    .A2(\design_top.MEM[2][2] ),
    .A3(\design_top.MEM[3][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02965_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17058_ (.A0(\design_top.MEM[4][2] ),
    .A1(\design_top.MEM[5][2] ),
    .A2(\design_top.MEM[6][2] ),
    .A3(\design_top.MEM[7][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02966_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17059_ (.A0(\design_top.MEM[8][2] ),
    .A1(\design_top.MEM[9][2] ),
    .A2(\design_top.MEM[10][2] ),
    .A3(\design_top.MEM[11][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02967_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17060_ (.A0(\design_top.MEM[12][2] ),
    .A1(\design_top.MEM[13][2] ),
    .A2(\design_top.MEM[14][2] ),
    .A3(\design_top.MEM[15][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02968_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17061_ (.A0(_02965_),
    .A1(_02966_),
    .A2(_02967_),
    .A3(_02968_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_02969_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17062_ (.A0(\design_top.MEM[16][2] ),
    .A1(\design_top.MEM[17][2] ),
    .A2(\design_top.MEM[18][2] ),
    .A3(\design_top.MEM[19][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02970_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17063_ (.A0(\design_top.MEM[20][2] ),
    .A1(\design_top.MEM[21][2] ),
    .A2(\design_top.MEM[22][2] ),
    .A3(\design_top.MEM[23][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02971_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17064_ (.A0(\design_top.MEM[24][2] ),
    .A1(\design_top.MEM[25][2] ),
    .A2(\design_top.MEM[26][2] ),
    .A3(\design_top.MEM[27][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02972_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17065_ (.A0(\design_top.MEM[28][2] ),
    .A1(\design_top.MEM[29][2] ),
    .A2(\design_top.MEM[30][2] ),
    .A3(\design_top.MEM[31][2] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02973_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17066_ (.A0(_02970_),
    .A1(_02971_),
    .A2(_02972_),
    .A3(_02973_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_02974_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17067_ (.A0(\design_top.MEM[0][1] ),
    .A1(\design_top.MEM[1][1] ),
    .A2(\design_top.MEM[2][1] ),
    .A3(\design_top.MEM[3][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02955_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17068_ (.A0(\design_top.MEM[4][1] ),
    .A1(\design_top.MEM[5][1] ),
    .A2(\design_top.MEM[6][1] ),
    .A3(\design_top.MEM[7][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02956_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17069_ (.A0(\design_top.MEM[8][1] ),
    .A1(\design_top.MEM[9][1] ),
    .A2(\design_top.MEM[10][1] ),
    .A3(\design_top.MEM[11][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02957_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17070_ (.A0(\design_top.MEM[12][1] ),
    .A1(\design_top.MEM[13][1] ),
    .A2(\design_top.MEM[14][1] ),
    .A3(\design_top.MEM[15][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02958_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17071_ (.A0(_02955_),
    .A1(_02956_),
    .A2(_02957_),
    .A3(_02958_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_02959_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17072_ (.A0(\design_top.MEM[16][1] ),
    .A1(\design_top.MEM[17][1] ),
    .A2(\design_top.MEM[18][1] ),
    .A3(\design_top.MEM[19][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02960_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17073_ (.A0(\design_top.MEM[20][1] ),
    .A1(\design_top.MEM[21][1] ),
    .A2(\design_top.MEM[22][1] ),
    .A3(\design_top.MEM[23][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02961_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17074_ (.A0(\design_top.MEM[24][1] ),
    .A1(\design_top.MEM[25][1] ),
    .A2(\design_top.MEM[26][1] ),
    .A3(\design_top.MEM[27][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02962_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17075_ (.A0(\design_top.MEM[28][1] ),
    .A1(\design_top.MEM[29][1] ),
    .A2(\design_top.MEM[30][1] ),
    .A3(\design_top.MEM[31][1] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02963_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17076_ (.A0(_02960_),
    .A1(_02961_),
    .A2(_02962_),
    .A3(_02963_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_02964_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17077_ (.A0(\design_top.MEM[0][0] ),
    .A1(\design_top.MEM[1][0] ),
    .A2(\design_top.MEM[2][0] ),
    .A3(\design_top.MEM[3][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02945_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17078_ (.A0(\design_top.MEM[4][0] ),
    .A1(\design_top.MEM[5][0] ),
    .A2(\design_top.MEM[6][0] ),
    .A3(\design_top.MEM[7][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02946_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17079_ (.A0(\design_top.MEM[8][0] ),
    .A1(\design_top.MEM[9][0] ),
    .A2(\design_top.MEM[10][0] ),
    .A3(\design_top.MEM[11][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02947_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17080_ (.A0(\design_top.MEM[12][0] ),
    .A1(\design_top.MEM[13][0] ),
    .A2(\design_top.MEM[14][0] ),
    .A3(\design_top.MEM[15][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02948_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17081_ (.A0(_02945_),
    .A1(_02946_),
    .A2(_02947_),
    .A3(_02948_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_02949_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17082_ (.A0(\design_top.MEM[16][0] ),
    .A1(\design_top.MEM[17][0] ),
    .A2(\design_top.MEM[18][0] ),
    .A3(\design_top.MEM[19][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02950_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17083_ (.A0(\design_top.MEM[20][0] ),
    .A1(\design_top.MEM[21][0] ),
    .A2(\design_top.MEM[22][0] ),
    .A3(\design_top.MEM[23][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02951_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17084_ (.A0(\design_top.MEM[24][0] ),
    .A1(\design_top.MEM[25][0] ),
    .A2(\design_top.MEM[26][0] ),
    .A3(\design_top.MEM[27][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02952_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17085_ (.A0(\design_top.MEM[28][0] ),
    .A1(\design_top.MEM[29][0] ),
    .A2(\design_top.MEM[30][0] ),
    .A3(\design_top.MEM[31][0] ),
    .S0(io_out[18]),
    .S1(io_out[19]),
    .X(_02953_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17086_ (.A0(_02950_),
    .A1(_02951_),
    .A2(_02952_),
    .A3(_02953_),
    .S0(\design_top.IADDR[4] ),
    .S1(\design_top.IADDR[5] ),
    .X(_02954_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17087_ (.A0(\design_top.MEM[31][31] ),
    .A1(\design_top.MEM[30][31] ),
    .A2(\design_top.MEM[29][31] ),
    .A3(\design_top.MEM[28][31] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02910_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17088_ (.A0(\design_top.MEM[27][31] ),
    .A1(\design_top.MEM[26][31] ),
    .A2(\design_top.MEM[25][31] ),
    .A3(\design_top.MEM[24][31] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02909_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17089_ (.A0(\design_top.MEM[23][31] ),
    .A1(\design_top.MEM[22][31] ),
    .A2(\design_top.MEM[21][31] ),
    .A3(\design_top.MEM[20][31] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02908_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17090_ (.A0(\design_top.MEM[19][31] ),
    .A1(\design_top.MEM[18][31] ),
    .A2(\design_top.MEM[17][31] ),
    .A3(\design_top.MEM[16][31] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02907_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17091_ (.A0(_02910_),
    .A1(_02909_),
    .A2(_02908_),
    .A3(_02907_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02911_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17092_ (.A0(\design_top.MEM[15][31] ),
    .A1(\design_top.MEM[14][31] ),
    .A2(\design_top.MEM[13][31] ),
    .A3(\design_top.MEM[12][31] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02905_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17093_ (.A0(\design_top.MEM[11][31] ),
    .A1(\design_top.MEM[10][31] ),
    .A2(\design_top.MEM[9][31] ),
    .A3(\design_top.MEM[8][31] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02904_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17094_ (.A0(\design_top.MEM[7][31] ),
    .A1(\design_top.MEM[6][31] ),
    .A2(\design_top.MEM[5][31] ),
    .A3(\design_top.MEM[4][31] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02903_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17095_ (.A0(\design_top.MEM[3][31] ),
    .A1(\design_top.MEM[2][31] ),
    .A2(\design_top.MEM[1][31] ),
    .A3(\design_top.MEM[0][31] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02902_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17096_ (.A0(_02905_),
    .A1(_02904_),
    .A2(_02903_),
    .A3(_02902_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02906_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17097_ (.A0(\design_top.MEM[31][30] ),
    .A1(\design_top.MEM[30][30] ),
    .A2(\design_top.MEM[29][30] ),
    .A3(\design_top.MEM[28][30] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02900_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17098_ (.A0(\design_top.MEM[27][30] ),
    .A1(\design_top.MEM[26][30] ),
    .A2(\design_top.MEM[25][30] ),
    .A3(\design_top.MEM[24][30] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02899_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17099_ (.A0(\design_top.MEM[23][30] ),
    .A1(\design_top.MEM[22][30] ),
    .A2(\design_top.MEM[21][30] ),
    .A3(\design_top.MEM[20][30] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02898_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17100_ (.A0(\design_top.MEM[19][30] ),
    .A1(\design_top.MEM[18][30] ),
    .A2(\design_top.MEM[17][30] ),
    .A3(\design_top.MEM[16][30] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02897_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17101_ (.A0(_02900_),
    .A1(_02899_),
    .A2(_02898_),
    .A3(_02897_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02901_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17102_ (.A0(\design_top.MEM[15][30] ),
    .A1(\design_top.MEM[14][30] ),
    .A2(\design_top.MEM[13][30] ),
    .A3(\design_top.MEM[12][30] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02895_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17103_ (.A0(\design_top.MEM[11][30] ),
    .A1(\design_top.MEM[10][30] ),
    .A2(\design_top.MEM[9][30] ),
    .A3(\design_top.MEM[8][30] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02894_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17104_ (.A0(\design_top.MEM[7][30] ),
    .A1(\design_top.MEM[6][30] ),
    .A2(\design_top.MEM[5][30] ),
    .A3(\design_top.MEM[4][30] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02893_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17105_ (.A0(\design_top.MEM[3][30] ),
    .A1(\design_top.MEM[2][30] ),
    .A2(\design_top.MEM[1][30] ),
    .A3(\design_top.MEM[0][30] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02892_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17106_ (.A0(_02895_),
    .A1(_02894_),
    .A2(_02893_),
    .A3(_02892_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02896_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17107_ (.A0(\design_top.MEM[31][29] ),
    .A1(\design_top.MEM[30][29] ),
    .A2(\design_top.MEM[29][29] ),
    .A3(\design_top.MEM[28][29] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02890_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17108_ (.A0(\design_top.MEM[27][29] ),
    .A1(\design_top.MEM[26][29] ),
    .A2(\design_top.MEM[25][29] ),
    .A3(\design_top.MEM[24][29] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02889_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17109_ (.A0(\design_top.MEM[23][29] ),
    .A1(\design_top.MEM[22][29] ),
    .A2(\design_top.MEM[21][29] ),
    .A3(\design_top.MEM[20][29] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02888_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17110_ (.A0(\design_top.MEM[19][29] ),
    .A1(\design_top.MEM[18][29] ),
    .A2(\design_top.MEM[17][29] ),
    .A3(\design_top.MEM[16][29] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02887_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17111_ (.A0(_02890_),
    .A1(_02889_),
    .A2(_02888_),
    .A3(_02887_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02891_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17112_ (.A0(\design_top.MEM[15][29] ),
    .A1(\design_top.MEM[14][29] ),
    .A2(\design_top.MEM[13][29] ),
    .A3(\design_top.MEM[12][29] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02885_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17113_ (.A0(\design_top.MEM[11][29] ),
    .A1(\design_top.MEM[10][29] ),
    .A2(\design_top.MEM[9][29] ),
    .A3(\design_top.MEM[8][29] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02884_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17114_ (.A0(\design_top.MEM[7][29] ),
    .A1(\design_top.MEM[6][29] ),
    .A2(\design_top.MEM[5][29] ),
    .A3(\design_top.MEM[4][29] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02883_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17115_ (.A0(\design_top.MEM[3][29] ),
    .A1(\design_top.MEM[2][29] ),
    .A2(\design_top.MEM[1][29] ),
    .A3(\design_top.MEM[0][29] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02882_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17116_ (.A0(_02885_),
    .A1(_02884_),
    .A2(_02883_),
    .A3(_02882_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02886_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17117_ (.A0(\design_top.MEM[31][28] ),
    .A1(\design_top.MEM[30][28] ),
    .A2(\design_top.MEM[29][28] ),
    .A3(\design_top.MEM[28][28] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02880_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17118_ (.A0(\design_top.MEM[27][28] ),
    .A1(\design_top.MEM[26][28] ),
    .A2(\design_top.MEM[25][28] ),
    .A3(\design_top.MEM[24][28] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02879_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17119_ (.A0(\design_top.MEM[23][28] ),
    .A1(\design_top.MEM[22][28] ),
    .A2(\design_top.MEM[21][28] ),
    .A3(\design_top.MEM[20][28] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02878_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17120_ (.A0(\design_top.MEM[19][28] ),
    .A1(\design_top.MEM[18][28] ),
    .A2(\design_top.MEM[17][28] ),
    .A3(\design_top.MEM[16][28] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02877_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17121_ (.A0(_02880_),
    .A1(_02879_),
    .A2(_02878_),
    .A3(_02877_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02881_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17122_ (.A0(\design_top.MEM[15][28] ),
    .A1(\design_top.MEM[14][28] ),
    .A2(\design_top.MEM[13][28] ),
    .A3(\design_top.MEM[12][28] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02875_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17123_ (.A0(\design_top.MEM[11][28] ),
    .A1(\design_top.MEM[10][28] ),
    .A2(\design_top.MEM[9][28] ),
    .A3(\design_top.MEM[8][28] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02874_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17124_ (.A0(\design_top.MEM[7][28] ),
    .A1(\design_top.MEM[6][28] ),
    .A2(\design_top.MEM[5][28] ),
    .A3(\design_top.MEM[4][28] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02873_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17125_ (.A0(\design_top.MEM[3][28] ),
    .A1(\design_top.MEM[2][28] ),
    .A2(\design_top.MEM[1][28] ),
    .A3(\design_top.MEM[0][28] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02872_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17126_ (.A0(_02875_),
    .A1(_02874_),
    .A2(_02873_),
    .A3(_02872_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02876_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17127_ (.A0(\design_top.MEM[31][27] ),
    .A1(\design_top.MEM[30][27] ),
    .A2(\design_top.MEM[29][27] ),
    .A3(\design_top.MEM[28][27] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02870_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17128_ (.A0(\design_top.MEM[27][27] ),
    .A1(\design_top.MEM[26][27] ),
    .A2(\design_top.MEM[25][27] ),
    .A3(\design_top.MEM[24][27] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02869_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17129_ (.A0(\design_top.MEM[23][27] ),
    .A1(\design_top.MEM[22][27] ),
    .A2(\design_top.MEM[21][27] ),
    .A3(\design_top.MEM[20][27] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02868_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17130_ (.A0(\design_top.MEM[19][27] ),
    .A1(\design_top.MEM[18][27] ),
    .A2(\design_top.MEM[17][27] ),
    .A3(\design_top.MEM[16][27] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02867_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17131_ (.A0(_02870_),
    .A1(_02869_),
    .A2(_02868_),
    .A3(_02867_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02871_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17132_ (.A0(\design_top.MEM[15][27] ),
    .A1(\design_top.MEM[14][27] ),
    .A2(\design_top.MEM[13][27] ),
    .A3(\design_top.MEM[12][27] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02865_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17133_ (.A0(\design_top.MEM[11][27] ),
    .A1(\design_top.MEM[10][27] ),
    .A2(\design_top.MEM[9][27] ),
    .A3(\design_top.MEM[8][27] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02864_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17134_ (.A0(\design_top.MEM[7][27] ),
    .A1(\design_top.MEM[6][27] ),
    .A2(\design_top.MEM[5][27] ),
    .A3(\design_top.MEM[4][27] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02863_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17135_ (.A0(\design_top.MEM[3][27] ),
    .A1(\design_top.MEM[2][27] ),
    .A2(\design_top.MEM[1][27] ),
    .A3(\design_top.MEM[0][27] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02862_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17136_ (.A0(_02865_),
    .A1(_02864_),
    .A2(_02863_),
    .A3(_02862_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02866_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17137_ (.A0(\design_top.MEM[31][26] ),
    .A1(\design_top.MEM[30][26] ),
    .A2(\design_top.MEM[29][26] ),
    .A3(\design_top.MEM[28][26] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02860_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17138_ (.A0(\design_top.MEM[27][26] ),
    .A1(\design_top.MEM[26][26] ),
    .A2(\design_top.MEM[25][26] ),
    .A3(\design_top.MEM[24][26] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02859_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17139_ (.A0(\design_top.MEM[23][26] ),
    .A1(\design_top.MEM[22][26] ),
    .A2(\design_top.MEM[21][26] ),
    .A3(\design_top.MEM[20][26] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02858_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17140_ (.A0(\design_top.MEM[19][26] ),
    .A1(\design_top.MEM[18][26] ),
    .A2(\design_top.MEM[17][26] ),
    .A3(\design_top.MEM[16][26] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02857_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17141_ (.A0(_02860_),
    .A1(_02859_),
    .A2(_02858_),
    .A3(_02857_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02861_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17142_ (.A0(\design_top.MEM[15][26] ),
    .A1(\design_top.MEM[14][26] ),
    .A2(\design_top.MEM[13][26] ),
    .A3(\design_top.MEM[12][26] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02855_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17143_ (.A0(\design_top.MEM[11][26] ),
    .A1(\design_top.MEM[10][26] ),
    .A2(\design_top.MEM[9][26] ),
    .A3(\design_top.MEM[8][26] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02854_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17144_ (.A0(\design_top.MEM[7][26] ),
    .A1(\design_top.MEM[6][26] ),
    .A2(\design_top.MEM[5][26] ),
    .A3(\design_top.MEM[4][26] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02853_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17145_ (.A0(\design_top.MEM[3][26] ),
    .A1(\design_top.MEM[2][26] ),
    .A2(\design_top.MEM[1][26] ),
    .A3(\design_top.MEM[0][26] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02852_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17146_ (.A0(_02855_),
    .A1(_02854_),
    .A2(_02853_),
    .A3(_02852_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02856_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17147_ (.A0(\design_top.MEM[31][25] ),
    .A1(\design_top.MEM[30][25] ),
    .A2(\design_top.MEM[29][25] ),
    .A3(\design_top.MEM[28][25] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02850_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17148_ (.A0(\design_top.MEM[27][25] ),
    .A1(\design_top.MEM[26][25] ),
    .A2(\design_top.MEM[25][25] ),
    .A3(\design_top.MEM[24][25] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02849_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17149_ (.A0(\design_top.MEM[23][25] ),
    .A1(\design_top.MEM[22][25] ),
    .A2(\design_top.MEM[21][25] ),
    .A3(\design_top.MEM[20][25] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02848_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17150_ (.A0(\design_top.MEM[19][25] ),
    .A1(\design_top.MEM[18][25] ),
    .A2(\design_top.MEM[17][25] ),
    .A3(\design_top.MEM[16][25] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02847_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17151_ (.A0(_02850_),
    .A1(_02849_),
    .A2(_02848_),
    .A3(_02847_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02851_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17152_ (.A0(\design_top.MEM[15][25] ),
    .A1(\design_top.MEM[14][25] ),
    .A2(\design_top.MEM[13][25] ),
    .A3(\design_top.MEM[12][25] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02845_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17153_ (.A0(\design_top.MEM[11][25] ),
    .A1(\design_top.MEM[10][25] ),
    .A2(\design_top.MEM[9][25] ),
    .A3(\design_top.MEM[8][25] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02844_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17154_ (.A0(\design_top.MEM[7][25] ),
    .A1(\design_top.MEM[6][25] ),
    .A2(\design_top.MEM[5][25] ),
    .A3(\design_top.MEM[4][25] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02843_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17155_ (.A0(\design_top.MEM[3][25] ),
    .A1(\design_top.MEM[2][25] ),
    .A2(\design_top.MEM[1][25] ),
    .A3(\design_top.MEM[0][25] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02842_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17156_ (.A0(_02845_),
    .A1(_02844_),
    .A2(_02843_),
    .A3(_02842_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02846_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17157_ (.A0(\design_top.MEM[31][24] ),
    .A1(\design_top.MEM[30][24] ),
    .A2(\design_top.MEM[29][24] ),
    .A3(\design_top.MEM[28][24] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02840_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17158_ (.A0(\design_top.MEM[27][24] ),
    .A1(\design_top.MEM[26][24] ),
    .A2(\design_top.MEM[25][24] ),
    .A3(\design_top.MEM[24][24] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02839_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17159_ (.A0(\design_top.MEM[23][24] ),
    .A1(\design_top.MEM[22][24] ),
    .A2(\design_top.MEM[21][24] ),
    .A3(\design_top.MEM[20][24] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02838_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17160_ (.A0(\design_top.MEM[19][24] ),
    .A1(\design_top.MEM[18][24] ),
    .A2(\design_top.MEM[17][24] ),
    .A3(\design_top.MEM[16][24] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02837_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17161_ (.A0(_02840_),
    .A1(_02839_),
    .A2(_02838_),
    .A3(_02837_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02841_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17162_ (.A0(\design_top.MEM[15][24] ),
    .A1(\design_top.MEM[14][24] ),
    .A2(\design_top.MEM[13][24] ),
    .A3(\design_top.MEM[12][24] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02835_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17163_ (.A0(\design_top.MEM[11][24] ),
    .A1(\design_top.MEM[10][24] ),
    .A2(\design_top.MEM[9][24] ),
    .A3(\design_top.MEM[8][24] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02834_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17164_ (.A0(\design_top.MEM[7][24] ),
    .A1(\design_top.MEM[6][24] ),
    .A2(\design_top.MEM[5][24] ),
    .A3(\design_top.MEM[4][24] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02833_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17165_ (.A0(\design_top.MEM[3][24] ),
    .A1(\design_top.MEM[2][24] ),
    .A2(\design_top.MEM[1][24] ),
    .A3(\design_top.MEM[0][24] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02832_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17166_ (.A0(_02835_),
    .A1(_02834_),
    .A2(_02833_),
    .A3(_02832_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02836_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17167_ (.A0(\design_top.MEM[31][23] ),
    .A1(\design_top.MEM[30][23] ),
    .A2(\design_top.MEM[29][23] ),
    .A3(\design_top.MEM[28][23] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02830_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17168_ (.A0(\design_top.MEM[27][23] ),
    .A1(\design_top.MEM[26][23] ),
    .A2(\design_top.MEM[25][23] ),
    .A3(\design_top.MEM[24][23] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02829_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17169_ (.A0(\design_top.MEM[23][23] ),
    .A1(\design_top.MEM[22][23] ),
    .A2(\design_top.MEM[21][23] ),
    .A3(\design_top.MEM[20][23] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02828_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17170_ (.A0(\design_top.MEM[19][23] ),
    .A1(\design_top.MEM[18][23] ),
    .A2(\design_top.MEM[17][23] ),
    .A3(\design_top.MEM[16][23] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02827_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17171_ (.A0(_02830_),
    .A1(_02829_),
    .A2(_02828_),
    .A3(_02827_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02831_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17172_ (.A0(\design_top.MEM[15][23] ),
    .A1(\design_top.MEM[14][23] ),
    .A2(\design_top.MEM[13][23] ),
    .A3(\design_top.MEM[12][23] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02825_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17173_ (.A0(\design_top.MEM[11][23] ),
    .A1(\design_top.MEM[10][23] ),
    .A2(\design_top.MEM[9][23] ),
    .A3(\design_top.MEM[8][23] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02824_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17174_ (.A0(\design_top.MEM[7][23] ),
    .A1(\design_top.MEM[6][23] ),
    .A2(\design_top.MEM[5][23] ),
    .A3(\design_top.MEM[4][23] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02823_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17175_ (.A0(\design_top.MEM[3][23] ),
    .A1(\design_top.MEM[2][23] ),
    .A2(\design_top.MEM[1][23] ),
    .A3(\design_top.MEM[0][23] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02822_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17176_ (.A0(_02825_),
    .A1(_02824_),
    .A2(_02823_),
    .A3(_02822_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02826_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17177_ (.A0(\design_top.MEM[31][22] ),
    .A1(\design_top.MEM[30][22] ),
    .A2(\design_top.MEM[29][22] ),
    .A3(\design_top.MEM[28][22] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02820_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17178_ (.A0(\design_top.MEM[27][22] ),
    .A1(\design_top.MEM[26][22] ),
    .A2(\design_top.MEM[25][22] ),
    .A3(\design_top.MEM[24][22] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02819_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17179_ (.A0(\design_top.MEM[23][22] ),
    .A1(\design_top.MEM[22][22] ),
    .A2(\design_top.MEM[21][22] ),
    .A3(\design_top.MEM[20][22] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02818_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17180_ (.A0(\design_top.MEM[19][22] ),
    .A1(\design_top.MEM[18][22] ),
    .A2(\design_top.MEM[17][22] ),
    .A3(\design_top.MEM[16][22] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02817_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17181_ (.A0(_02820_),
    .A1(_02819_),
    .A2(_02818_),
    .A3(_02817_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02821_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17182_ (.A0(\design_top.MEM[15][22] ),
    .A1(\design_top.MEM[14][22] ),
    .A2(\design_top.MEM[13][22] ),
    .A3(\design_top.MEM[12][22] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02815_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17183_ (.A0(\design_top.MEM[11][22] ),
    .A1(\design_top.MEM[10][22] ),
    .A2(\design_top.MEM[9][22] ),
    .A3(\design_top.MEM[8][22] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02814_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17184_ (.A0(\design_top.MEM[7][22] ),
    .A1(\design_top.MEM[6][22] ),
    .A2(\design_top.MEM[5][22] ),
    .A3(\design_top.MEM[4][22] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02813_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17185_ (.A0(\design_top.MEM[3][22] ),
    .A1(\design_top.MEM[2][22] ),
    .A2(\design_top.MEM[1][22] ),
    .A3(\design_top.MEM[0][22] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02812_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17186_ (.A0(_02815_),
    .A1(_02814_),
    .A2(_02813_),
    .A3(_02812_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02816_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17187_ (.A0(\design_top.MEM[31][21] ),
    .A1(\design_top.MEM[30][21] ),
    .A2(\design_top.MEM[29][21] ),
    .A3(\design_top.MEM[28][21] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02810_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17188_ (.A0(\design_top.MEM[27][21] ),
    .A1(\design_top.MEM[26][21] ),
    .A2(\design_top.MEM[25][21] ),
    .A3(\design_top.MEM[24][21] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02809_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17189_ (.A0(\design_top.MEM[23][21] ),
    .A1(\design_top.MEM[22][21] ),
    .A2(\design_top.MEM[21][21] ),
    .A3(\design_top.MEM[20][21] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02808_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17190_ (.A0(\design_top.MEM[19][21] ),
    .A1(\design_top.MEM[18][21] ),
    .A2(\design_top.MEM[17][21] ),
    .A3(\design_top.MEM[16][21] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02807_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17191_ (.A0(_02810_),
    .A1(_02809_),
    .A2(_02808_),
    .A3(_02807_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02811_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17192_ (.A0(\design_top.MEM[15][21] ),
    .A1(\design_top.MEM[14][21] ),
    .A2(\design_top.MEM[13][21] ),
    .A3(\design_top.MEM[12][21] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02805_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17193_ (.A0(\design_top.MEM[11][21] ),
    .A1(\design_top.MEM[10][21] ),
    .A2(\design_top.MEM[9][21] ),
    .A3(\design_top.MEM[8][21] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02804_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17194_ (.A0(\design_top.MEM[7][21] ),
    .A1(\design_top.MEM[6][21] ),
    .A2(\design_top.MEM[5][21] ),
    .A3(\design_top.MEM[4][21] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02803_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17195_ (.A0(\design_top.MEM[3][21] ),
    .A1(\design_top.MEM[2][21] ),
    .A2(\design_top.MEM[1][21] ),
    .A3(\design_top.MEM[0][21] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02802_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17196_ (.A0(_02805_),
    .A1(_02804_),
    .A2(_02803_),
    .A3(_02802_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02806_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17197_ (.A0(\design_top.MEM[31][20] ),
    .A1(\design_top.MEM[30][20] ),
    .A2(\design_top.MEM[29][20] ),
    .A3(\design_top.MEM[28][20] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02800_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17198_ (.A0(\design_top.MEM[27][20] ),
    .A1(\design_top.MEM[26][20] ),
    .A2(\design_top.MEM[25][20] ),
    .A3(\design_top.MEM[24][20] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02799_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17199_ (.A0(\design_top.MEM[23][20] ),
    .A1(\design_top.MEM[22][20] ),
    .A2(\design_top.MEM[21][20] ),
    .A3(\design_top.MEM[20][20] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02798_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17200_ (.A0(\design_top.MEM[19][20] ),
    .A1(\design_top.MEM[18][20] ),
    .A2(\design_top.MEM[17][20] ),
    .A3(\design_top.MEM[16][20] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02797_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17201_ (.A0(_02800_),
    .A1(_02799_),
    .A2(_02798_),
    .A3(_02797_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02801_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17202_ (.A0(\design_top.MEM[15][20] ),
    .A1(\design_top.MEM[14][20] ),
    .A2(\design_top.MEM[13][20] ),
    .A3(\design_top.MEM[12][20] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02795_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17203_ (.A0(\design_top.MEM[11][20] ),
    .A1(\design_top.MEM[10][20] ),
    .A2(\design_top.MEM[9][20] ),
    .A3(\design_top.MEM[8][20] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02794_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17204_ (.A0(\design_top.MEM[7][20] ),
    .A1(\design_top.MEM[6][20] ),
    .A2(\design_top.MEM[5][20] ),
    .A3(\design_top.MEM[4][20] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02793_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17205_ (.A0(\design_top.MEM[3][20] ),
    .A1(\design_top.MEM[2][20] ),
    .A2(\design_top.MEM[1][20] ),
    .A3(\design_top.MEM[0][20] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02792_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17206_ (.A0(_02795_),
    .A1(_02794_),
    .A2(_02793_),
    .A3(_02792_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02796_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17207_ (.A0(\design_top.MEM[31][19] ),
    .A1(\design_top.MEM[30][19] ),
    .A2(\design_top.MEM[29][19] ),
    .A3(\design_top.MEM[28][19] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02790_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17208_ (.A0(\design_top.MEM[27][19] ),
    .A1(\design_top.MEM[26][19] ),
    .A2(\design_top.MEM[25][19] ),
    .A3(\design_top.MEM[24][19] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02789_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17209_ (.A0(\design_top.MEM[23][19] ),
    .A1(\design_top.MEM[22][19] ),
    .A2(\design_top.MEM[21][19] ),
    .A3(\design_top.MEM[20][19] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02788_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17210_ (.A0(\design_top.MEM[19][19] ),
    .A1(\design_top.MEM[18][19] ),
    .A2(\design_top.MEM[17][19] ),
    .A3(\design_top.MEM[16][19] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02787_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17211_ (.A0(_02790_),
    .A1(_02789_),
    .A2(_02788_),
    .A3(_02787_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02791_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17212_ (.A0(\design_top.MEM[15][19] ),
    .A1(\design_top.MEM[14][19] ),
    .A2(\design_top.MEM[13][19] ),
    .A3(\design_top.MEM[12][19] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02785_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17213_ (.A0(\design_top.MEM[11][19] ),
    .A1(\design_top.MEM[10][19] ),
    .A2(\design_top.MEM[9][19] ),
    .A3(\design_top.MEM[8][19] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02784_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17214_ (.A0(\design_top.MEM[7][19] ),
    .A1(\design_top.MEM[6][19] ),
    .A2(\design_top.MEM[5][19] ),
    .A3(\design_top.MEM[4][19] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02783_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17215_ (.A0(\design_top.MEM[3][19] ),
    .A1(\design_top.MEM[2][19] ),
    .A2(\design_top.MEM[1][19] ),
    .A3(\design_top.MEM[0][19] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02782_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17216_ (.A0(_02785_),
    .A1(_02784_),
    .A2(_02783_),
    .A3(_02782_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02786_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17217_ (.A0(\design_top.MEM[31][18] ),
    .A1(\design_top.MEM[30][18] ),
    .A2(\design_top.MEM[29][18] ),
    .A3(\design_top.MEM[28][18] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02780_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17218_ (.A0(\design_top.MEM[27][18] ),
    .A1(\design_top.MEM[26][18] ),
    .A2(\design_top.MEM[25][18] ),
    .A3(\design_top.MEM[24][18] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02779_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17219_ (.A0(\design_top.MEM[23][18] ),
    .A1(\design_top.MEM[22][18] ),
    .A2(\design_top.MEM[21][18] ),
    .A3(\design_top.MEM[20][18] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02778_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17220_ (.A0(\design_top.MEM[19][18] ),
    .A1(\design_top.MEM[18][18] ),
    .A2(\design_top.MEM[17][18] ),
    .A3(\design_top.MEM[16][18] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02777_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17221_ (.A0(_02780_),
    .A1(_02779_),
    .A2(_02778_),
    .A3(_02777_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02781_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17222_ (.A0(\design_top.MEM[15][18] ),
    .A1(\design_top.MEM[14][18] ),
    .A2(\design_top.MEM[13][18] ),
    .A3(\design_top.MEM[12][18] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02775_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17223_ (.A0(\design_top.MEM[11][18] ),
    .A1(\design_top.MEM[10][18] ),
    .A2(\design_top.MEM[9][18] ),
    .A3(\design_top.MEM[8][18] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02774_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17224_ (.A0(\design_top.MEM[7][18] ),
    .A1(\design_top.MEM[6][18] ),
    .A2(\design_top.MEM[5][18] ),
    .A3(\design_top.MEM[4][18] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02773_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17225_ (.A0(\design_top.MEM[3][18] ),
    .A1(\design_top.MEM[2][18] ),
    .A2(\design_top.MEM[1][18] ),
    .A3(\design_top.MEM[0][18] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02772_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17226_ (.A0(_02775_),
    .A1(_02774_),
    .A2(_02773_),
    .A3(_02772_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02776_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17227_ (.A0(\design_top.MEM[31][17] ),
    .A1(\design_top.MEM[30][17] ),
    .A2(\design_top.MEM[29][17] ),
    .A3(\design_top.MEM[28][17] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02770_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17228_ (.A0(\design_top.MEM[27][17] ),
    .A1(\design_top.MEM[26][17] ),
    .A2(\design_top.MEM[25][17] ),
    .A3(\design_top.MEM[24][17] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02769_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17229_ (.A0(\design_top.MEM[23][17] ),
    .A1(\design_top.MEM[22][17] ),
    .A2(\design_top.MEM[21][17] ),
    .A3(\design_top.MEM[20][17] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02768_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17230_ (.A0(\design_top.MEM[19][17] ),
    .A1(\design_top.MEM[18][17] ),
    .A2(\design_top.MEM[17][17] ),
    .A3(\design_top.MEM[16][17] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02767_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17231_ (.A0(_02770_),
    .A1(_02769_),
    .A2(_02768_),
    .A3(_02767_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02771_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17232_ (.A0(\design_top.MEM[15][17] ),
    .A1(\design_top.MEM[14][17] ),
    .A2(\design_top.MEM[13][17] ),
    .A3(\design_top.MEM[12][17] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02765_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17233_ (.A0(\design_top.MEM[11][17] ),
    .A1(\design_top.MEM[10][17] ),
    .A2(\design_top.MEM[9][17] ),
    .A3(\design_top.MEM[8][17] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02764_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17234_ (.A0(\design_top.MEM[7][17] ),
    .A1(\design_top.MEM[6][17] ),
    .A2(\design_top.MEM[5][17] ),
    .A3(\design_top.MEM[4][17] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02763_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17235_ (.A0(\design_top.MEM[3][17] ),
    .A1(\design_top.MEM[2][17] ),
    .A2(\design_top.MEM[1][17] ),
    .A3(\design_top.MEM[0][17] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02762_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17236_ (.A0(_02765_),
    .A1(_02764_),
    .A2(_02763_),
    .A3(_02762_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02766_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17237_ (.A0(\design_top.MEM[31][16] ),
    .A1(\design_top.MEM[30][16] ),
    .A2(\design_top.MEM[29][16] ),
    .A3(\design_top.MEM[28][16] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02760_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17238_ (.A0(\design_top.MEM[27][16] ),
    .A1(\design_top.MEM[26][16] ),
    .A2(\design_top.MEM[25][16] ),
    .A3(\design_top.MEM[24][16] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02759_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17239_ (.A0(\design_top.MEM[23][16] ),
    .A1(\design_top.MEM[22][16] ),
    .A2(\design_top.MEM[21][16] ),
    .A3(\design_top.MEM[20][16] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02758_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17240_ (.A0(\design_top.MEM[19][16] ),
    .A1(\design_top.MEM[18][16] ),
    .A2(\design_top.MEM[17][16] ),
    .A3(\design_top.MEM[16][16] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02757_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17241_ (.A0(_02760_),
    .A1(_02759_),
    .A2(_02758_),
    .A3(_02757_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02761_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17242_ (.A0(\design_top.MEM[15][16] ),
    .A1(\design_top.MEM[14][16] ),
    .A2(\design_top.MEM[13][16] ),
    .A3(\design_top.MEM[12][16] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02755_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17243_ (.A0(\design_top.MEM[11][16] ),
    .A1(\design_top.MEM[10][16] ),
    .A2(\design_top.MEM[9][16] ),
    .A3(\design_top.MEM[8][16] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02754_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17244_ (.A0(\design_top.MEM[7][16] ),
    .A1(\design_top.MEM[6][16] ),
    .A2(\design_top.MEM[5][16] ),
    .A3(\design_top.MEM[4][16] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02753_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17245_ (.A0(\design_top.MEM[3][16] ),
    .A1(\design_top.MEM[2][16] ),
    .A2(\design_top.MEM[1][16] ),
    .A3(\design_top.MEM[0][16] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02752_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17246_ (.A0(_02755_),
    .A1(_02754_),
    .A2(_02753_),
    .A3(_02752_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02756_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17247_ (.A0(\design_top.MEM[31][15] ),
    .A1(\design_top.MEM[30][15] ),
    .A2(\design_top.MEM[29][15] ),
    .A3(\design_top.MEM[28][15] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02750_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17248_ (.A0(\design_top.MEM[27][15] ),
    .A1(\design_top.MEM[26][15] ),
    .A2(\design_top.MEM[25][15] ),
    .A3(\design_top.MEM[24][15] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02749_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17249_ (.A0(\design_top.MEM[23][15] ),
    .A1(\design_top.MEM[22][15] ),
    .A2(\design_top.MEM[21][15] ),
    .A3(\design_top.MEM[20][15] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02748_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17250_ (.A0(\design_top.MEM[19][15] ),
    .A1(\design_top.MEM[18][15] ),
    .A2(\design_top.MEM[17][15] ),
    .A3(\design_top.MEM[16][15] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02747_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17251_ (.A0(_02750_),
    .A1(_02749_),
    .A2(_02748_),
    .A3(_02747_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02751_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17252_ (.A0(\design_top.MEM[15][15] ),
    .A1(\design_top.MEM[14][15] ),
    .A2(\design_top.MEM[13][15] ),
    .A3(\design_top.MEM[12][15] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02745_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17253_ (.A0(\design_top.MEM[11][15] ),
    .A1(\design_top.MEM[10][15] ),
    .A2(\design_top.MEM[9][15] ),
    .A3(\design_top.MEM[8][15] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02744_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17254_ (.A0(\design_top.MEM[7][15] ),
    .A1(\design_top.MEM[6][15] ),
    .A2(\design_top.MEM[5][15] ),
    .A3(\design_top.MEM[4][15] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02743_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17255_ (.A0(\design_top.MEM[3][15] ),
    .A1(\design_top.MEM[2][15] ),
    .A2(\design_top.MEM[1][15] ),
    .A3(\design_top.MEM[0][15] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02742_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17256_ (.A0(_02745_),
    .A1(_02744_),
    .A2(_02743_),
    .A3(_02742_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02746_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17257_ (.A0(\design_top.MEM[31][14] ),
    .A1(\design_top.MEM[30][14] ),
    .A2(\design_top.MEM[29][14] ),
    .A3(\design_top.MEM[28][14] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02740_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17258_ (.A0(\design_top.MEM[27][14] ),
    .A1(\design_top.MEM[26][14] ),
    .A2(\design_top.MEM[25][14] ),
    .A3(\design_top.MEM[24][14] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02739_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17259_ (.A0(\design_top.MEM[23][14] ),
    .A1(\design_top.MEM[22][14] ),
    .A2(\design_top.MEM[21][14] ),
    .A3(\design_top.MEM[20][14] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02738_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17260_ (.A0(\design_top.MEM[19][14] ),
    .A1(\design_top.MEM[18][14] ),
    .A2(\design_top.MEM[17][14] ),
    .A3(\design_top.MEM[16][14] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02737_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17261_ (.A0(_02740_),
    .A1(_02739_),
    .A2(_02738_),
    .A3(_02737_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02741_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17262_ (.A0(\design_top.MEM[15][14] ),
    .A1(\design_top.MEM[14][14] ),
    .A2(\design_top.MEM[13][14] ),
    .A3(\design_top.MEM[12][14] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02735_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17263_ (.A0(\design_top.MEM[11][14] ),
    .A1(\design_top.MEM[10][14] ),
    .A2(\design_top.MEM[9][14] ),
    .A3(\design_top.MEM[8][14] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02734_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17264_ (.A0(\design_top.MEM[7][14] ),
    .A1(\design_top.MEM[6][14] ),
    .A2(\design_top.MEM[5][14] ),
    .A3(\design_top.MEM[4][14] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02733_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17265_ (.A0(\design_top.MEM[3][14] ),
    .A1(\design_top.MEM[2][14] ),
    .A2(\design_top.MEM[1][14] ),
    .A3(\design_top.MEM[0][14] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02732_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17266_ (.A0(_02735_),
    .A1(_02734_),
    .A2(_02733_),
    .A3(_02732_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02736_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17267_ (.A0(\design_top.MEM[31][13] ),
    .A1(\design_top.MEM[30][13] ),
    .A2(\design_top.MEM[29][13] ),
    .A3(\design_top.MEM[28][13] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02730_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17268_ (.A0(\design_top.MEM[27][13] ),
    .A1(\design_top.MEM[26][13] ),
    .A2(\design_top.MEM[25][13] ),
    .A3(\design_top.MEM[24][13] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02729_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17269_ (.A0(\design_top.MEM[23][13] ),
    .A1(\design_top.MEM[22][13] ),
    .A2(\design_top.MEM[21][13] ),
    .A3(\design_top.MEM[20][13] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02728_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17270_ (.A0(\design_top.MEM[19][13] ),
    .A1(\design_top.MEM[18][13] ),
    .A2(\design_top.MEM[17][13] ),
    .A3(\design_top.MEM[16][13] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02727_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17271_ (.A0(_02730_),
    .A1(_02729_),
    .A2(_02728_),
    .A3(_02727_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02731_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17272_ (.A0(\design_top.MEM[15][13] ),
    .A1(\design_top.MEM[14][13] ),
    .A2(\design_top.MEM[13][13] ),
    .A3(\design_top.MEM[12][13] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02725_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17273_ (.A0(\design_top.MEM[11][13] ),
    .A1(\design_top.MEM[10][13] ),
    .A2(\design_top.MEM[9][13] ),
    .A3(\design_top.MEM[8][13] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02724_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17274_ (.A0(\design_top.MEM[7][13] ),
    .A1(\design_top.MEM[6][13] ),
    .A2(\design_top.MEM[5][13] ),
    .A3(\design_top.MEM[4][13] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02723_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17275_ (.A0(\design_top.MEM[3][13] ),
    .A1(\design_top.MEM[2][13] ),
    .A2(\design_top.MEM[1][13] ),
    .A3(\design_top.MEM[0][13] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02722_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17276_ (.A0(_02725_),
    .A1(_02724_),
    .A2(_02723_),
    .A3(_02722_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02726_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17277_ (.A0(\design_top.MEM[31][12] ),
    .A1(\design_top.MEM[30][12] ),
    .A2(\design_top.MEM[29][12] ),
    .A3(\design_top.MEM[28][12] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02720_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17278_ (.A0(\design_top.MEM[27][12] ),
    .A1(\design_top.MEM[26][12] ),
    .A2(\design_top.MEM[25][12] ),
    .A3(\design_top.MEM[24][12] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02719_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17279_ (.A0(\design_top.MEM[23][12] ),
    .A1(\design_top.MEM[22][12] ),
    .A2(\design_top.MEM[21][12] ),
    .A3(\design_top.MEM[20][12] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02718_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17280_ (.A0(\design_top.MEM[19][12] ),
    .A1(\design_top.MEM[18][12] ),
    .A2(\design_top.MEM[17][12] ),
    .A3(\design_top.MEM[16][12] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02717_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17281_ (.A0(_02720_),
    .A1(_02719_),
    .A2(_02718_),
    .A3(_02717_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02721_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17282_ (.A0(\design_top.MEM[15][12] ),
    .A1(\design_top.MEM[14][12] ),
    .A2(\design_top.MEM[13][12] ),
    .A3(\design_top.MEM[12][12] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02715_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17283_ (.A0(\design_top.MEM[11][12] ),
    .A1(\design_top.MEM[10][12] ),
    .A2(\design_top.MEM[9][12] ),
    .A3(\design_top.MEM[8][12] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02714_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17284_ (.A0(\design_top.MEM[7][12] ),
    .A1(\design_top.MEM[6][12] ),
    .A2(\design_top.MEM[5][12] ),
    .A3(\design_top.MEM[4][12] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02713_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17285_ (.A0(\design_top.MEM[3][12] ),
    .A1(\design_top.MEM[2][12] ),
    .A2(\design_top.MEM[1][12] ),
    .A3(\design_top.MEM[0][12] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02712_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17286_ (.A0(_02715_),
    .A1(_02714_),
    .A2(_02713_),
    .A3(_02712_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02716_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17287_ (.A0(\design_top.MEM[31][11] ),
    .A1(\design_top.MEM[30][11] ),
    .A2(\design_top.MEM[29][11] ),
    .A3(\design_top.MEM[28][11] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02710_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17288_ (.A0(\design_top.MEM[27][11] ),
    .A1(\design_top.MEM[26][11] ),
    .A2(\design_top.MEM[25][11] ),
    .A3(\design_top.MEM[24][11] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02709_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17289_ (.A0(\design_top.MEM[23][11] ),
    .A1(\design_top.MEM[22][11] ),
    .A2(\design_top.MEM[21][11] ),
    .A3(\design_top.MEM[20][11] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02708_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17290_ (.A0(\design_top.MEM[19][11] ),
    .A1(\design_top.MEM[18][11] ),
    .A2(\design_top.MEM[17][11] ),
    .A3(\design_top.MEM[16][11] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02707_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17291_ (.A0(_02710_),
    .A1(_02709_),
    .A2(_02708_),
    .A3(_02707_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02711_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17292_ (.A0(\design_top.MEM[15][11] ),
    .A1(\design_top.MEM[14][11] ),
    .A2(\design_top.MEM[13][11] ),
    .A3(\design_top.MEM[12][11] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02705_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17293_ (.A0(\design_top.MEM[11][11] ),
    .A1(\design_top.MEM[10][11] ),
    .A2(\design_top.MEM[9][11] ),
    .A3(\design_top.MEM[8][11] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02704_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17294_ (.A0(\design_top.MEM[7][11] ),
    .A1(\design_top.MEM[6][11] ),
    .A2(\design_top.MEM[5][11] ),
    .A3(\design_top.MEM[4][11] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02703_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17295_ (.A0(\design_top.MEM[3][11] ),
    .A1(\design_top.MEM[2][11] ),
    .A2(\design_top.MEM[1][11] ),
    .A3(\design_top.MEM[0][11] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02702_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17296_ (.A0(_02705_),
    .A1(_02704_),
    .A2(_02703_),
    .A3(_02702_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02706_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17297_ (.A0(\design_top.MEM[31][10] ),
    .A1(\design_top.MEM[30][10] ),
    .A2(\design_top.MEM[29][10] ),
    .A3(\design_top.MEM[28][10] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02700_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17298_ (.A0(\design_top.MEM[27][10] ),
    .A1(\design_top.MEM[26][10] ),
    .A2(\design_top.MEM[25][10] ),
    .A3(\design_top.MEM[24][10] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02699_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17299_ (.A0(\design_top.MEM[23][10] ),
    .A1(\design_top.MEM[22][10] ),
    .A2(\design_top.MEM[21][10] ),
    .A3(\design_top.MEM[20][10] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02698_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17300_ (.A0(\design_top.MEM[19][10] ),
    .A1(\design_top.MEM[18][10] ),
    .A2(\design_top.MEM[17][10] ),
    .A3(\design_top.MEM[16][10] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02697_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17301_ (.A0(_02700_),
    .A1(_02699_),
    .A2(_02698_),
    .A3(_02697_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02701_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17302_ (.A0(\design_top.MEM[15][10] ),
    .A1(\design_top.MEM[14][10] ),
    .A2(\design_top.MEM[13][10] ),
    .A3(\design_top.MEM[12][10] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02695_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17303_ (.A0(\design_top.MEM[11][10] ),
    .A1(\design_top.MEM[10][10] ),
    .A2(\design_top.MEM[9][10] ),
    .A3(\design_top.MEM[8][10] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02694_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17304_ (.A0(\design_top.MEM[7][10] ),
    .A1(\design_top.MEM[6][10] ),
    .A2(\design_top.MEM[5][10] ),
    .A3(\design_top.MEM[4][10] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02693_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17305_ (.A0(\design_top.MEM[3][10] ),
    .A1(\design_top.MEM[2][10] ),
    .A2(\design_top.MEM[1][10] ),
    .A3(\design_top.MEM[0][10] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02692_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17306_ (.A0(_02695_),
    .A1(_02694_),
    .A2(_02693_),
    .A3(_02692_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02696_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17307_ (.A0(\design_top.MEM[31][9] ),
    .A1(\design_top.MEM[30][9] ),
    .A2(\design_top.MEM[29][9] ),
    .A3(\design_top.MEM[28][9] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02690_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17308_ (.A0(\design_top.MEM[27][9] ),
    .A1(\design_top.MEM[26][9] ),
    .A2(\design_top.MEM[25][9] ),
    .A3(\design_top.MEM[24][9] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02689_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17309_ (.A0(\design_top.MEM[23][9] ),
    .A1(\design_top.MEM[22][9] ),
    .A2(\design_top.MEM[21][9] ),
    .A3(\design_top.MEM[20][9] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02688_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17310_ (.A0(\design_top.MEM[19][9] ),
    .A1(\design_top.MEM[18][9] ),
    .A2(\design_top.MEM[17][9] ),
    .A3(\design_top.MEM[16][9] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02687_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17311_ (.A0(_02690_),
    .A1(_02689_),
    .A2(_02688_),
    .A3(_02687_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02691_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17312_ (.A0(\design_top.MEM[15][9] ),
    .A1(\design_top.MEM[14][9] ),
    .A2(\design_top.MEM[13][9] ),
    .A3(\design_top.MEM[12][9] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02685_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17313_ (.A0(\design_top.MEM[11][9] ),
    .A1(\design_top.MEM[10][9] ),
    .A2(\design_top.MEM[9][9] ),
    .A3(\design_top.MEM[8][9] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02684_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17314_ (.A0(\design_top.MEM[7][9] ),
    .A1(\design_top.MEM[6][9] ),
    .A2(\design_top.MEM[5][9] ),
    .A3(\design_top.MEM[4][9] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02683_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17315_ (.A0(\design_top.MEM[3][9] ),
    .A1(\design_top.MEM[2][9] ),
    .A2(\design_top.MEM[1][9] ),
    .A3(\design_top.MEM[0][9] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02682_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17316_ (.A0(_02685_),
    .A1(_02684_),
    .A2(_02683_),
    .A3(_02682_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02686_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17317_ (.A0(\design_top.MEM[31][8] ),
    .A1(\design_top.MEM[30][8] ),
    .A2(\design_top.MEM[29][8] ),
    .A3(\design_top.MEM[28][8] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02680_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17318_ (.A0(\design_top.MEM[27][8] ),
    .A1(\design_top.MEM[26][8] ),
    .A2(\design_top.MEM[25][8] ),
    .A3(\design_top.MEM[24][8] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02679_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17319_ (.A0(\design_top.MEM[23][8] ),
    .A1(\design_top.MEM[22][8] ),
    .A2(\design_top.MEM[21][8] ),
    .A3(\design_top.MEM[20][8] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02678_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17320_ (.A0(\design_top.MEM[19][8] ),
    .A1(\design_top.MEM[18][8] ),
    .A2(\design_top.MEM[17][8] ),
    .A3(\design_top.MEM[16][8] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02677_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17321_ (.A0(_02680_),
    .A1(_02679_),
    .A2(_02678_),
    .A3(_02677_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02681_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17322_ (.A0(\design_top.MEM[15][8] ),
    .A1(\design_top.MEM[14][8] ),
    .A2(\design_top.MEM[13][8] ),
    .A3(\design_top.MEM[12][8] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02675_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17323_ (.A0(\design_top.MEM[11][8] ),
    .A1(\design_top.MEM[10][8] ),
    .A2(\design_top.MEM[9][8] ),
    .A3(\design_top.MEM[8][8] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02674_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17324_ (.A0(\design_top.MEM[7][8] ),
    .A1(\design_top.MEM[6][8] ),
    .A2(\design_top.MEM[5][8] ),
    .A3(\design_top.MEM[4][8] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02673_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17325_ (.A0(\design_top.MEM[3][8] ),
    .A1(\design_top.MEM[2][8] ),
    .A2(\design_top.MEM[1][8] ),
    .A3(\design_top.MEM[0][8] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02672_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17326_ (.A0(_02675_),
    .A1(_02674_),
    .A2(_02673_),
    .A3(_02672_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02676_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17327_ (.A0(\design_top.MEM[31][7] ),
    .A1(\design_top.MEM[30][7] ),
    .A2(\design_top.MEM[29][7] ),
    .A3(\design_top.MEM[28][7] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02670_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17328_ (.A0(\design_top.MEM[27][7] ),
    .A1(\design_top.MEM[26][7] ),
    .A2(\design_top.MEM[25][7] ),
    .A3(\design_top.MEM[24][7] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02669_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17329_ (.A0(\design_top.MEM[23][7] ),
    .A1(\design_top.MEM[22][7] ),
    .A2(\design_top.MEM[21][7] ),
    .A3(\design_top.MEM[20][7] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02668_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17330_ (.A0(\design_top.MEM[19][7] ),
    .A1(\design_top.MEM[18][7] ),
    .A2(\design_top.MEM[17][7] ),
    .A3(\design_top.MEM[16][7] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02667_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17331_ (.A0(_02670_),
    .A1(_02669_),
    .A2(_02668_),
    .A3(_02667_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02671_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17332_ (.A0(\design_top.MEM[15][7] ),
    .A1(\design_top.MEM[14][7] ),
    .A2(\design_top.MEM[13][7] ),
    .A3(\design_top.MEM[12][7] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02665_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17333_ (.A0(\design_top.MEM[11][7] ),
    .A1(\design_top.MEM[10][7] ),
    .A2(\design_top.MEM[9][7] ),
    .A3(\design_top.MEM[8][7] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02664_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17334_ (.A0(\design_top.MEM[7][7] ),
    .A1(\design_top.MEM[6][7] ),
    .A2(\design_top.MEM[5][7] ),
    .A3(\design_top.MEM[4][7] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02663_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17335_ (.A0(\design_top.MEM[3][7] ),
    .A1(\design_top.MEM[2][7] ),
    .A2(\design_top.MEM[1][7] ),
    .A3(\design_top.MEM[0][7] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02662_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17336_ (.A0(_02665_),
    .A1(_02664_),
    .A2(_02663_),
    .A3(_02662_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02666_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17337_ (.A0(\design_top.MEM[31][6] ),
    .A1(\design_top.MEM[30][6] ),
    .A2(\design_top.MEM[29][6] ),
    .A3(\design_top.MEM[28][6] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02660_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17338_ (.A0(\design_top.MEM[27][6] ),
    .A1(\design_top.MEM[26][6] ),
    .A2(\design_top.MEM[25][6] ),
    .A3(\design_top.MEM[24][6] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02659_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17339_ (.A0(\design_top.MEM[23][6] ),
    .A1(\design_top.MEM[22][6] ),
    .A2(\design_top.MEM[21][6] ),
    .A3(\design_top.MEM[20][6] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02658_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17340_ (.A0(\design_top.MEM[19][6] ),
    .A1(\design_top.MEM[18][6] ),
    .A2(\design_top.MEM[17][6] ),
    .A3(\design_top.MEM[16][6] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02657_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17341_ (.A0(_02660_),
    .A1(_02659_),
    .A2(_02658_),
    .A3(_02657_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02661_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17342_ (.A0(\design_top.MEM[15][6] ),
    .A1(\design_top.MEM[14][6] ),
    .A2(\design_top.MEM[13][6] ),
    .A3(\design_top.MEM[12][6] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02655_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17343_ (.A0(\design_top.MEM[11][6] ),
    .A1(\design_top.MEM[10][6] ),
    .A2(\design_top.MEM[9][6] ),
    .A3(\design_top.MEM[8][6] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02654_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17344_ (.A0(\design_top.MEM[7][6] ),
    .A1(\design_top.MEM[6][6] ),
    .A2(\design_top.MEM[5][6] ),
    .A3(\design_top.MEM[4][6] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02653_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17345_ (.A0(\design_top.MEM[3][6] ),
    .A1(\design_top.MEM[2][6] ),
    .A2(\design_top.MEM[1][6] ),
    .A3(\design_top.MEM[0][6] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02652_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17346_ (.A0(_02655_),
    .A1(_02654_),
    .A2(_02653_),
    .A3(_02652_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02656_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17347_ (.A0(\design_top.MEM[31][5] ),
    .A1(\design_top.MEM[30][5] ),
    .A2(\design_top.MEM[29][5] ),
    .A3(\design_top.MEM[28][5] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02650_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17348_ (.A0(\design_top.MEM[27][5] ),
    .A1(\design_top.MEM[26][5] ),
    .A2(\design_top.MEM[25][5] ),
    .A3(\design_top.MEM[24][5] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02649_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17349_ (.A0(\design_top.MEM[23][5] ),
    .A1(\design_top.MEM[22][5] ),
    .A2(\design_top.MEM[21][5] ),
    .A3(\design_top.MEM[20][5] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02648_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17350_ (.A0(\design_top.MEM[19][5] ),
    .A1(\design_top.MEM[18][5] ),
    .A2(\design_top.MEM[17][5] ),
    .A3(\design_top.MEM[16][5] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02647_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17351_ (.A0(_02650_),
    .A1(_02649_),
    .A2(_02648_),
    .A3(_02647_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02651_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17352_ (.A0(\design_top.MEM[15][5] ),
    .A1(\design_top.MEM[14][5] ),
    .A2(\design_top.MEM[13][5] ),
    .A3(\design_top.MEM[12][5] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02645_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17353_ (.A0(\design_top.MEM[11][5] ),
    .A1(\design_top.MEM[10][5] ),
    .A2(\design_top.MEM[9][5] ),
    .A3(\design_top.MEM[8][5] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02644_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17354_ (.A0(\design_top.MEM[7][5] ),
    .A1(\design_top.MEM[6][5] ),
    .A2(\design_top.MEM[5][5] ),
    .A3(\design_top.MEM[4][5] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02643_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17355_ (.A0(\design_top.MEM[3][5] ),
    .A1(\design_top.MEM[2][5] ),
    .A2(\design_top.MEM[1][5] ),
    .A3(\design_top.MEM[0][5] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02642_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17356_ (.A0(_02645_),
    .A1(_02644_),
    .A2(_02643_),
    .A3(_02642_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02646_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17357_ (.A0(\design_top.MEM[31][4] ),
    .A1(\design_top.MEM[30][4] ),
    .A2(\design_top.MEM[29][4] ),
    .A3(\design_top.MEM[28][4] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02640_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17358_ (.A0(\design_top.MEM[27][4] ),
    .A1(\design_top.MEM[26][4] ),
    .A2(\design_top.MEM[25][4] ),
    .A3(\design_top.MEM[24][4] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02639_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17359_ (.A0(\design_top.MEM[23][4] ),
    .A1(\design_top.MEM[22][4] ),
    .A2(\design_top.MEM[21][4] ),
    .A3(\design_top.MEM[20][4] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02638_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17360_ (.A0(\design_top.MEM[19][4] ),
    .A1(\design_top.MEM[18][4] ),
    .A2(\design_top.MEM[17][4] ),
    .A3(\design_top.MEM[16][4] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02637_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17361_ (.A0(_02640_),
    .A1(_02639_),
    .A2(_02638_),
    .A3(_02637_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02641_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17362_ (.A0(\design_top.MEM[15][4] ),
    .A1(\design_top.MEM[14][4] ),
    .A2(\design_top.MEM[13][4] ),
    .A3(\design_top.MEM[12][4] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02635_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17363_ (.A0(\design_top.MEM[11][4] ),
    .A1(\design_top.MEM[10][4] ),
    .A2(\design_top.MEM[9][4] ),
    .A3(\design_top.MEM[8][4] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02634_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17364_ (.A0(\design_top.MEM[7][4] ),
    .A1(\design_top.MEM[6][4] ),
    .A2(\design_top.MEM[5][4] ),
    .A3(\design_top.MEM[4][4] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02633_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17365_ (.A0(\design_top.MEM[3][4] ),
    .A1(\design_top.MEM[2][4] ),
    .A2(\design_top.MEM[1][4] ),
    .A3(\design_top.MEM[0][4] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02632_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17366_ (.A0(_02635_),
    .A1(_02634_),
    .A2(_02633_),
    .A3(_02632_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02636_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17367_ (.A0(\design_top.MEM[31][3] ),
    .A1(\design_top.MEM[30][3] ),
    .A2(\design_top.MEM[29][3] ),
    .A3(\design_top.MEM[28][3] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02630_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17368_ (.A0(\design_top.MEM[27][3] ),
    .A1(\design_top.MEM[26][3] ),
    .A2(\design_top.MEM[25][3] ),
    .A3(\design_top.MEM[24][3] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02629_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17369_ (.A0(\design_top.MEM[23][3] ),
    .A1(\design_top.MEM[22][3] ),
    .A2(\design_top.MEM[21][3] ),
    .A3(\design_top.MEM[20][3] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02628_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17370_ (.A0(\design_top.MEM[19][3] ),
    .A1(\design_top.MEM[18][3] ),
    .A2(\design_top.MEM[17][3] ),
    .A3(\design_top.MEM[16][3] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02627_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17371_ (.A0(_02630_),
    .A1(_02629_),
    .A2(_02628_),
    .A3(_02627_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02631_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17372_ (.A0(\design_top.MEM[15][3] ),
    .A1(\design_top.MEM[14][3] ),
    .A2(\design_top.MEM[13][3] ),
    .A3(\design_top.MEM[12][3] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02625_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17373_ (.A0(\design_top.MEM[11][3] ),
    .A1(\design_top.MEM[10][3] ),
    .A2(\design_top.MEM[9][3] ),
    .A3(\design_top.MEM[8][3] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02624_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17374_ (.A0(\design_top.MEM[7][3] ),
    .A1(\design_top.MEM[6][3] ),
    .A2(\design_top.MEM[5][3] ),
    .A3(\design_top.MEM[4][3] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02623_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17375_ (.A0(\design_top.MEM[3][3] ),
    .A1(\design_top.MEM[2][3] ),
    .A2(\design_top.MEM[1][3] ),
    .A3(\design_top.MEM[0][3] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02622_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17376_ (.A0(_02625_),
    .A1(_02624_),
    .A2(_02623_),
    .A3(_02622_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02626_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17377_ (.A0(\design_top.MEM[31][2] ),
    .A1(\design_top.MEM[30][2] ),
    .A2(\design_top.MEM[29][2] ),
    .A3(\design_top.MEM[28][2] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02620_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17378_ (.A0(\design_top.MEM[27][2] ),
    .A1(\design_top.MEM[26][2] ),
    .A2(\design_top.MEM[25][2] ),
    .A3(\design_top.MEM[24][2] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02619_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17379_ (.A0(\design_top.MEM[23][2] ),
    .A1(\design_top.MEM[22][2] ),
    .A2(\design_top.MEM[21][2] ),
    .A3(\design_top.MEM[20][2] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02618_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17380_ (.A0(\design_top.MEM[19][2] ),
    .A1(\design_top.MEM[18][2] ),
    .A2(\design_top.MEM[17][2] ),
    .A3(\design_top.MEM[16][2] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02617_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17381_ (.A0(_02620_),
    .A1(_02619_),
    .A2(_02618_),
    .A3(_02617_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02621_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17382_ (.A0(\design_top.MEM[15][2] ),
    .A1(\design_top.MEM[14][2] ),
    .A2(\design_top.MEM[13][2] ),
    .A3(\design_top.MEM[12][2] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02615_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17383_ (.A0(\design_top.MEM[11][2] ),
    .A1(\design_top.MEM[10][2] ),
    .A2(\design_top.MEM[9][2] ),
    .A3(\design_top.MEM[8][2] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02614_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17384_ (.A0(\design_top.MEM[7][2] ),
    .A1(\design_top.MEM[6][2] ),
    .A2(\design_top.MEM[5][2] ),
    .A3(\design_top.MEM[4][2] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02613_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17385_ (.A0(\design_top.MEM[3][2] ),
    .A1(\design_top.MEM[2][2] ),
    .A2(\design_top.MEM[1][2] ),
    .A3(\design_top.MEM[0][2] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02612_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17386_ (.A0(_02615_),
    .A1(_02614_),
    .A2(_02613_),
    .A3(_02612_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02616_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17387_ (.A0(\design_top.MEM[31][1] ),
    .A1(\design_top.MEM[30][1] ),
    .A2(\design_top.MEM[29][1] ),
    .A3(\design_top.MEM[28][1] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02610_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17388_ (.A0(\design_top.MEM[27][1] ),
    .A1(\design_top.MEM[26][1] ),
    .A2(\design_top.MEM[25][1] ),
    .A3(\design_top.MEM[24][1] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02609_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17389_ (.A0(\design_top.MEM[23][1] ),
    .A1(\design_top.MEM[22][1] ),
    .A2(\design_top.MEM[21][1] ),
    .A3(\design_top.MEM[20][1] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02608_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17390_ (.A0(\design_top.MEM[19][1] ),
    .A1(\design_top.MEM[18][1] ),
    .A2(\design_top.MEM[17][1] ),
    .A3(\design_top.MEM[16][1] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02607_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17391_ (.A0(_02610_),
    .A1(_02609_),
    .A2(_02608_),
    .A3(_02607_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02611_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17392_ (.A0(\design_top.MEM[15][1] ),
    .A1(\design_top.MEM[14][1] ),
    .A2(\design_top.MEM[13][1] ),
    .A3(\design_top.MEM[12][1] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02605_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17393_ (.A0(\design_top.MEM[11][1] ),
    .A1(\design_top.MEM[10][1] ),
    .A2(\design_top.MEM[9][1] ),
    .A3(\design_top.MEM[8][1] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02604_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17394_ (.A0(\design_top.MEM[7][1] ),
    .A1(\design_top.MEM[6][1] ),
    .A2(\design_top.MEM[5][1] ),
    .A3(\design_top.MEM[4][1] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02603_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17395_ (.A0(\design_top.MEM[3][1] ),
    .A1(\design_top.MEM[2][1] ),
    .A2(\design_top.MEM[1][1] ),
    .A3(\design_top.MEM[0][1] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02602_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17396_ (.A0(_02605_),
    .A1(_02604_),
    .A2(_02603_),
    .A3(_02602_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02606_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17397_ (.A0(\design_top.MEM[31][0] ),
    .A1(\design_top.MEM[30][0] ),
    .A2(\design_top.MEM[29][0] ),
    .A3(\design_top.MEM[28][0] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02600_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17398_ (.A0(\design_top.MEM[27][0] ),
    .A1(\design_top.MEM[26][0] ),
    .A2(\design_top.MEM[25][0] ),
    .A3(\design_top.MEM[24][0] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02599_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17399_ (.A0(\design_top.MEM[23][0] ),
    .A1(\design_top.MEM[22][0] ),
    .A2(\design_top.MEM[21][0] ),
    .A3(\design_top.MEM[20][0] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02598_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17400_ (.A0(\design_top.MEM[19][0] ),
    .A1(\design_top.MEM[18][0] ),
    .A2(\design_top.MEM[17][0] ),
    .A3(\design_top.MEM[16][0] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02597_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17401_ (.A0(_02600_),
    .A1(_02599_),
    .A2(_02598_),
    .A3(_02597_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02601_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17402_ (.A0(\design_top.MEM[15][0] ),
    .A1(\design_top.MEM[14][0] ),
    .A2(\design_top.MEM[13][0] ),
    .A3(\design_top.MEM[12][0] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02595_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17403_ (.A0(\design_top.MEM[11][0] ),
    .A1(\design_top.MEM[10][0] ),
    .A2(\design_top.MEM[9][0] ),
    .A3(\design_top.MEM[8][0] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02594_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17404_ (.A0(\design_top.MEM[7][0] ),
    .A1(\design_top.MEM[6][0] ),
    .A2(\design_top.MEM[5][0] ),
    .A3(\design_top.MEM[4][0] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02593_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17405_ (.A0(\design_top.MEM[3][0] ),
    .A1(\design_top.MEM[2][0] ),
    .A2(\design_top.MEM[1][0] ),
    .A3(\design_top.MEM[0][0] ),
    .S0(_00810_),
    .S1(_00820_),
    .X(_02592_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux4_1 _17406_ (.A0(_02595_),
    .A1(_02594_),
    .A2(_02593_),
    .A3(_02592_),
    .S0(_01333_),
    .S1(_01335_),
    .X(_02596_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17407_ (.D(_00046_),
    .Q(\design_top.core0.XRES ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17408_ (.D(io_in[1]),
    .Q(\design_top.uart0.UART_RXDFF[0] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17409_ (.D(\design_top.uart0.UART_RXDFF[0] ),
    .Q(\design_top.uart0.UART_RXDFF[1] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17410_ (.D(\design_top.uart0.UART_RXDFF[1] ),
    .Q(\design_top.uart0.UART_RXDFF[2] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17411_ (.D(\design_top.XRES_reg ),
    .Q(\design_top.XRES ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17412_ (.D(io_in[0]),
    .Q(\design_top.XRES_reg ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17413_ (.D(\design_top.HLT ),
    .Q(\design_top.HLT2 ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17414_ (.D(\design_top.DADDR[2] ),
    .Q(\design_top.XADDR[2] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17415_ (.D(\design_top.DADDR[3] ),
    .Q(\design_top.XADDR[3] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17416_ (.D(\design_top.DADDR[31] ),
    .Q(\design_top.XADDR[31] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17417_ (.D(_00109_),
    .Q(\design_top.RAMFF[0] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17418_ (.D(_00120_),
    .Q(\design_top.RAMFF[1] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17419_ (.D(_00131_),
    .Q(\design_top.RAMFF[2] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17420_ (.D(_00134_),
    .Q(\design_top.RAMFF[3] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17421_ (.D(_00135_),
    .Q(\design_top.RAMFF[4] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17422_ (.D(_00136_),
    .Q(\design_top.RAMFF[5] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17423_ (.D(_00137_),
    .Q(\design_top.RAMFF[6] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17424_ (.D(_00138_),
    .Q(\design_top.RAMFF[7] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17425_ (.D(_00139_),
    .Q(\design_top.RAMFF[8] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17426_ (.D(_00140_),
    .Q(\design_top.RAMFF[9] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17427_ (.D(_00110_),
    .Q(\design_top.RAMFF[10] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17428_ (.D(_00111_),
    .Q(\design_top.RAMFF[11] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17429_ (.D(_00112_),
    .Q(\design_top.RAMFF[12] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17430_ (.D(_00113_),
    .Q(\design_top.RAMFF[13] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17431_ (.D(_00114_),
    .Q(\design_top.RAMFF[14] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17432_ (.D(_00115_),
    .Q(\design_top.RAMFF[15] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17433_ (.D(_00116_),
    .Q(\design_top.RAMFF[16] ),
    .CLK(clknet_leaf_270_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17434_ (.D(_00117_),
    .Q(\design_top.RAMFF[17] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17435_ (.D(_00118_),
    .Q(\design_top.RAMFF[18] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17436_ (.D(_00119_),
    .Q(\design_top.RAMFF[19] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17437_ (.D(_00121_),
    .Q(\design_top.RAMFF[20] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17438_ (.D(_00122_),
    .Q(\design_top.RAMFF[21] ),
    .CLK(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17439_ (.D(_00123_),
    .Q(\design_top.RAMFF[22] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17440_ (.D(_00124_),
    .Q(\design_top.RAMFF[23] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17441_ (.D(_00125_),
    .Q(\design_top.RAMFF[24] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17442_ (.D(_00126_),
    .Q(\design_top.RAMFF[25] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17443_ (.D(_00127_),
    .Q(\design_top.RAMFF[26] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17444_ (.D(_00128_),
    .Q(\design_top.RAMFF[27] ),
    .CLK(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17445_ (.D(_00129_),
    .Q(\design_top.RAMFF[28] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17446_ (.D(_00130_),
    .Q(\design_top.RAMFF[29] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17447_ (.D(_00132_),
    .Q(\design_top.RAMFF[30] ),
    .CLK(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17448_ (.D(_00133_),
    .Q(\design_top.RAMFF[31] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17449_ (.D(_00141_),
    .Q(\design_top.ROMFF[0] ),
    .CLK(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17450_ (.D(_00152_),
    .Q(\design_top.ROMFF[1] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17451_ (.D(_00163_),
    .Q(\design_top.ROMFF[2] ),
    .CLK(clknet_leaf_264_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17452_ (.D(_00166_),
    .Q(\design_top.ROMFF[3] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17453_ (.D(_00167_),
    .Q(\design_top.ROMFF[4] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17454_ (.D(_00168_),
    .Q(\design_top.ROMFF[5] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17455_ (.D(_00169_),
    .Q(\design_top.ROMFF[6] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17456_ (.D(_00170_),
    .Q(\design_top.ROMFF[7] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17457_ (.D(_00171_),
    .Q(\design_top.ROMFF[8] ),
    .CLK(clknet_leaf_271_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17458_ (.D(_00172_),
    .Q(\design_top.ROMFF[9] ),
    .CLK(clknet_leaf_290_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17459_ (.D(_00142_),
    .Q(\design_top.ROMFF[10] ),
    .CLK(clknet_leaf_270_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17460_ (.D(_00143_),
    .Q(\design_top.ROMFF[11] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17461_ (.D(_00144_),
    .Q(\design_top.ROMFF[12] ),
    .CLK(clknet_leaf_298_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17462_ (.D(_00145_),
    .Q(\design_top.ROMFF[13] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17463_ (.D(_00146_),
    .Q(\design_top.ROMFF[14] ),
    .CLK(clknet_leaf_298_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17464_ (.D(_00147_),
    .Q(\design_top.ROMFF[15] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17465_ (.D(_00148_),
    .Q(\design_top.ROMFF[16] ),
    .CLK(clknet_leaf_270_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17466_ (.D(_00149_),
    .Q(\design_top.ROMFF[17] ),
    .CLK(clknet_leaf_270_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17467_ (.D(_00150_),
    .Q(\design_top.ROMFF[18] ),
    .CLK(clknet_leaf_264_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17468_ (.D(_00151_),
    .Q(\design_top.ROMFF[19] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17469_ (.D(_00153_),
    .Q(\design_top.ROMFF[20] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17470_ (.D(_00154_),
    .Q(\design_top.ROMFF[21] ),
    .CLK(clknet_leaf_272_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17471_ (.D(_00155_),
    .Q(\design_top.ROMFF[22] ),
    .CLK(clknet_leaf_272_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17472_ (.D(_00156_),
    .Q(\design_top.ROMFF[23] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17473_ (.D(_00157_),
    .Q(\design_top.ROMFF[24] ),
    .CLK(clknet_leaf_286_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17474_ (.D(_00158_),
    .Q(\design_top.ROMFF[25] ),
    .CLK(clknet_leaf_271_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17475_ (.D(_00159_),
    .Q(\design_top.ROMFF[26] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17476_ (.D(_00160_),
    .Q(\design_top.ROMFF[27] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17477_ (.D(_00161_),
    .Q(\design_top.ROMFF[28] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17478_ (.D(_00162_),
    .Q(\design_top.ROMFF[29] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17479_ (.D(_00164_),
    .Q(\design_top.ROMFF[30] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17480_ (.D(_00165_),
    .Q(\design_top.ROMFF[31] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17481_ (.D(_03059_),
    .Q(\design_top.core0.REG2[9][0] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17482_ (.D(_03060_),
    .Q(\design_top.core0.REG2[9][1] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17483_ (.D(_03061_),
    .Q(\design_top.core0.REG2[9][2] ),
    .CLK(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17484_ (.D(_03062_),
    .Q(\design_top.core0.REG2[9][3] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17485_ (.D(_03063_),
    .Q(\design_top.core0.REG2[9][4] ),
    .CLK(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17486_ (.D(_03064_),
    .Q(\design_top.core0.REG2[9][5] ),
    .CLK(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17487_ (.D(_03065_),
    .Q(\design_top.core0.REG2[9][6] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17488_ (.D(_03066_),
    .Q(\design_top.core0.REG2[9][7] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17489_ (.D(_03067_),
    .Q(\design_top.core0.REG2[9][8] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17490_ (.D(_03068_),
    .Q(\design_top.core0.REG2[9][9] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17491_ (.D(_03069_),
    .Q(\design_top.core0.REG2[9][10] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17492_ (.D(_03070_),
    .Q(\design_top.core0.REG2[9][11] ),
    .CLK(clknet_leaf_76_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17493_ (.D(_03071_),
    .Q(\design_top.core0.REG2[9][12] ),
    .CLK(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17494_ (.D(_03072_),
    .Q(\design_top.core0.REG2[9][13] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17495_ (.D(_03073_),
    .Q(\design_top.core0.REG2[9][14] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17496_ (.D(_03074_),
    .Q(\design_top.core0.REG2[9][15] ),
    .CLK(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17497_ (.D(_03075_),
    .Q(\design_top.core0.REG2[9][16] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17498_ (.D(_03076_),
    .Q(\design_top.core0.REG2[9][17] ),
    .CLK(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17499_ (.D(_03077_),
    .Q(\design_top.core0.REG2[9][18] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17500_ (.D(_03078_),
    .Q(\design_top.core0.REG2[9][19] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17501_ (.D(_03079_),
    .Q(\design_top.core0.REG2[9][20] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17502_ (.D(_03080_),
    .Q(\design_top.core0.REG2[9][21] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17503_ (.D(_03081_),
    .Q(\design_top.core0.REG2[9][22] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17504_ (.D(_03082_),
    .Q(\design_top.core0.REG2[9][23] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17505_ (.D(_03083_),
    .Q(\design_top.core0.REG2[9][24] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17506_ (.D(_03084_),
    .Q(\design_top.core0.REG2[9][25] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17507_ (.D(_03085_),
    .Q(\design_top.core0.REG2[9][26] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17508_ (.D(_03086_),
    .Q(\design_top.core0.REG2[9][27] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17509_ (.D(_03087_),
    .Q(\design_top.core0.REG2[9][28] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17510_ (.D(_03088_),
    .Q(\design_top.core0.REG2[9][29] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17511_ (.D(_03089_),
    .Q(\design_top.core0.REG2[9][30] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17512_ (.D(_03090_),
    .Q(\design_top.core0.REG2[9][31] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17513_ (.D(_03091_),
    .Q(\design_top.core0.NXPC[0] ),
    .CLK(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17514_ (.D(_03092_),
    .Q(\design_top.core0.NXPC[1] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17515_ (.D(_03093_),
    .Q(\design_top.core0.NXPC[2] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17516_ (.D(_03094_),
    .Q(\design_top.core0.NXPC[3] ),
    .CLK(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17517_ (.D(_03095_),
    .Q(\design_top.core0.NXPC[4] ),
    .CLK(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17518_ (.D(_03096_),
    .Q(\design_top.core0.NXPC[5] ),
    .CLK(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17519_ (.D(_03097_),
    .Q(\design_top.core0.NXPC[6] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17520_ (.D(_03098_),
    .Q(\design_top.core0.NXPC[7] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17521_ (.D(_03099_),
    .Q(\design_top.core0.NXPC[8] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17522_ (.D(_03100_),
    .Q(\design_top.core0.NXPC[9] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17523_ (.D(_03101_),
    .Q(\design_top.core0.NXPC[10] ),
    .CLK(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17524_ (.D(_03102_),
    .Q(\design_top.core0.NXPC[11] ),
    .CLK(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17525_ (.D(_03103_),
    .Q(\design_top.core0.NXPC[12] ),
    .CLK(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17526_ (.D(_03104_),
    .Q(\design_top.core0.NXPC[13] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17527_ (.D(_03105_),
    .Q(\design_top.core0.NXPC[14] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17528_ (.D(_03106_),
    .Q(\design_top.core0.NXPC[15] ),
    .CLK(clknet_leaf_172_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17529_ (.D(_03107_),
    .Q(\design_top.core0.NXPC[16] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17530_ (.D(_03108_),
    .Q(\design_top.core0.NXPC[17] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17531_ (.D(_03109_),
    .Q(\design_top.core0.NXPC[18] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17532_ (.D(_03110_),
    .Q(\design_top.core0.NXPC[19] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17533_ (.D(_03111_),
    .Q(\design_top.core0.NXPC[20] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17534_ (.D(_03112_),
    .Q(\design_top.core0.NXPC[21] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17535_ (.D(_03113_),
    .Q(\design_top.core0.NXPC[22] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17536_ (.D(_03114_),
    .Q(\design_top.core0.NXPC[23] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17537_ (.D(_03115_),
    .Q(\design_top.core0.NXPC[24] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17538_ (.D(_03116_),
    .Q(\design_top.core0.NXPC[25] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17539_ (.D(_03117_),
    .Q(\design_top.core0.NXPC[26] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17540_ (.D(_03118_),
    .Q(\design_top.core0.NXPC[27] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17541_ (.D(_03119_),
    .Q(\design_top.core0.NXPC[28] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17542_ (.D(_03120_),
    .Q(\design_top.core0.NXPC[29] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17543_ (.D(_03121_),
    .Q(\design_top.core0.NXPC[30] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17544_ (.D(_03122_),
    .Q(\design_top.core0.NXPC[31] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17545_ (.D(_03123_),
    .Q(\design_top.MEM[12][0] ),
    .CLK(clknet_leaf_250_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17546_ (.D(_03124_),
    .Q(\design_top.MEM[12][1] ),
    .CLK(clknet_leaf_250_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17547_ (.D(_03125_),
    .Q(\design_top.MEM[12][2] ),
    .CLK(clknet_leaf_246_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17548_ (.D(_03126_),
    .Q(\design_top.MEM[12][3] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17549_ (.D(_03127_),
    .Q(\design_top.MEM[12][4] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17550_ (.D(_03128_),
    .Q(\design_top.MEM[12][5] ),
    .CLK(clknet_leaf_244_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17551_ (.D(_03129_),
    .Q(\design_top.MEM[12][6] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17552_ (.D(_03130_),
    .Q(\design_top.MEM[12][7] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17553_ (.D(_03131_),
    .Q(\design_top.core0.PC[0] ),
    .CLK(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17554_ (.D(_03132_),
    .Q(\design_top.core0.PC[1] ),
    .CLK(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17555_ (.D(_03133_),
    .Q(\design_top.core0.PC[2] ),
    .CLK(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17556_ (.D(_03134_),
    .Q(\design_top.core0.PC[3] ),
    .CLK(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17557_ (.D(_03135_),
    .Q(\design_top.core0.PC[4] ),
    .CLK(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17558_ (.D(_03136_),
    .Q(\design_top.core0.PC[5] ),
    .CLK(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17559_ (.D(_03137_),
    .Q(\design_top.core0.PC[6] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17560_ (.D(_03138_),
    .Q(\design_top.core0.PC[7] ),
    .CLK(clknet_5_27_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17561_ (.D(_03139_),
    .Q(\design_top.core0.PC[8] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17562_ (.D(_03140_),
    .Q(\design_top.core0.PC[9] ),
    .CLK(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17563_ (.D(_03141_),
    .Q(\design_top.core0.PC[10] ),
    .CLK(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17564_ (.D(_03142_),
    .Q(\design_top.core0.PC[11] ),
    .CLK(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17565_ (.D(_03143_),
    .Q(\design_top.core0.PC[12] ),
    .CLK(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17566_ (.D(_03144_),
    .Q(\design_top.core0.PC[13] ),
    .CLK(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17567_ (.D(_03145_),
    .Q(\design_top.core0.PC[14] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17568_ (.D(_03146_),
    .Q(\design_top.core0.PC[15] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17569_ (.D(_03147_),
    .Q(\design_top.core0.PC[16] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17570_ (.D(_03148_),
    .Q(\design_top.core0.PC[17] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17571_ (.D(_03149_),
    .Q(\design_top.core0.PC[18] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17572_ (.D(_03150_),
    .Q(\design_top.core0.PC[19] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17573_ (.D(_03151_),
    .Q(\design_top.core0.PC[20] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17574_ (.D(_03152_),
    .Q(\design_top.core0.PC[21] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17575_ (.D(_03153_),
    .Q(\design_top.core0.PC[22] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17576_ (.D(_03154_),
    .Q(\design_top.core0.PC[23] ),
    .CLK(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17577_ (.D(_03155_),
    .Q(\design_top.core0.PC[24] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17578_ (.D(_03156_),
    .Q(\design_top.core0.PC[25] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17579_ (.D(_03157_),
    .Q(\design_top.core0.PC[26] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17580_ (.D(_03158_),
    .Q(\design_top.core0.PC[27] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17581_ (.D(_03159_),
    .Q(\design_top.core0.PC[28] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17582_ (.D(_03160_),
    .Q(\design_top.core0.PC[29] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17583_ (.D(_03161_),
    .Q(\design_top.core0.PC[30] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17584_ (.D(_03162_),
    .Q(\design_top.core0.PC[31] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17585_ (.D(_03163_),
    .Q(\design_top.uart0.UART_RFIFO[0] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17586_ (.D(_03164_),
    .Q(\design_top.uart0.UART_RFIFO[1] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17587_ (.D(_03165_),
    .Q(\design_top.uart0.UART_RFIFO[2] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17588_ (.D(_03166_),
    .Q(\design_top.uart0.UART_RFIFO[3] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17589_ (.D(_03167_),
    .Q(\design_top.uart0.UART_RFIFO[4] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17590_ (.D(_03168_),
    .Q(\design_top.uart0.UART_RFIFO[5] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17591_ (.D(_03169_),
    .Q(\design_top.uart0.UART_RFIFO[6] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17592_ (.D(_03170_),
    .Q(\design_top.uart0.UART_RFIFO[7] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17593_ (.D(_03171_),
    .Q(\design_top.uart0.UART_RREQ ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17594_ (.D(_03172_),
    .Q(\design_top.uart0.UART_XACK ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17595_ (.D(_03173_),
    .Q(\design_top.ROMFF2[0] ),
    .CLK(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17596_ (.D(_03174_),
    .Q(\design_top.ROMFF2[1] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17597_ (.D(_03175_),
    .Q(\design_top.ROMFF2[2] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17598_ (.D(_03176_),
    .Q(\design_top.ROMFF2[3] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17599_ (.D(_03177_),
    .Q(\design_top.ROMFF2[4] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17600_ (.D(_03178_),
    .Q(\design_top.ROMFF2[5] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17601_ (.D(_03179_),
    .Q(\design_top.ROMFF2[6] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17602_ (.D(_03180_),
    .Q(\design_top.ROMFF2[7] ),
    .CLK(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17603_ (.D(_03181_),
    .Q(\design_top.ROMFF2[8] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17604_ (.D(_03182_),
    .Q(\design_top.ROMFF2[9] ),
    .CLK(clknet_leaf_271_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17605_ (.D(_03183_),
    .Q(\design_top.ROMFF2[10] ),
    .CLK(clknet_leaf_271_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17606_ (.D(_03184_),
    .Q(\design_top.ROMFF2[11] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17607_ (.D(_03185_),
    .Q(\design_top.ROMFF2[12] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17608_ (.D(_03186_),
    .Q(\design_top.ROMFF2[13] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17609_ (.D(_03187_),
    .Q(\design_top.ROMFF2[14] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17610_ (.D(_03188_),
    .Q(\design_top.ROMFF2[15] ),
    .CLK(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17611_ (.D(_03189_),
    .Q(\design_top.ROMFF2[16] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17612_ (.D(_03190_),
    .Q(\design_top.ROMFF2[17] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17613_ (.D(_03191_),
    .Q(\design_top.ROMFF2[18] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17614_ (.D(_03192_),
    .Q(\design_top.ROMFF2[19] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17615_ (.D(_03193_),
    .Q(\design_top.ROMFF2[20] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17616_ (.D(_03194_),
    .Q(\design_top.ROMFF2[21] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17617_ (.D(_03195_),
    .Q(\design_top.ROMFF2[22] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17618_ (.D(_03196_),
    .Q(\design_top.ROMFF2[23] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17619_ (.D(_03197_),
    .Q(\design_top.ROMFF2[24] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17620_ (.D(_03198_),
    .Q(\design_top.ROMFF2[25] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17621_ (.D(_03199_),
    .Q(\design_top.ROMFF2[26] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17622_ (.D(_03200_),
    .Q(\design_top.ROMFF2[27] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17623_ (.D(_03201_),
    .Q(\design_top.ROMFF2[28] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17624_ (.D(_03202_),
    .Q(\design_top.ROMFF2[29] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17625_ (.D(_03203_),
    .Q(\design_top.ROMFF2[30] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17626_ (.D(_03204_),
    .Q(\design_top.ROMFF2[31] ),
    .CLK(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17627_ (.D(_03205_),
    .Q(io_out[8]),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17628_ (.D(_03206_),
    .Q(io_out[9]),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17629_ (.D(_03207_),
    .Q(io_out[10]),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17630_ (.D(_03208_),
    .Q(io_out[11]),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17631_ (.D(_03209_),
    .Q(\design_top.LEDFF[4] ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17632_ (.D(_03210_),
    .Q(\design_top.LEDFF[5] ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17633_ (.D(_03211_),
    .Q(\design_top.LEDFF[6] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17634_ (.D(_03212_),
    .Q(\design_top.LEDFF[7] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17635_ (.D(_03213_),
    .Q(\design_top.LEDFF[8] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17636_ (.D(_03214_),
    .Q(\design_top.LEDFF[9] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17637_ (.D(_03215_),
    .Q(\design_top.LEDFF[10] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17638_ (.D(_03216_),
    .Q(\design_top.LEDFF[11] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17639_ (.D(_03217_),
    .Q(\design_top.LEDFF[12] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17640_ (.D(_03218_),
    .Q(\design_top.LEDFF[13] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17641_ (.D(_03219_),
    .Q(\design_top.LEDFF[14] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17642_ (.D(_03220_),
    .Q(\design_top.LEDFF[15] ),
    .CLK(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17643_ (.D(_03221_),
    .Q(io_out[15]),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17644_ (.D(_03222_),
    .Q(\design_top.GPIOFF[1] ),
    .CLK(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17645_ (.D(_03223_),
    .Q(\design_top.GPIOFF[2] ),
    .CLK(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17646_ (.D(_03224_),
    .Q(\design_top.GPIOFF[3] ),
    .CLK(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17647_ (.D(_03225_),
    .Q(\design_top.GPIOFF[4] ),
    .CLK(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17648_ (.D(_03226_),
    .Q(\design_top.GPIOFF[5] ),
    .CLK(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17649_ (.D(_03227_),
    .Q(\design_top.GPIOFF[6] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17650_ (.D(_03228_),
    .Q(\design_top.GPIOFF[7] ),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17651_ (.D(_03229_),
    .Q(\design_top.GPIOFF[8] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17652_ (.D(_03230_),
    .Q(\design_top.GPIOFF[9] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17653_ (.D(_03231_),
    .Q(\design_top.GPIOFF[10] ),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17654_ (.D(_03232_),
    .Q(\design_top.GPIOFF[11] ),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17655_ (.D(_03233_),
    .Q(\design_top.GPIOFF[12] ),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17656_ (.D(_03234_),
    .Q(\design_top.GPIOFF[13] ),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17657_ (.D(_03235_),
    .Q(\design_top.GPIOFF[14] ),
    .CLK(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17658_ (.D(_03236_),
    .Q(\design_top.GPIOFF[15] ),
    .CLK(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17659_ (.D(_03237_),
    .Q(\design_top.MEM[13][0] ),
    .CLK(clknet_leaf_249_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17660_ (.D(_03238_),
    .Q(\design_top.MEM[13][1] ),
    .CLK(clknet_leaf_250_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17661_ (.D(_03239_),
    .Q(\design_top.MEM[13][2] ),
    .CLK(clknet_leaf_249_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17662_ (.D(_03240_),
    .Q(\design_top.MEM[13][3] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17663_ (.D(_03241_),
    .Q(\design_top.MEM[13][4] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17664_ (.D(_03242_),
    .Q(\design_top.MEM[13][5] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17665_ (.D(_03243_),
    .Q(\design_top.MEM[13][6] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17666_ (.D(_03244_),
    .Q(\design_top.MEM[13][7] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17667_ (.D(_03245_),
    .Q(\design_top.MEM[2][0] ),
    .CLK(clknet_leaf_251_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17668_ (.D(_03246_),
    .Q(\design_top.MEM[2][1] ),
    .CLK(clknet_leaf_251_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17669_ (.D(_03247_),
    .Q(\design_top.MEM[2][2] ),
    .CLK(clknet_leaf_248_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17670_ (.D(_03248_),
    .Q(\design_top.MEM[2][3] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17671_ (.D(_03249_),
    .Q(\design_top.MEM[2][4] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17672_ (.D(_03250_),
    .Q(\design_top.MEM[2][5] ),
    .CLK(clknet_leaf_247_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17673_ (.D(_03251_),
    .Q(\design_top.MEM[2][6] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17674_ (.D(_03252_),
    .Q(\design_top.MEM[2][7] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17675_ (.D(_03253_),
    .Q(\design_top.MEM[29][0] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17676_ (.D(_03254_),
    .Q(\design_top.MEM[29][1] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17677_ (.D(_03255_),
    .Q(\design_top.MEM[29][2] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17678_ (.D(_03256_),
    .Q(\design_top.MEM[29][3] ),
    .CLK(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17679_ (.D(_03257_),
    .Q(\design_top.MEM[29][4] ),
    .CLK(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17680_ (.D(_03258_),
    .Q(\design_top.MEM[29][5] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17681_ (.D(_03259_),
    .Q(\design_top.MEM[29][6] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17682_ (.D(_03260_),
    .Q(\design_top.MEM[29][7] ),
    .CLK(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17683_ (.D(_03261_),
    .Q(\design_top.MEM[28][0] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17684_ (.D(_03262_),
    .Q(\design_top.MEM[28][1] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17685_ (.D(_03263_),
    .Q(\design_top.MEM[28][2] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17686_ (.D(_03264_),
    .Q(\design_top.MEM[28][3] ),
    .CLK(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17687_ (.D(_03265_),
    .Q(\design_top.MEM[28][4] ),
    .CLK(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17688_ (.D(_03266_),
    .Q(\design_top.MEM[28][5] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17689_ (.D(_03267_),
    .Q(\design_top.MEM[28][6] ),
    .CLK(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17690_ (.D(_03268_),
    .Q(\design_top.MEM[28][7] ),
    .CLK(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17691_ (.D(_03269_),
    .Q(\design_top.MEM[23][0] ),
    .CLK(clknet_leaf_259_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17692_ (.D(_03270_),
    .Q(\design_top.MEM[23][1] ),
    .CLK(clknet_leaf_258_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17693_ (.D(_03271_),
    .Q(\design_top.MEM[23][2] ),
    .CLK(clknet_leaf_258_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17694_ (.D(_03272_),
    .Q(\design_top.MEM[23][3] ),
    .CLK(clknet_leaf_263_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17695_ (.D(_03273_),
    .Q(\design_top.MEM[23][4] ),
    .CLK(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17696_ (.D(_03274_),
    .Q(\design_top.MEM[23][5] ),
    .CLK(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17697_ (.D(_03275_),
    .Q(\design_top.MEM[23][6] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17698_ (.D(_03276_),
    .Q(\design_top.MEM[23][7] ),
    .CLK(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17699_ (.D(_03277_),
    .Q(\design_top.MEM[27][0] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17700_ (.D(_03278_),
    .Q(\design_top.MEM[27][1] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17701_ (.D(_03279_),
    .Q(\design_top.MEM[27][2] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17702_ (.D(_03280_),
    .Q(\design_top.MEM[27][3] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17703_ (.D(_03281_),
    .Q(\design_top.MEM[27][4] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17704_ (.D(_03282_),
    .Q(\design_top.MEM[27][5] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17705_ (.D(_03283_),
    .Q(\design_top.MEM[27][6] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17706_ (.D(_03284_),
    .Q(\design_top.MEM[27][7] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17707_ (.D(_03285_),
    .Q(\design_top.MEM[26][0] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17708_ (.D(_03286_),
    .Q(\design_top.MEM[26][1] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17709_ (.D(_03287_),
    .Q(\design_top.MEM[26][2] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17710_ (.D(_03288_),
    .Q(\design_top.MEM[26][3] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17711_ (.D(_03289_),
    .Q(\design_top.MEM[26][4] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17712_ (.D(_03290_),
    .Q(\design_top.MEM[26][5] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17713_ (.D(_03291_),
    .Q(\design_top.MEM[26][6] ),
    .CLK(clknet_leaf_260_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17714_ (.D(_03292_),
    .Q(\design_top.MEM[26][7] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17715_ (.D(_03293_),
    .Q(\design_top.MEM[25][0] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17716_ (.D(_03294_),
    .Q(\design_top.MEM[25][1] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17717_ (.D(_03295_),
    .Q(\design_top.MEM[25][2] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17718_ (.D(_03296_),
    .Q(\design_top.MEM[25][3] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17719_ (.D(_03297_),
    .Q(\design_top.MEM[25][4] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17720_ (.D(_03298_),
    .Q(\design_top.MEM[25][5] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17721_ (.D(_03299_),
    .Q(\design_top.MEM[25][6] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17722_ (.D(_03300_),
    .Q(\design_top.MEM[25][7] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17723_ (.D(_03301_),
    .Q(\design_top.MEM[24][0] ),
    .CLK(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17724_ (.D(_03302_),
    .Q(\design_top.MEM[24][1] ),
    .CLK(clknet_leaf_260_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17725_ (.D(_03303_),
    .Q(\design_top.MEM[24][2] ),
    .CLK(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17726_ (.D(_03304_),
    .Q(\design_top.MEM[24][3] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17727_ (.D(_03305_),
    .Q(\design_top.MEM[24][4] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17728_ (.D(_03306_),
    .Q(\design_top.MEM[24][5] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17729_ (.D(_03307_),
    .Q(\design_top.MEM[24][6] ),
    .CLK(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17730_ (.D(_03308_),
    .Q(\design_top.MEM[24][7] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17731_ (.D(_03309_),
    .Q(\design_top.MEM[9][0] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17732_ (.D(_03310_),
    .Q(\design_top.MEM[9][1] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17733_ (.D(_03311_),
    .Q(\design_top.MEM[9][2] ),
    .CLK(clknet_leaf_248_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17734_ (.D(_03312_),
    .Q(\design_top.MEM[9][3] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17735_ (.D(_03313_),
    .Q(\design_top.MEM[9][4] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17736_ (.D(_03314_),
    .Q(\design_top.MEM[9][5] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17737_ (.D(_03315_),
    .Q(\design_top.MEM[9][6] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17738_ (.D(_03316_),
    .Q(\design_top.MEM[9][7] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17739_ (.D(_03317_),
    .Q(\design_top.MEM[8][0] ),
    .CLK(clknet_leaf_253_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17740_ (.D(_03318_),
    .Q(\design_top.MEM[8][1] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17741_ (.D(_03319_),
    .Q(\design_top.MEM[8][2] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17742_ (.D(_03320_),
    .Q(\design_top.MEM[8][3] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17743_ (.D(_03321_),
    .Q(\design_top.MEM[8][4] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17744_ (.D(_03322_),
    .Q(\design_top.MEM[8][5] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17745_ (.D(_03323_),
    .Q(\design_top.MEM[8][6] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17746_ (.D(_03324_),
    .Q(\design_top.MEM[8][7] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17747_ (.D(_03325_),
    .Q(\design_top.core0.REG2[14][0] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17748_ (.D(_03326_),
    .Q(\design_top.core0.REG2[14][1] ),
    .CLK(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17749_ (.D(_03327_),
    .Q(\design_top.core0.REG2[14][2] ),
    .CLK(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17750_ (.D(_03328_),
    .Q(\design_top.core0.REG2[14][3] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17751_ (.D(_03329_),
    .Q(\design_top.core0.REG2[14][4] ),
    .CLK(clknet_leaf_48_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17752_ (.D(_03330_),
    .Q(\design_top.core0.REG2[14][5] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17753_ (.D(_03331_),
    .Q(\design_top.core0.REG2[14][6] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17754_ (.D(_03332_),
    .Q(\design_top.core0.REG2[14][7] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17755_ (.D(_03333_),
    .Q(\design_top.core0.REG2[14][8] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17756_ (.D(_03334_),
    .Q(\design_top.core0.REG2[14][9] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17757_ (.D(_03335_),
    .Q(\design_top.core0.REG2[14][10] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17758_ (.D(_03336_),
    .Q(\design_top.core0.REG2[14][11] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17759_ (.D(_03337_),
    .Q(\design_top.core0.REG2[14][12] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17760_ (.D(_03338_),
    .Q(\design_top.core0.REG2[14][13] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17761_ (.D(_03339_),
    .Q(\design_top.core0.REG2[14][14] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17762_ (.D(_03340_),
    .Q(\design_top.core0.REG2[14][15] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17763_ (.D(_03341_),
    .Q(\design_top.core0.REG2[14][16] ),
    .CLK(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17764_ (.D(_03342_),
    .Q(\design_top.core0.REG2[14][17] ),
    .CLK(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17765_ (.D(_03343_),
    .Q(\design_top.core0.REG2[14][18] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17766_ (.D(_03344_),
    .Q(\design_top.core0.REG2[14][19] ),
    .CLK(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17767_ (.D(_03345_),
    .Q(\design_top.core0.REG2[14][20] ),
    .CLK(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17768_ (.D(_03346_),
    .Q(\design_top.core0.REG2[14][21] ),
    .CLK(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17769_ (.D(_03347_),
    .Q(\design_top.core0.REG2[14][22] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17770_ (.D(_03348_),
    .Q(\design_top.core0.REG2[14][23] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17771_ (.D(_03349_),
    .Q(\design_top.core0.REG2[14][24] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17772_ (.D(_03350_),
    .Q(\design_top.core0.REG2[14][25] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17773_ (.D(_03351_),
    .Q(\design_top.core0.REG2[14][26] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17774_ (.D(_03352_),
    .Q(\design_top.core0.REG2[14][27] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17775_ (.D(_03353_),
    .Q(\design_top.core0.REG2[14][28] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17776_ (.D(_03354_),
    .Q(\design_top.core0.REG2[14][29] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17777_ (.D(_03355_),
    .Q(\design_top.core0.REG2[14][30] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17778_ (.D(_03356_),
    .Q(\design_top.core0.REG2[14][31] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17779_ (.D(_03357_),
    .Q(\design_top.core0.REG2[13][0] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17780_ (.D(_03358_),
    .Q(\design_top.core0.REG2[13][1] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17781_ (.D(_03359_),
    .Q(\design_top.core0.REG2[13][2] ),
    .CLK(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17782_ (.D(_03360_),
    .Q(\design_top.core0.REG2[13][3] ),
    .CLK(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17783_ (.D(_03361_),
    .Q(\design_top.core0.REG2[13][4] ),
    .CLK(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17784_ (.D(_03362_),
    .Q(\design_top.core0.REG2[13][5] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17785_ (.D(_03363_),
    .Q(\design_top.core0.REG2[13][6] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17786_ (.D(_03364_),
    .Q(\design_top.core0.REG2[13][7] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17787_ (.D(_03365_),
    .Q(\design_top.core0.REG2[13][8] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17788_ (.D(_03366_),
    .Q(\design_top.core0.REG2[13][9] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17789_ (.D(_03367_),
    .Q(\design_top.core0.REG2[13][10] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17790_ (.D(_03368_),
    .Q(\design_top.core0.REG2[13][11] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17791_ (.D(_03369_),
    .Q(\design_top.core0.REG2[13][12] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17792_ (.D(_03370_),
    .Q(\design_top.core0.REG2[13][13] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17793_ (.D(_03371_),
    .Q(\design_top.core0.REG2[13][14] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17794_ (.D(_03372_),
    .Q(\design_top.core0.REG2[13][15] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17795_ (.D(_03373_),
    .Q(\design_top.core0.REG2[13][16] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17796_ (.D(_03374_),
    .Q(\design_top.core0.REG2[13][17] ),
    .CLK(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17797_ (.D(_03375_),
    .Q(\design_top.core0.REG2[13][18] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17798_ (.D(_03376_),
    .Q(\design_top.core0.REG2[13][19] ),
    .CLK(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17799_ (.D(_03377_),
    .Q(\design_top.core0.REG2[13][20] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17800_ (.D(_03378_),
    .Q(\design_top.core0.REG2[13][21] ),
    .CLK(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17801_ (.D(_03379_),
    .Q(\design_top.core0.REG2[13][22] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17802_ (.D(_03380_),
    .Q(\design_top.core0.REG2[13][23] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17803_ (.D(_03381_),
    .Q(\design_top.core0.REG2[13][24] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17804_ (.D(_03382_),
    .Q(\design_top.core0.REG2[13][25] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17805_ (.D(_03383_),
    .Q(\design_top.core0.REG2[13][26] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17806_ (.D(_03384_),
    .Q(\design_top.core0.REG2[13][27] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17807_ (.D(_03385_),
    .Q(\design_top.core0.REG2[13][28] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17808_ (.D(_03386_),
    .Q(\design_top.core0.REG2[13][29] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17809_ (.D(_03387_),
    .Q(\design_top.core0.REG2[13][30] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17810_ (.D(_03388_),
    .Q(\design_top.core0.REG2[13][31] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17811_ (.D(_03389_),
    .Q(\design_top.core0.REG2[12][0] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17812_ (.D(_03390_),
    .Q(\design_top.core0.REG2[12][1] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17813_ (.D(_03391_),
    .Q(\design_top.core0.REG2[12][2] ),
    .CLK(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17814_ (.D(_03392_),
    .Q(\design_top.core0.REG2[12][3] ),
    .CLK(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17815_ (.D(_03393_),
    .Q(\design_top.core0.REG2[12][4] ),
    .CLK(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17816_ (.D(_03394_),
    .Q(\design_top.core0.REG2[12][5] ),
    .CLK(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17817_ (.D(_03395_),
    .Q(\design_top.core0.REG2[12][6] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17818_ (.D(_03396_),
    .Q(\design_top.core0.REG2[12][7] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17819_ (.D(_03397_),
    .Q(\design_top.core0.REG2[12][8] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17820_ (.D(_03398_),
    .Q(\design_top.core0.REG2[12][9] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17821_ (.D(_03399_),
    .Q(\design_top.core0.REG2[12][10] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17822_ (.D(_03400_),
    .Q(\design_top.core0.REG2[12][11] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17823_ (.D(_03401_),
    .Q(\design_top.core0.REG2[12][12] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17824_ (.D(_03402_),
    .Q(\design_top.core0.REG2[12][13] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17825_ (.D(_03403_),
    .Q(\design_top.core0.REG2[12][14] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17826_ (.D(_03404_),
    .Q(\design_top.core0.REG2[12][15] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17827_ (.D(_03405_),
    .Q(\design_top.core0.REG2[12][16] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17828_ (.D(_03406_),
    .Q(\design_top.core0.REG2[12][17] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17829_ (.D(_03407_),
    .Q(\design_top.core0.REG2[12][18] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17830_ (.D(_03408_),
    .Q(\design_top.core0.REG2[12][19] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17831_ (.D(_03409_),
    .Q(\design_top.core0.REG2[12][20] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17832_ (.D(_03410_),
    .Q(\design_top.core0.REG2[12][21] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17833_ (.D(_03411_),
    .Q(\design_top.core0.REG2[12][22] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17834_ (.D(_03412_),
    .Q(\design_top.core0.REG2[12][23] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17835_ (.D(_03413_),
    .Q(\design_top.core0.REG2[12][24] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17836_ (.D(_03414_),
    .Q(\design_top.core0.REG2[12][25] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17837_ (.D(_03415_),
    .Q(\design_top.core0.REG2[12][26] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17838_ (.D(_03416_),
    .Q(\design_top.core0.REG2[12][27] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17839_ (.D(_03417_),
    .Q(\design_top.core0.REG2[12][28] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17840_ (.D(_03418_),
    .Q(\design_top.core0.REG2[12][29] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17841_ (.D(_03419_),
    .Q(\design_top.core0.REG2[12][30] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17842_ (.D(_03420_),
    .Q(\design_top.core0.REG2[12][31] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17843_ (.D(_03421_),
    .Q(\design_top.core0.REG2[11][0] ),
    .CLK(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17844_ (.D(_03422_),
    .Q(\design_top.core0.REG2[11][1] ),
    .CLK(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17845_ (.D(_03423_),
    .Q(\design_top.core0.REG2[11][2] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17846_ (.D(_03424_),
    .Q(\design_top.core0.REG2[11][3] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17847_ (.D(_03425_),
    .Q(\design_top.core0.REG2[11][4] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17848_ (.D(_03426_),
    .Q(\design_top.core0.REG2[11][5] ),
    .CLK(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17849_ (.D(_03427_),
    .Q(\design_top.core0.REG2[11][6] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17850_ (.D(_03428_),
    .Q(\design_top.core0.REG2[11][7] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17851_ (.D(_03429_),
    .Q(\design_top.core0.REG2[11][8] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17852_ (.D(_03430_),
    .Q(\design_top.core0.REG2[11][9] ),
    .CLK(clknet_leaf_76_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17853_ (.D(_03431_),
    .Q(\design_top.core0.REG2[11][10] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17854_ (.D(_03432_),
    .Q(\design_top.core0.REG2[11][11] ),
    .CLK(clknet_leaf_76_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17855_ (.D(_03433_),
    .Q(\design_top.core0.REG2[11][12] ),
    .CLK(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17856_ (.D(_03434_),
    .Q(\design_top.core0.REG2[11][13] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17857_ (.D(_03435_),
    .Q(\design_top.core0.REG2[11][14] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17858_ (.D(_03436_),
    .Q(\design_top.core0.REG2[11][15] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17859_ (.D(_03437_),
    .Q(\design_top.core0.REG2[11][16] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17860_ (.D(_03438_),
    .Q(\design_top.core0.REG2[11][17] ),
    .CLK(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17861_ (.D(_03439_),
    .Q(\design_top.core0.REG2[11][18] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17862_ (.D(_03440_),
    .Q(\design_top.core0.REG2[11][19] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17863_ (.D(_03441_),
    .Q(\design_top.core0.REG2[11][20] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17864_ (.D(_03442_),
    .Q(\design_top.core0.REG2[11][21] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17865_ (.D(_03443_),
    .Q(\design_top.core0.REG2[11][22] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17866_ (.D(_03444_),
    .Q(\design_top.core0.REG2[11][23] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17867_ (.D(_03445_),
    .Q(\design_top.core0.REG2[11][24] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17868_ (.D(_03446_),
    .Q(\design_top.core0.REG2[11][25] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17869_ (.D(_03447_),
    .Q(\design_top.core0.REG2[11][26] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17870_ (.D(_03448_),
    .Q(\design_top.core0.REG2[11][27] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17871_ (.D(_03449_),
    .Q(\design_top.core0.REG2[11][28] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17872_ (.D(_03450_),
    .Q(\design_top.core0.REG2[11][29] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17873_ (.D(_03451_),
    .Q(\design_top.core0.REG2[11][30] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17874_ (.D(_03452_),
    .Q(\design_top.core0.REG2[11][31] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17875_ (.D(_03453_),
    .Q(\design_top.core0.REG2[10][0] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17876_ (.D(_03454_),
    .Q(\design_top.core0.REG2[10][1] ),
    .CLK(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17877_ (.D(_03455_),
    .Q(\design_top.core0.REG2[10][2] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17878_ (.D(_03456_),
    .Q(\design_top.core0.REG2[10][3] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17879_ (.D(_03457_),
    .Q(\design_top.core0.REG2[10][4] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17880_ (.D(_03458_),
    .Q(\design_top.core0.REG2[10][5] ),
    .CLK(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17881_ (.D(_03459_),
    .Q(\design_top.core0.REG2[10][6] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17882_ (.D(_03460_),
    .Q(\design_top.core0.REG2[10][7] ),
    .CLK(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17883_ (.D(_03461_),
    .Q(\design_top.core0.REG2[10][8] ),
    .CLK(clknet_leaf_76_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17884_ (.D(_03462_),
    .Q(\design_top.core0.REG2[10][9] ),
    .CLK(clknet_leaf_76_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17885_ (.D(_03463_),
    .Q(\design_top.core0.REG2[10][10] ),
    .CLK(clknet_leaf_79_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17886_ (.D(_03464_),
    .Q(\design_top.core0.REG2[10][11] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17887_ (.D(_03465_),
    .Q(\design_top.core0.REG2[10][12] ),
    .CLK(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17888_ (.D(_03466_),
    .Q(\design_top.core0.REG2[10][13] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17889_ (.D(_03467_),
    .Q(\design_top.core0.REG2[10][14] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17890_ (.D(_03468_),
    .Q(\design_top.core0.REG2[10][15] ),
    .CLK(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17891_ (.D(_03469_),
    .Q(\design_top.core0.REG2[10][16] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17892_ (.D(_03470_),
    .Q(\design_top.core0.REG2[10][17] ),
    .CLK(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17893_ (.D(_03471_),
    .Q(\design_top.core0.REG2[10][18] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17894_ (.D(_03472_),
    .Q(\design_top.core0.REG2[10][19] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17895_ (.D(_03473_),
    .Q(\design_top.core0.REG2[10][20] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17896_ (.D(_03474_),
    .Q(\design_top.core0.REG2[10][21] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17897_ (.D(_03475_),
    .Q(\design_top.core0.REG2[10][22] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17898_ (.D(_03476_),
    .Q(\design_top.core0.REG2[10][23] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17899_ (.D(_03477_),
    .Q(\design_top.core0.REG2[10][24] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17900_ (.D(_03478_),
    .Q(\design_top.core0.REG2[10][25] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17901_ (.D(_03479_),
    .Q(\design_top.core0.REG2[10][26] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17902_ (.D(_03480_),
    .Q(\design_top.core0.REG2[10][27] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17903_ (.D(_03481_),
    .Q(\design_top.core0.REG2[10][28] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17904_ (.D(_03482_),
    .Q(\design_top.core0.REG2[10][29] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17905_ (.D(_03483_),
    .Q(\design_top.core0.REG2[10][30] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17906_ (.D(_03484_),
    .Q(\design_top.core0.REG2[10][31] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17907_ (.D(_03485_),
    .Q(\design_top.core0.REG2[0][0] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17908_ (.D(_03486_),
    .Q(\design_top.core0.REG2[0][1] ),
    .CLK(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17909_ (.D(_03487_),
    .Q(\design_top.core0.REG2[0][2] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17910_ (.D(_03488_),
    .Q(\design_top.core0.REG2[0][3] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17911_ (.D(_03489_),
    .Q(\design_top.core0.REG2[0][4] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17912_ (.D(_03490_),
    .Q(\design_top.core0.REG2[0][5] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17913_ (.D(_03491_),
    .Q(\design_top.core0.REG2[0][6] ),
    .CLK(clknet_leaf_79_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17914_ (.D(_03492_),
    .Q(\design_top.core0.REG2[0][7] ),
    .CLK(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17915_ (.D(_03493_),
    .Q(\design_top.core0.REG2[0][8] ),
    .CLK(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17916_ (.D(_03494_),
    .Q(\design_top.core0.REG2[0][9] ),
    .CLK(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17917_ (.D(_03495_),
    .Q(\design_top.core0.REG2[0][10] ),
    .CLK(clknet_leaf_79_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17918_ (.D(_03496_),
    .Q(\design_top.core0.REG2[0][11] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17919_ (.D(_03497_),
    .Q(\design_top.core0.REG2[0][12] ),
    .CLK(clknet_leaf_84_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17920_ (.D(_03498_),
    .Q(\design_top.core0.REG2[0][13] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17921_ (.D(_03499_),
    .Q(\design_top.core0.REG2[0][14] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17922_ (.D(_03500_),
    .Q(\design_top.core0.REG2[0][15] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17923_ (.D(_03501_),
    .Q(\design_top.core0.REG2[0][16] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17924_ (.D(_03502_),
    .Q(\design_top.core0.REG2[0][17] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17925_ (.D(_03503_),
    .Q(\design_top.core0.REG2[0][18] ),
    .CLK(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17926_ (.D(_03504_),
    .Q(\design_top.core0.REG2[0][19] ),
    .CLK(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17927_ (.D(_03505_),
    .Q(\design_top.core0.REG2[0][20] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17928_ (.D(_03506_),
    .Q(\design_top.core0.REG2[0][21] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17929_ (.D(_03507_),
    .Q(\design_top.core0.REG2[0][22] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17930_ (.D(_03508_),
    .Q(\design_top.core0.REG2[0][23] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17931_ (.D(_03509_),
    .Q(\design_top.core0.REG2[0][24] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17932_ (.D(_03510_),
    .Q(\design_top.core0.REG2[0][25] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17933_ (.D(_03511_),
    .Q(\design_top.core0.REG2[0][26] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17934_ (.D(_03512_),
    .Q(\design_top.core0.REG2[0][27] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17935_ (.D(_03513_),
    .Q(\design_top.core0.REG2[0][28] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17936_ (.D(_03514_),
    .Q(\design_top.core0.REG2[0][29] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17937_ (.D(_03515_),
    .Q(\design_top.core0.REG2[0][30] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17938_ (.D(_03516_),
    .Q(\design_top.core0.REG2[0][31] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17939_ (.D(_03517_),
    .Q(\design_top.MEM[22][0] ),
    .CLK(clknet_leaf_258_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17940_ (.D(_03518_),
    .Q(\design_top.MEM[22][1] ),
    .CLK(clknet_leaf_258_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17941_ (.D(_03519_),
    .Q(\design_top.MEM[22][2] ),
    .CLK(clknet_leaf_256_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17942_ (.D(_03520_),
    .Q(\design_top.MEM[22][3] ),
    .CLK(clknet_leaf_262_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17943_ (.D(_03521_),
    .Q(\design_top.MEM[22][4] ),
    .CLK(clknet_leaf_263_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17944_ (.D(_03522_),
    .Q(\design_top.MEM[22][5] ),
    .CLK(clknet_leaf_263_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17945_ (.D(_03523_),
    .Q(\design_top.MEM[22][6] ),
    .CLK(clknet_leaf_263_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17946_ (.D(_03524_),
    .Q(\design_top.MEM[22][7] ),
    .CLK(clknet_leaf_263_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17947_ (.D(_03525_),
    .Q(\design_top.MEM[21][0] ),
    .CLK(clknet_leaf_258_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17948_ (.D(_03526_),
    .Q(\design_top.MEM[21][1] ),
    .CLK(clknet_leaf_260_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17949_ (.D(_03527_),
    .Q(\design_top.MEM[21][2] ),
    .CLK(clknet_leaf_259_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17950_ (.D(_03528_),
    .Q(\design_top.MEM[21][3] ),
    .CLK(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17951_ (.D(_03529_),
    .Q(\design_top.MEM[21][4] ),
    .CLK(clknet_leaf_270_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17952_ (.D(_03530_),
    .Q(\design_top.MEM[21][5] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17953_ (.D(_03531_),
    .Q(\design_top.MEM[21][6] ),
    .CLK(clknet_leaf_261_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17954_ (.D(_03532_),
    .Q(\design_top.MEM[21][7] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17955_ (.D(_03533_),
    .Q(\design_top.MEM[20][0] ),
    .CLK(clknet_leaf_259_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17956_ (.D(_03534_),
    .Q(\design_top.MEM[20][1] ),
    .CLK(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17957_ (.D(_03535_),
    .Q(\design_top.MEM[20][2] ),
    .CLK(clknet_leaf_260_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17958_ (.D(_03536_),
    .Q(\design_top.MEM[20][3] ),
    .CLK(clknet_leaf_264_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17959_ (.D(_03537_),
    .Q(\design_top.MEM[20][4] ),
    .CLK(clknet_leaf_264_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17960_ (.D(_03538_),
    .Q(\design_top.MEM[20][5] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17961_ (.D(_03539_),
    .Q(\design_top.MEM[20][6] ),
    .CLK(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17962_ (.D(_03540_),
    .Q(\design_top.MEM[20][7] ),
    .CLK(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17963_ (.D(_03541_),
    .Q(\design_top.core0.REG2[8][0] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17964_ (.D(_03542_),
    .Q(\design_top.core0.REG2[8][1] ),
    .CLK(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17965_ (.D(_03543_),
    .Q(\design_top.core0.REG2[8][2] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17966_ (.D(_03544_),
    .Q(\design_top.core0.REG2[8][3] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17967_ (.D(_03545_),
    .Q(\design_top.core0.REG2[8][4] ),
    .CLK(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17968_ (.D(_03546_),
    .Q(\design_top.core0.REG2[8][5] ),
    .CLK(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17969_ (.D(_03547_),
    .Q(\design_top.core0.REG2[8][6] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17970_ (.D(_03548_),
    .Q(\design_top.core0.REG2[8][7] ),
    .CLK(clknet_leaf_76_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17971_ (.D(_03549_),
    .Q(\design_top.core0.REG2[8][8] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17972_ (.D(_03550_),
    .Q(\design_top.core0.REG2[8][9] ),
    .CLK(clknet_leaf_76_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17973_ (.D(_03551_),
    .Q(\design_top.core0.REG2[8][10] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17974_ (.D(_03552_),
    .Q(\design_top.core0.REG2[8][11] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17975_ (.D(_03553_),
    .Q(\design_top.core0.REG2[8][12] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17976_ (.D(_03554_),
    .Q(\design_top.core0.REG2[8][13] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17977_ (.D(_03555_),
    .Q(\design_top.core0.REG2[8][14] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17978_ (.D(_03556_),
    .Q(\design_top.core0.REG2[8][15] ),
    .CLK(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17979_ (.D(_03557_),
    .Q(\design_top.core0.REG2[8][16] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17980_ (.D(_03558_),
    .Q(\design_top.core0.REG2[8][17] ),
    .CLK(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17981_ (.D(_03559_),
    .Q(\design_top.core0.REG2[8][18] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17982_ (.D(_03560_),
    .Q(\design_top.core0.REG2[8][19] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17983_ (.D(_03561_),
    .Q(\design_top.core0.REG2[8][20] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17984_ (.D(_03562_),
    .Q(\design_top.core0.REG2[8][21] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17985_ (.D(_03563_),
    .Q(\design_top.core0.REG2[8][22] ),
    .CLK(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17986_ (.D(_03564_),
    .Q(\design_top.core0.REG2[8][23] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17987_ (.D(_03565_),
    .Q(\design_top.core0.REG2[8][24] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17988_ (.D(_03566_),
    .Q(\design_top.core0.REG2[8][25] ),
    .CLK(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17989_ (.D(_03567_),
    .Q(\design_top.core0.REG2[8][26] ),
    .CLK(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17990_ (.D(_03568_),
    .Q(\design_top.core0.REG2[8][27] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17991_ (.D(_03569_),
    .Q(\design_top.core0.REG2[8][28] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17992_ (.D(_03570_),
    .Q(\design_top.core0.REG2[8][29] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17993_ (.D(_03571_),
    .Q(\design_top.core0.REG2[8][30] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17994_ (.D(_03572_),
    .Q(\design_top.core0.REG2[8][31] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17995_ (.D(_03573_),
    .Q(\design_top.core0.REG2[7][0] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17996_ (.D(_03574_),
    .Q(\design_top.core0.REG2[7][1] ),
    .CLK(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17997_ (.D(_03575_),
    .Q(\design_top.core0.REG2[7][2] ),
    .CLK(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17998_ (.D(_03576_),
    .Q(\design_top.core0.REG2[7][3] ),
    .CLK(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _17999_ (.D(_03577_),
    .Q(\design_top.core0.REG2[7][4] ),
    .CLK(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18000_ (.D(_03578_),
    .Q(\design_top.core0.REG2[7][5] ),
    .CLK(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18001_ (.D(_03579_),
    .Q(\design_top.core0.REG2[7][6] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18002_ (.D(_03580_),
    .Q(\design_top.core0.REG2[7][7] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18003_ (.D(_03581_),
    .Q(\design_top.core0.REG2[7][8] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18004_ (.D(_03582_),
    .Q(\design_top.core0.REG2[7][9] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18005_ (.D(_03583_),
    .Q(\design_top.core0.REG2[7][10] ),
    .CLK(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18006_ (.D(_03584_),
    .Q(\design_top.core0.REG2[7][11] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18007_ (.D(_03585_),
    .Q(\design_top.core0.REG2[7][12] ),
    .CLK(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18008_ (.D(_03586_),
    .Q(\design_top.core0.REG2[7][13] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18009_ (.D(_03587_),
    .Q(\design_top.core0.REG2[7][14] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18010_ (.D(_03588_),
    .Q(\design_top.core0.REG2[7][15] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18011_ (.D(_03589_),
    .Q(\design_top.core0.REG2[7][16] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18012_ (.D(_03590_),
    .Q(\design_top.core0.REG2[7][17] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18013_ (.D(_03591_),
    .Q(\design_top.core0.REG2[7][18] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18014_ (.D(_03592_),
    .Q(\design_top.core0.REG2[7][19] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18015_ (.D(_03593_),
    .Q(\design_top.core0.REG2[7][20] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18016_ (.D(_03594_),
    .Q(\design_top.core0.REG2[7][21] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18017_ (.D(_03595_),
    .Q(\design_top.core0.REG2[7][22] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18018_ (.D(_03596_),
    .Q(\design_top.core0.REG2[7][23] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18019_ (.D(_03597_),
    .Q(\design_top.core0.REG2[7][24] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18020_ (.D(_03598_),
    .Q(\design_top.core0.REG2[7][25] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18021_ (.D(_03599_),
    .Q(\design_top.core0.REG2[7][26] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18022_ (.D(_03600_),
    .Q(\design_top.core0.REG2[7][27] ),
    .CLK(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18023_ (.D(_03601_),
    .Q(\design_top.core0.REG2[7][28] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18024_ (.D(_03602_),
    .Q(\design_top.core0.REG2[7][29] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18025_ (.D(_03603_),
    .Q(\design_top.core0.REG2[7][30] ),
    .CLK(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18026_ (.D(_03604_),
    .Q(\design_top.core0.REG2[7][31] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18027_ (.D(_03605_),
    .Q(\design_top.core0.REG2[6][0] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18028_ (.D(_03606_),
    .Q(\design_top.core0.REG2[6][1] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18029_ (.D(_03607_),
    .Q(\design_top.core0.REG2[6][2] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18030_ (.D(_03608_),
    .Q(\design_top.core0.REG2[6][3] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18031_ (.D(_03609_),
    .Q(\design_top.core0.REG2[6][4] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18032_ (.D(_03610_),
    .Q(\design_top.core0.REG2[6][5] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18033_ (.D(_03611_),
    .Q(\design_top.core0.REG2[6][6] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18034_ (.D(_03612_),
    .Q(\design_top.core0.REG2[6][7] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18035_ (.D(_03613_),
    .Q(\design_top.core0.REG2[6][8] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18036_ (.D(_03614_),
    .Q(\design_top.core0.REG2[6][9] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18037_ (.D(_03615_),
    .Q(\design_top.core0.REG2[6][10] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18038_ (.D(_03616_),
    .Q(\design_top.core0.REG2[6][11] ),
    .CLK(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18039_ (.D(_03617_),
    .Q(\design_top.core0.REG2[6][12] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18040_ (.D(_03618_),
    .Q(\design_top.core0.REG2[6][13] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18041_ (.D(_03619_),
    .Q(\design_top.core0.REG2[6][14] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18042_ (.D(_03620_),
    .Q(\design_top.core0.REG2[6][15] ),
    .CLK(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18043_ (.D(_03621_),
    .Q(\design_top.core0.REG2[6][16] ),
    .CLK(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18044_ (.D(_03622_),
    .Q(\design_top.core0.REG2[6][17] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18045_ (.D(_03623_),
    .Q(\design_top.core0.REG2[6][18] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18046_ (.D(_03624_),
    .Q(\design_top.core0.REG2[6][19] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18047_ (.D(_03625_),
    .Q(\design_top.core0.REG2[6][20] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18048_ (.D(_03626_),
    .Q(\design_top.core0.REG2[6][21] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18049_ (.D(_03627_),
    .Q(\design_top.core0.REG2[6][22] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18050_ (.D(_03628_),
    .Q(\design_top.core0.REG2[6][23] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18051_ (.D(_03629_),
    .Q(\design_top.core0.REG2[6][24] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18052_ (.D(_03630_),
    .Q(\design_top.core0.REG2[6][25] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18053_ (.D(_03631_),
    .Q(\design_top.core0.REG2[6][26] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18054_ (.D(_03632_),
    .Q(\design_top.core0.REG2[6][27] ),
    .CLK(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18055_ (.D(_03633_),
    .Q(\design_top.core0.REG2[6][28] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18056_ (.D(_03634_),
    .Q(\design_top.core0.REG2[6][29] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18057_ (.D(_03635_),
    .Q(\design_top.core0.REG2[6][30] ),
    .CLK(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18058_ (.D(_03636_),
    .Q(\design_top.core0.REG2[6][31] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18059_ (.D(_03637_),
    .Q(\design_top.core0.REG2[5][0] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18060_ (.D(_03638_),
    .Q(\design_top.core0.REG2[5][1] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18061_ (.D(_03639_),
    .Q(\design_top.core0.REG2[5][2] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18062_ (.D(_03640_),
    .Q(\design_top.core0.REG2[5][3] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18063_ (.D(_03641_),
    .Q(\design_top.core0.REG2[5][4] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18064_ (.D(_03642_),
    .Q(\design_top.core0.REG2[5][5] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18065_ (.D(_03643_),
    .Q(\design_top.core0.REG2[5][6] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18066_ (.D(_03644_),
    .Q(\design_top.core0.REG2[5][7] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18067_ (.D(_03645_),
    .Q(\design_top.core0.REG2[5][8] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18068_ (.D(_03646_),
    .Q(\design_top.core0.REG2[5][9] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18069_ (.D(_03647_),
    .Q(\design_top.core0.REG2[5][10] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18070_ (.D(_03648_),
    .Q(\design_top.core0.REG2[5][11] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18071_ (.D(_03649_),
    .Q(\design_top.core0.REG2[5][12] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18072_ (.D(_03650_),
    .Q(\design_top.core0.REG2[5][13] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18073_ (.D(_03651_),
    .Q(\design_top.core0.REG2[5][14] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18074_ (.D(_03652_),
    .Q(\design_top.core0.REG2[5][15] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18075_ (.D(_03653_),
    .Q(\design_top.core0.REG2[5][16] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18076_ (.D(_03654_),
    .Q(\design_top.core0.REG2[5][17] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18077_ (.D(_03655_),
    .Q(\design_top.core0.REG2[5][18] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18078_ (.D(_03656_),
    .Q(\design_top.core0.REG2[5][19] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18079_ (.D(_03657_),
    .Q(\design_top.core0.REG2[5][20] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18080_ (.D(_03658_),
    .Q(\design_top.core0.REG2[5][21] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18081_ (.D(_03659_),
    .Q(\design_top.core0.REG2[5][22] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18082_ (.D(_03660_),
    .Q(\design_top.core0.REG2[5][23] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18083_ (.D(_03661_),
    .Q(\design_top.core0.REG2[5][24] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18084_ (.D(_03662_),
    .Q(\design_top.core0.REG2[5][25] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18085_ (.D(_03663_),
    .Q(\design_top.core0.REG2[5][26] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18086_ (.D(_03664_),
    .Q(\design_top.core0.REG2[5][27] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18087_ (.D(_03665_),
    .Q(\design_top.core0.REG2[5][28] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18088_ (.D(_03666_),
    .Q(\design_top.core0.REG2[5][29] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18089_ (.D(_03667_),
    .Q(\design_top.core0.REG2[5][30] ),
    .CLK(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18090_ (.D(_03668_),
    .Q(\design_top.core0.REG2[5][31] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18091_ (.D(_03669_),
    .Q(\design_top.MEM[7][0] ),
    .CLK(clknet_leaf_250_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18092_ (.D(_03670_),
    .Q(\design_top.MEM[7][1] ),
    .CLK(clknet_leaf_250_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18093_ (.D(_03671_),
    .Q(\design_top.MEM[7][2] ),
    .CLK(clknet_leaf_249_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18094_ (.D(_03672_),
    .Q(\design_top.MEM[7][3] ),
    .CLK(clknet_leaf_245_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18095_ (.D(_03673_),
    .Q(\design_top.MEM[7][4] ),
    .CLK(clknet_leaf_246_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18096_ (.D(_03674_),
    .Q(\design_top.MEM[7][5] ),
    .CLK(clknet_leaf_246_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18097_ (.D(_03675_),
    .Q(\design_top.MEM[7][6] ),
    .CLK(clknet_leaf_244_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18098_ (.D(_03676_),
    .Q(\design_top.MEM[7][7] ),
    .CLK(clknet_leaf_244_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18099_ (.D(_03677_),
    .Q(\design_top.core0.REG2[4][0] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18100_ (.D(_03678_),
    .Q(\design_top.core0.REG2[4][1] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18101_ (.D(_03679_),
    .Q(\design_top.core0.REG2[4][2] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18102_ (.D(_03680_),
    .Q(\design_top.core0.REG2[4][3] ),
    .CLK(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18103_ (.D(_03681_),
    .Q(\design_top.core0.REG2[4][4] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18104_ (.D(_03682_),
    .Q(\design_top.core0.REG2[4][5] ),
    .CLK(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18105_ (.D(_03683_),
    .Q(\design_top.core0.REG2[4][6] ),
    .CLK(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18106_ (.D(_03684_),
    .Q(\design_top.core0.REG2[4][7] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18107_ (.D(_03685_),
    .Q(\design_top.core0.REG2[4][8] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18108_ (.D(_03686_),
    .Q(\design_top.core0.REG2[4][9] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18109_ (.D(_03687_),
    .Q(\design_top.core0.REG2[4][10] ),
    .CLK(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18110_ (.D(_03688_),
    .Q(\design_top.core0.REG2[4][11] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18111_ (.D(_03689_),
    .Q(\design_top.core0.REG2[4][12] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18112_ (.D(_03690_),
    .Q(\design_top.core0.REG2[4][13] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18113_ (.D(_03691_),
    .Q(\design_top.core0.REG2[4][14] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18114_ (.D(_03692_),
    .Q(\design_top.core0.REG2[4][15] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18115_ (.D(_03693_),
    .Q(\design_top.core0.REG2[4][16] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18116_ (.D(_03694_),
    .Q(\design_top.core0.REG2[4][17] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18117_ (.D(_03695_),
    .Q(\design_top.core0.REG2[4][18] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18118_ (.D(_03696_),
    .Q(\design_top.core0.REG2[4][19] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18119_ (.D(_03697_),
    .Q(\design_top.core0.REG2[4][20] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18120_ (.D(_03698_),
    .Q(\design_top.core0.REG2[4][21] ),
    .CLK(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18121_ (.D(_03699_),
    .Q(\design_top.core0.REG2[4][22] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18122_ (.D(_03700_),
    .Q(\design_top.core0.REG2[4][23] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18123_ (.D(_03701_),
    .Q(\design_top.core0.REG2[4][24] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18124_ (.D(_03702_),
    .Q(\design_top.core0.REG2[4][25] ),
    .CLK(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18125_ (.D(_03703_),
    .Q(\design_top.core0.REG2[4][26] ),
    .CLK(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18126_ (.D(_03704_),
    .Q(\design_top.core0.REG2[4][27] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18127_ (.D(_03705_),
    .Q(\design_top.core0.REG2[4][28] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18128_ (.D(_03706_),
    .Q(\design_top.core0.REG2[4][29] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18129_ (.D(_03707_),
    .Q(\design_top.core0.REG2[4][30] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18130_ (.D(_03708_),
    .Q(\design_top.core0.REG2[4][31] ),
    .CLK(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18131_ (.D(_03709_),
    .Q(\design_top.core0.REG2[3][0] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18132_ (.D(_03710_),
    .Q(\design_top.core0.REG2[3][1] ),
    .CLK(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18133_ (.D(_03711_),
    .Q(\design_top.core0.REG2[3][2] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18134_ (.D(_03712_),
    .Q(\design_top.core0.REG2[3][3] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18135_ (.D(_03713_),
    .Q(\design_top.core0.REG2[3][4] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18136_ (.D(_03714_),
    .Q(\design_top.core0.REG2[3][5] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18137_ (.D(_03715_),
    .Q(\design_top.core0.REG2[3][6] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18138_ (.D(_03716_),
    .Q(\design_top.core0.REG2[3][7] ),
    .CLK(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18139_ (.D(_03717_),
    .Q(\design_top.core0.REG2[3][8] ),
    .CLK(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18140_ (.D(_03718_),
    .Q(\design_top.core0.REG2[3][9] ),
    .CLK(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18141_ (.D(_03719_),
    .Q(\design_top.core0.REG2[3][10] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18142_ (.D(_03720_),
    .Q(\design_top.core0.REG2[3][11] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18143_ (.D(_03721_),
    .Q(\design_top.core0.REG2[3][12] ),
    .CLK(clknet_leaf_84_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18144_ (.D(_03722_),
    .Q(\design_top.core0.REG2[3][13] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18145_ (.D(_03723_),
    .Q(\design_top.core0.REG2[3][14] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18146_ (.D(_03724_),
    .Q(\design_top.core0.REG2[3][15] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18147_ (.D(_03725_),
    .Q(\design_top.core0.REG2[3][16] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18148_ (.D(_03726_),
    .Q(\design_top.core0.REG2[3][17] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18149_ (.D(_03727_),
    .Q(\design_top.core0.REG2[3][18] ),
    .CLK(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18150_ (.D(_03728_),
    .Q(\design_top.core0.REG2[3][19] ),
    .CLK(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18151_ (.D(_03729_),
    .Q(\design_top.core0.REG2[3][20] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18152_ (.D(_03730_),
    .Q(\design_top.core0.REG2[3][21] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18153_ (.D(_03731_),
    .Q(\design_top.core0.REG2[3][22] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18154_ (.D(_03732_),
    .Q(\design_top.core0.REG2[3][23] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18155_ (.D(_03733_),
    .Q(\design_top.core0.REG2[3][24] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18156_ (.D(_03734_),
    .Q(\design_top.core0.REG2[3][25] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18157_ (.D(_03735_),
    .Q(\design_top.core0.REG2[3][26] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18158_ (.D(_03736_),
    .Q(\design_top.core0.REG2[3][27] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18159_ (.D(_03737_),
    .Q(\design_top.core0.REG2[3][28] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18160_ (.D(_03738_),
    .Q(\design_top.core0.REG2[3][29] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18161_ (.D(_03739_),
    .Q(\design_top.core0.REG2[3][30] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18162_ (.D(_03740_),
    .Q(\design_top.core0.REG2[3][31] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18163_ (.D(_03741_),
    .Q(\design_top.core0.REG2[2][0] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18164_ (.D(_03742_),
    .Q(\design_top.core0.REG2[2][1] ),
    .CLK(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18165_ (.D(_03743_),
    .Q(\design_top.core0.REG2[2][2] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18166_ (.D(_03744_),
    .Q(\design_top.core0.REG2[2][3] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18167_ (.D(_03745_),
    .Q(\design_top.core0.REG2[2][4] ),
    .CLK(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18168_ (.D(_03746_),
    .Q(\design_top.core0.REG2[2][5] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18169_ (.D(_03747_),
    .Q(\design_top.core0.REG2[2][6] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18170_ (.D(_03748_),
    .Q(\design_top.core0.REG2[2][7] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18171_ (.D(_03749_),
    .Q(\design_top.core0.REG2[2][8] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18172_ (.D(_03750_),
    .Q(\design_top.core0.REG2[2][9] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18173_ (.D(_03751_),
    .Q(\design_top.core0.REG2[2][10] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18174_ (.D(_03752_),
    .Q(\design_top.core0.REG2[2][11] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18175_ (.D(_03753_),
    .Q(\design_top.core0.REG2[2][12] ),
    .CLK(clknet_leaf_84_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18176_ (.D(_03754_),
    .Q(\design_top.core0.REG2[2][13] ),
    .CLK(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18177_ (.D(_03755_),
    .Q(\design_top.core0.REG2[2][14] ),
    .CLK(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18178_ (.D(_03756_),
    .Q(\design_top.core0.REG2[2][15] ),
    .CLK(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18179_ (.D(_03757_),
    .Q(\design_top.core0.REG2[2][16] ),
    .CLK(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18180_ (.D(_03758_),
    .Q(\design_top.core0.REG2[2][17] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18181_ (.D(_03759_),
    .Q(\design_top.core0.REG2[2][18] ),
    .CLK(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18182_ (.D(_03760_),
    .Q(\design_top.core0.REG2[2][19] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18183_ (.D(_03761_),
    .Q(\design_top.core0.REG2[2][20] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18184_ (.D(_03762_),
    .Q(\design_top.core0.REG2[2][21] ),
    .CLK(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18185_ (.D(_03763_),
    .Q(\design_top.core0.REG2[2][22] ),
    .CLK(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18186_ (.D(_03764_),
    .Q(\design_top.core0.REG2[2][23] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18187_ (.D(_03765_),
    .Q(\design_top.core0.REG2[2][24] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18188_ (.D(_03766_),
    .Q(\design_top.core0.REG2[2][25] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18189_ (.D(_03767_),
    .Q(\design_top.core0.REG2[2][26] ),
    .CLK(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18190_ (.D(_03768_),
    .Q(\design_top.core0.REG2[2][27] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18191_ (.D(_03769_),
    .Q(\design_top.core0.REG2[2][28] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18192_ (.D(_03770_),
    .Q(\design_top.core0.REG2[2][29] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18193_ (.D(_03771_),
    .Q(\design_top.core0.REG2[2][30] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18194_ (.D(_03772_),
    .Q(\design_top.core0.REG2[2][31] ),
    .CLK(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18195_ (.D(_03773_),
    .Q(\design_top.core0.REG2[1][0] ),
    .CLK(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18196_ (.D(_03774_),
    .Q(\design_top.core0.REG2[1][1] ),
    .CLK(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18197_ (.D(_03775_),
    .Q(\design_top.core0.REG2[1][2] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18198_ (.D(_03776_),
    .Q(\design_top.core0.REG2[1][3] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18199_ (.D(_03777_),
    .Q(\design_top.core0.REG2[1][4] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18200_ (.D(_03778_),
    .Q(\design_top.core0.REG2[1][5] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18201_ (.D(_03779_),
    .Q(\design_top.core0.REG2[1][6] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18202_ (.D(_03780_),
    .Q(\design_top.core0.REG2[1][7] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18203_ (.D(_03781_),
    .Q(\design_top.core0.REG2[1][8] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18204_ (.D(_03782_),
    .Q(\design_top.core0.REG2[1][9] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18205_ (.D(_03783_),
    .Q(\design_top.core0.REG2[1][10] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18206_ (.D(_03784_),
    .Q(\design_top.core0.REG2[1][11] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18207_ (.D(_03785_),
    .Q(\design_top.core0.REG2[1][12] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18208_ (.D(_03786_),
    .Q(\design_top.core0.REG2[1][13] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18209_ (.D(_03787_),
    .Q(\design_top.core0.REG2[1][14] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18210_ (.D(_03788_),
    .Q(\design_top.core0.REG2[1][15] ),
    .CLK(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18211_ (.D(_03789_),
    .Q(\design_top.core0.REG2[1][16] ),
    .CLK(clknet_5_22_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18212_ (.D(_03790_),
    .Q(\design_top.core0.REG2[1][17] ),
    .CLK(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18213_ (.D(_03791_),
    .Q(\design_top.core0.REG2[1][18] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18214_ (.D(_03792_),
    .Q(\design_top.core0.REG2[1][19] ),
    .CLK(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18215_ (.D(_03793_),
    .Q(\design_top.core0.REG2[1][20] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18216_ (.D(_03794_),
    .Q(\design_top.core0.REG2[1][21] ),
    .CLK(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18217_ (.D(_03795_),
    .Q(\design_top.core0.REG2[1][22] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18218_ (.D(_03796_),
    .Q(\design_top.core0.REG2[1][23] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18219_ (.D(_03797_),
    .Q(\design_top.core0.REG2[1][24] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18220_ (.D(_03798_),
    .Q(\design_top.core0.REG2[1][25] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18221_ (.D(_03799_),
    .Q(\design_top.core0.REG2[1][26] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18222_ (.D(_03800_),
    .Q(\design_top.core0.REG2[1][27] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18223_ (.D(_03801_),
    .Q(\design_top.core0.REG2[1][28] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18224_ (.D(_03802_),
    .Q(\design_top.core0.REG2[1][29] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18225_ (.D(_03803_),
    .Q(\design_top.core0.REG2[1][30] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18226_ (.D(_03804_),
    .Q(\design_top.core0.REG2[1][31] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18227_ (.D(_03805_),
    .Q(\design_top.core0.REG2[15][0] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18228_ (.D(_03806_),
    .Q(\design_top.core0.REG2[15][1] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18229_ (.D(_03807_),
    .Q(\design_top.core0.REG2[15][2] ),
    .CLK(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18230_ (.D(_03808_),
    .Q(\design_top.core0.REG2[15][3] ),
    .CLK(clknet_leaf_48_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18231_ (.D(_03809_),
    .Q(\design_top.core0.REG2[15][4] ),
    .CLK(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18232_ (.D(_03810_),
    .Q(\design_top.core0.REG2[15][5] ),
    .CLK(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18233_ (.D(_03811_),
    .Q(\design_top.core0.REG2[15][6] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18234_ (.D(_03812_),
    .Q(\design_top.core0.REG2[15][7] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18235_ (.D(_03813_),
    .Q(\design_top.core0.REG2[15][8] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18236_ (.D(_03814_),
    .Q(\design_top.core0.REG2[15][9] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18237_ (.D(_03815_),
    .Q(\design_top.core0.REG2[15][10] ),
    .CLK(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18238_ (.D(_03816_),
    .Q(\design_top.core0.REG2[15][11] ),
    .CLK(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18239_ (.D(_03817_),
    .Q(\design_top.core0.REG2[15][12] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18240_ (.D(_03818_),
    .Q(\design_top.core0.REG2[15][13] ),
    .CLK(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18241_ (.D(_03819_),
    .Q(\design_top.core0.REG2[15][14] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18242_ (.D(_03820_),
    .Q(\design_top.core0.REG2[15][15] ),
    .CLK(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18243_ (.D(_03821_),
    .Q(\design_top.core0.REG2[15][16] ),
    .CLK(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18244_ (.D(_03822_),
    .Q(\design_top.core0.REG2[15][17] ),
    .CLK(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18245_ (.D(_03823_),
    .Q(\design_top.core0.REG2[15][18] ),
    .CLK(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18246_ (.D(_03824_),
    .Q(\design_top.core0.REG2[15][19] ),
    .CLK(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18247_ (.D(_03825_),
    .Q(\design_top.core0.REG2[15][20] ),
    .CLK(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18248_ (.D(_03826_),
    .Q(\design_top.core0.REG2[15][21] ),
    .CLK(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18249_ (.D(_03827_),
    .Q(\design_top.core0.REG2[15][22] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18250_ (.D(_03828_),
    .Q(\design_top.core0.REG2[15][23] ),
    .CLK(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18251_ (.D(_03829_),
    .Q(\design_top.core0.REG2[15][24] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18252_ (.D(_03830_),
    .Q(\design_top.core0.REG2[15][25] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18253_ (.D(_03831_),
    .Q(\design_top.core0.REG2[15][26] ),
    .CLK(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18254_ (.D(_03832_),
    .Q(\design_top.core0.REG2[15][27] ),
    .CLK(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18255_ (.D(_03833_),
    .Q(\design_top.core0.REG2[15][28] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18256_ (.D(_03834_),
    .Q(\design_top.core0.REG2[15][29] ),
    .CLK(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18257_ (.D(_03835_),
    .Q(\design_top.core0.REG2[15][30] ),
    .CLK(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18258_ (.D(_03836_),
    .Q(\design_top.core0.REG2[15][31] ),
    .CLK(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18259_ (.D(_03837_),
    .Q(\design_top.MEM[1][0] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18260_ (.D(_03838_),
    .Q(\design_top.MEM[1][1] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18261_ (.D(_03839_),
    .Q(\design_top.MEM[1][2] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18262_ (.D(_03840_),
    .Q(\design_top.MEM[1][3] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18263_ (.D(_03841_),
    .Q(\design_top.MEM[1][4] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18264_ (.D(_03842_),
    .Q(\design_top.MEM[1][5] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18265_ (.D(_03843_),
    .Q(\design_top.MEM[1][6] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18266_ (.D(_03844_),
    .Q(\design_top.MEM[1][7] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18267_ (.D(_03845_),
    .Q(\design_top.MEM[19][0] ),
    .CLK(clknet_leaf_253_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18268_ (.D(_03846_),
    .Q(\design_top.MEM[19][1] ),
    .CLK(clknet_leaf_253_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18269_ (.D(_03847_),
    .Q(\design_top.MEM[19][2] ),
    .CLK(clknet_leaf_255_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18270_ (.D(_03848_),
    .Q(\design_top.MEM[19][3] ),
    .CLK(clknet_leaf_255_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18271_ (.D(_03849_),
    .Q(\design_top.MEM[19][4] ),
    .CLK(clknet_leaf_266_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18272_ (.D(_03850_),
    .Q(\design_top.MEM[19][5] ),
    .CLK(clknet_leaf_266_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18273_ (.D(_03851_),
    .Q(\design_top.MEM[19][6] ),
    .CLK(clknet_leaf_256_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18274_ (.D(_03852_),
    .Q(\design_top.MEM[19][7] ),
    .CLK(clknet_leaf_258_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18275_ (.D(_03853_),
    .Q(\design_top.MEM[18][0] ),
    .CLK(clknet_leaf_253_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18276_ (.D(_03854_),
    .Q(\design_top.MEM[18][1] ),
    .CLK(clknet_leaf_256_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18277_ (.D(_03855_),
    .Q(\design_top.MEM[18][2] ),
    .CLK(clknet_leaf_256_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18278_ (.D(_03856_),
    .Q(\design_top.MEM[18][3] ),
    .CLK(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18279_ (.D(_03857_),
    .Q(\design_top.MEM[18][4] ),
    .CLK(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18280_ (.D(_03858_),
    .Q(\design_top.MEM[18][5] ),
    .CLK(clknet_leaf_262_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18281_ (.D(_03859_),
    .Q(\design_top.MEM[18][6] ),
    .CLK(clknet_leaf_258_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18282_ (.D(_03860_),
    .Q(\design_top.MEM[18][7] ),
    .CLK(clknet_leaf_262_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18283_ (.D(_03861_),
    .Q(\design_top.MEM[17][0] ),
    .CLK(clknet_leaf_255_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18284_ (.D(_03862_),
    .Q(\design_top.MEM[17][1] ),
    .CLK(clknet_leaf_255_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18285_ (.D(_03863_),
    .Q(\design_top.MEM[17][2] ),
    .CLK(clknet_leaf_255_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18286_ (.D(_03864_),
    .Q(\design_top.MEM[17][3] ),
    .CLK(clknet_leaf_266_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18287_ (.D(_03865_),
    .Q(\design_top.MEM[17][4] ),
    .CLK(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18288_ (.D(_03866_),
    .Q(\design_top.MEM[17][5] ),
    .CLK(clknet_leaf_261_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18289_ (.D(_03867_),
    .Q(\design_top.MEM[17][6] ),
    .CLK(clknet_leaf_258_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18290_ (.D(_03868_),
    .Q(\design_top.MEM[17][7] ),
    .CLK(clknet_leaf_261_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18291_ (.D(_03869_),
    .Q(\design_top.MEM[16][0] ),
    .CLK(clknet_leaf_255_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18292_ (.D(_03870_),
    .Q(\design_top.MEM[16][1] ),
    .CLK(clknet_leaf_255_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18293_ (.D(_03871_),
    .Q(\design_top.MEM[16][2] ),
    .CLK(clknet_leaf_255_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18294_ (.D(_03872_),
    .Q(\design_top.MEM[16][3] ),
    .CLK(clknet_leaf_266_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18295_ (.D(_03873_),
    .Q(\design_top.MEM[16][4] ),
    .CLK(clknet_leaf_266_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18296_ (.D(_03874_),
    .Q(\design_top.MEM[16][5] ),
    .CLK(clknet_leaf_262_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18297_ (.D(_03875_),
    .Q(\design_top.MEM[16][6] ),
    .CLK(clknet_leaf_258_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18298_ (.D(_03876_),
    .Q(\design_top.MEM[16][7] ),
    .CLK(clknet_leaf_262_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18299_ (.D(_03877_),
    .Q(\design_top.MEM[15][0] ),
    .CLK(clknet_leaf_250_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18300_ (.D(_03878_),
    .Q(\design_top.MEM[15][1] ),
    .CLK(clknet_leaf_298_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18301_ (.D(_03879_),
    .Q(\design_top.MEM[15][2] ),
    .CLK(clknet_leaf_249_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18302_ (.D(_03880_),
    .Q(\design_top.MEM[15][3] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18303_ (.D(_03881_),
    .Q(\design_top.MEM[15][4] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18304_ (.D(_03882_),
    .Q(\design_top.MEM[15][5] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18305_ (.D(_03883_),
    .Q(\design_top.MEM[15][6] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18306_ (.D(_03884_),
    .Q(\design_top.MEM[15][7] ),
    .CLK(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18307_ (.D(_03885_),
    .Q(\design_top.MEM[14][0] ),
    .CLK(clknet_leaf_249_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18308_ (.D(_03886_),
    .Q(\design_top.MEM[14][1] ),
    .CLK(clknet_leaf_298_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18309_ (.D(_03887_),
    .Q(\design_top.MEM[14][2] ),
    .CLK(clknet_leaf_249_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18310_ (.D(_03888_),
    .Q(\design_top.MEM[14][3] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18311_ (.D(_03889_),
    .Q(\design_top.MEM[14][4] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18312_ (.D(_03890_),
    .Q(\design_top.MEM[14][5] ),
    .CLK(clknet_leaf_244_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18313_ (.D(_03891_),
    .Q(\design_top.MEM[14][6] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18314_ (.D(_03892_),
    .Q(\design_top.MEM[14][7] ),
    .CLK(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18315_ (.D(_03893_),
    .Q(\design_top.core0.REG1[9][0] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18316_ (.D(_03894_),
    .Q(\design_top.core0.REG1[9][1] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18317_ (.D(_03895_),
    .Q(\design_top.core0.REG1[9][2] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18318_ (.D(_03896_),
    .Q(\design_top.core0.REG1[9][3] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18319_ (.D(_03897_),
    .Q(\design_top.core0.REG1[9][4] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18320_ (.D(_03898_),
    .Q(\design_top.core0.REG1[9][5] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18321_ (.D(_03899_),
    .Q(\design_top.core0.REG1[9][6] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18322_ (.D(_03900_),
    .Q(\design_top.core0.REG1[9][7] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18323_ (.D(_03901_),
    .Q(\design_top.core0.REG1[9][8] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18324_ (.D(_03902_),
    .Q(\design_top.core0.REG1[9][9] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18325_ (.D(_03903_),
    .Q(\design_top.core0.REG1[9][10] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18326_ (.D(_03904_),
    .Q(\design_top.core0.REG1[9][11] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18327_ (.D(_03905_),
    .Q(\design_top.core0.REG1[9][12] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18328_ (.D(_03906_),
    .Q(\design_top.core0.REG1[9][13] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18329_ (.D(_03907_),
    .Q(\design_top.core0.REG1[9][14] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18330_ (.D(_03908_),
    .Q(\design_top.core0.REG1[9][15] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18331_ (.D(_03909_),
    .Q(\design_top.core0.REG1[9][16] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18332_ (.D(_03910_),
    .Q(\design_top.core0.REG1[9][17] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18333_ (.D(_03911_),
    .Q(\design_top.core0.REG1[9][18] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18334_ (.D(_03912_),
    .Q(\design_top.core0.REG1[9][19] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18335_ (.D(_03913_),
    .Q(\design_top.core0.REG1[9][20] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18336_ (.D(_03914_),
    .Q(\design_top.core0.REG1[9][21] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18337_ (.D(_03915_),
    .Q(\design_top.core0.REG1[9][22] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18338_ (.D(_03916_),
    .Q(\design_top.core0.REG1[9][23] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18339_ (.D(_03917_),
    .Q(\design_top.core0.REG1[9][24] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18340_ (.D(_03918_),
    .Q(\design_top.core0.REG1[9][25] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18341_ (.D(_03919_),
    .Q(\design_top.core0.REG1[9][26] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18342_ (.D(_03920_),
    .Q(\design_top.core0.REG1[9][27] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18343_ (.D(_03921_),
    .Q(\design_top.core0.REG1[9][28] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18344_ (.D(_03922_),
    .Q(\design_top.core0.REG1[9][29] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18345_ (.D(_03923_),
    .Q(\design_top.core0.REG1[9][30] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18346_ (.D(_03924_),
    .Q(\design_top.core0.REG1[9][31] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18347_ (.D(_03925_),
    .Q(\design_top.MEM[6][0] ),
    .CLK(clknet_leaf_250_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18348_ (.D(_03926_),
    .Q(\design_top.MEM[6][1] ),
    .CLK(clknet_leaf_250_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18349_ (.D(_03927_),
    .Q(\design_top.MEM[6][2] ),
    .CLK(clknet_leaf_249_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18350_ (.D(_03928_),
    .Q(\design_top.MEM[6][3] ),
    .CLK(clknet_leaf_246_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18351_ (.D(_03929_),
    .Q(\design_top.MEM[6][4] ),
    .CLK(clknet_leaf_246_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18352_ (.D(_03930_),
    .Q(\design_top.MEM[6][5] ),
    .CLK(clknet_leaf_246_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18353_ (.D(_03931_),
    .Q(\design_top.MEM[6][6] ),
    .CLK(clknet_leaf_246_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18354_ (.D(_03932_),
    .Q(\design_top.MEM[6][7] ),
    .CLK(clknet_leaf_246_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18355_ (.D(_03933_),
    .Q(\design_top.MEM[5][0] ),
    .CLK(clknet_leaf_249_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18356_ (.D(_03934_),
    .Q(\design_top.MEM[5][1] ),
    .CLK(clknet_leaf_250_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18357_ (.D(_03935_),
    .Q(\design_top.MEM[5][2] ),
    .CLK(clknet_leaf_249_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18358_ (.D(_03936_),
    .Q(\design_top.MEM[5][3] ),
    .CLK(clknet_leaf_245_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18359_ (.D(_03937_),
    .Q(\design_top.MEM[5][4] ),
    .CLK(clknet_leaf_247_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18360_ (.D(_03938_),
    .Q(\design_top.MEM[5][5] ),
    .CLK(clknet_leaf_245_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18361_ (.D(_03939_),
    .Q(\design_top.MEM[5][6] ),
    .CLK(clknet_leaf_245_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18362_ (.D(_03940_),
    .Q(\design_top.MEM[5][7] ),
    .CLK(clknet_leaf_245_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18363_ (.D(_03941_),
    .Q(\design_top.core0.REG1[14][0] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18364_ (.D(_03942_),
    .Q(\design_top.core0.REG1[14][1] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18365_ (.D(_03943_),
    .Q(\design_top.core0.REG1[14][2] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18366_ (.D(_03944_),
    .Q(\design_top.core0.REG1[14][3] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18367_ (.D(_03945_),
    .Q(\design_top.core0.REG1[14][4] ),
    .CLK(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18368_ (.D(_03946_),
    .Q(\design_top.core0.REG1[14][5] ),
    .CLK(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18369_ (.D(_03947_),
    .Q(\design_top.core0.REG1[14][6] ),
    .CLK(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18370_ (.D(_03948_),
    .Q(\design_top.core0.REG1[14][7] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18371_ (.D(_03949_),
    .Q(\design_top.core0.REG1[14][8] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18372_ (.D(_03950_),
    .Q(\design_top.core0.REG1[14][9] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18373_ (.D(_03951_),
    .Q(\design_top.core0.REG1[14][10] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18374_ (.D(_03952_),
    .Q(\design_top.core0.REG1[14][11] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18375_ (.D(_03953_),
    .Q(\design_top.core0.REG1[14][12] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18376_ (.D(_03954_),
    .Q(\design_top.core0.REG1[14][13] ),
    .CLK(clknet_leaf_155_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18377_ (.D(_03955_),
    .Q(\design_top.core0.REG1[14][14] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18378_ (.D(_03956_),
    .Q(\design_top.core0.REG1[14][15] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18379_ (.D(_03957_),
    .Q(\design_top.core0.REG1[14][16] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18380_ (.D(_03958_),
    .Q(\design_top.core0.REG1[14][17] ),
    .CLK(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18381_ (.D(_03959_),
    .Q(\design_top.core0.REG1[14][18] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18382_ (.D(_03960_),
    .Q(\design_top.core0.REG1[14][19] ),
    .CLK(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18383_ (.D(_03961_),
    .Q(\design_top.core0.REG1[14][20] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18384_ (.D(_03962_),
    .Q(\design_top.core0.REG1[14][21] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18385_ (.D(_03963_),
    .Q(\design_top.core0.REG1[14][22] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18386_ (.D(_03964_),
    .Q(\design_top.core0.REG1[14][23] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18387_ (.D(_03965_),
    .Q(\design_top.core0.REG1[14][24] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18388_ (.D(_03966_),
    .Q(\design_top.core0.REG1[14][25] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18389_ (.D(_03967_),
    .Q(\design_top.core0.REG1[14][26] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18390_ (.D(_03968_),
    .Q(\design_top.core0.REG1[14][27] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18391_ (.D(_03969_),
    .Q(\design_top.core0.REG1[14][28] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18392_ (.D(_03970_),
    .Q(\design_top.core0.REG1[14][29] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18393_ (.D(_03971_),
    .Q(\design_top.core0.REG1[14][30] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18394_ (.D(_03972_),
    .Q(\design_top.core0.REG1[14][31] ),
    .CLK(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18395_ (.D(_03973_),
    .Q(\design_top.core0.REG1[13][0] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18396_ (.D(_03974_),
    .Q(\design_top.core0.REG1[13][1] ),
    .CLK(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18397_ (.D(_03975_),
    .Q(\design_top.core0.REG1[13][2] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18398_ (.D(_03976_),
    .Q(\design_top.core0.REG1[13][3] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18399_ (.D(_03977_),
    .Q(\design_top.core0.REG1[13][4] ),
    .CLK(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18400_ (.D(_03978_),
    .Q(\design_top.core0.REG1[13][5] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18401_ (.D(_03979_),
    .Q(\design_top.core0.REG1[13][6] ),
    .CLK(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18402_ (.D(_03980_),
    .Q(\design_top.core0.REG1[13][7] ),
    .CLK(clknet_leaf_48_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18403_ (.D(_03981_),
    .Q(\design_top.core0.REG1[13][8] ),
    .CLK(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18404_ (.D(_03982_),
    .Q(\design_top.core0.REG1[13][9] ),
    .CLK(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18405_ (.D(_03983_),
    .Q(\design_top.core0.REG1[13][10] ),
    .CLK(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18406_ (.D(_03984_),
    .Q(\design_top.core0.REG1[13][11] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18407_ (.D(_03985_),
    .Q(\design_top.core0.REG1[13][12] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18408_ (.D(_03986_),
    .Q(\design_top.core0.REG1[13][13] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18409_ (.D(_03987_),
    .Q(\design_top.core0.REG1[13][14] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18410_ (.D(_03988_),
    .Q(\design_top.core0.REG1[13][15] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18411_ (.D(_03989_),
    .Q(\design_top.core0.REG1[13][16] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18412_ (.D(_03990_),
    .Q(\design_top.core0.REG1[13][17] ),
    .CLK(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18413_ (.D(_03991_),
    .Q(\design_top.core0.REG1[13][18] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18414_ (.D(_03992_),
    .Q(\design_top.core0.REG1[13][19] ),
    .CLK(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18415_ (.D(_03993_),
    .Q(\design_top.core0.REG1[13][20] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18416_ (.D(_03994_),
    .Q(\design_top.core0.REG1[13][21] ),
    .CLK(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18417_ (.D(_03995_),
    .Q(\design_top.core0.REG1[13][22] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18418_ (.D(_03996_),
    .Q(\design_top.core0.REG1[13][23] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18419_ (.D(_03997_),
    .Q(\design_top.core0.REG1[13][24] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18420_ (.D(_03998_),
    .Q(\design_top.core0.REG1[13][25] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18421_ (.D(_03999_),
    .Q(\design_top.core0.REG1[13][26] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18422_ (.D(_04000_),
    .Q(\design_top.core0.REG1[13][27] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18423_ (.D(_04001_),
    .Q(\design_top.core0.REG1[13][28] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18424_ (.D(_04002_),
    .Q(\design_top.core0.REG1[13][29] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18425_ (.D(_04003_),
    .Q(\design_top.core0.REG1[13][30] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18426_ (.D(_04004_),
    .Q(\design_top.core0.REG1[13][31] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18427_ (.D(_04005_),
    .Q(\design_top.core0.REG1[12][0] ),
    .CLK(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18428_ (.D(_04006_),
    .Q(\design_top.core0.REG1[12][1] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18429_ (.D(_04007_),
    .Q(\design_top.core0.REG1[12][2] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18430_ (.D(_04008_),
    .Q(\design_top.core0.REG1[12][3] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18431_ (.D(_04009_),
    .Q(\design_top.core0.REG1[12][4] ),
    .CLK(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18432_ (.D(_04010_),
    .Q(\design_top.core0.REG1[12][5] ),
    .CLK(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18433_ (.D(_04011_),
    .Q(\design_top.core0.REG1[12][6] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18434_ (.D(_04012_),
    .Q(\design_top.core0.REG1[12][7] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18435_ (.D(_04013_),
    .Q(\design_top.core0.REG1[12][8] ),
    .CLK(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18436_ (.D(_04014_),
    .Q(\design_top.core0.REG1[12][9] ),
    .CLK(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18437_ (.D(_04015_),
    .Q(\design_top.core0.REG1[12][10] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18438_ (.D(_04016_),
    .Q(\design_top.core0.REG1[12][11] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18439_ (.D(_04017_),
    .Q(\design_top.core0.REG1[12][12] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18440_ (.D(_04018_),
    .Q(\design_top.core0.REG1[12][13] ),
    .CLK(clknet_leaf_155_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18441_ (.D(_04019_),
    .Q(\design_top.core0.REG1[12][14] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18442_ (.D(_04020_),
    .Q(\design_top.core0.REG1[12][15] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18443_ (.D(_04021_),
    .Q(\design_top.core0.REG1[12][16] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18444_ (.D(_04022_),
    .Q(\design_top.core0.REG1[12][17] ),
    .CLK(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18445_ (.D(_04023_),
    .Q(\design_top.core0.REG1[12][18] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18446_ (.D(_04024_),
    .Q(\design_top.core0.REG1[12][19] ),
    .CLK(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18447_ (.D(_04025_),
    .Q(\design_top.core0.REG1[12][20] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18448_ (.D(_04026_),
    .Q(\design_top.core0.REG1[12][21] ),
    .CLK(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18449_ (.D(_04027_),
    .Q(\design_top.core0.REG1[12][22] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18450_ (.D(_04028_),
    .Q(\design_top.core0.REG1[12][23] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18451_ (.D(_04029_),
    .Q(\design_top.core0.REG1[12][24] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18452_ (.D(_04030_),
    .Q(\design_top.core0.REG1[12][25] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18453_ (.D(_04031_),
    .Q(\design_top.core0.REG1[12][26] ),
    .CLK(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18454_ (.D(_04032_),
    .Q(\design_top.core0.REG1[12][27] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18455_ (.D(_04033_),
    .Q(\design_top.core0.REG1[12][28] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18456_ (.D(_04034_),
    .Q(\design_top.core0.REG1[12][29] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18457_ (.D(_04035_),
    .Q(\design_top.core0.REG1[12][30] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18458_ (.D(_04036_),
    .Q(\design_top.core0.REG1[12][31] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18459_ (.D(_04037_),
    .Q(\design_top.core0.REG1[11][0] ),
    .CLK(clknet_leaf_155_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18460_ (.D(_04038_),
    .Q(\design_top.core0.REG1[11][1] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18461_ (.D(_04039_),
    .Q(\design_top.core0.REG1[11][2] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18462_ (.D(_04040_),
    .Q(\design_top.core0.REG1[11][3] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18463_ (.D(_04041_),
    .Q(\design_top.core0.REG1[11][4] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18464_ (.D(_04042_),
    .Q(\design_top.core0.REG1[11][5] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18465_ (.D(_04043_),
    .Q(\design_top.core0.REG1[11][6] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18466_ (.D(_04044_),
    .Q(\design_top.core0.REG1[11][7] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18467_ (.D(_04045_),
    .Q(\design_top.core0.REG1[11][8] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18468_ (.D(_04046_),
    .Q(\design_top.core0.REG1[11][9] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18469_ (.D(_04047_),
    .Q(\design_top.core0.REG1[11][10] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18470_ (.D(_04048_),
    .Q(\design_top.core0.REG1[11][11] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18471_ (.D(_04049_),
    .Q(\design_top.core0.REG1[11][12] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18472_ (.D(_04050_),
    .Q(\design_top.core0.REG1[11][13] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18473_ (.D(_04051_),
    .Q(\design_top.core0.REG1[11][14] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18474_ (.D(_04052_),
    .Q(\design_top.core0.REG1[11][15] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18475_ (.D(_04053_),
    .Q(\design_top.core0.REG1[11][16] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18476_ (.D(_04054_),
    .Q(\design_top.core0.REG1[11][17] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18477_ (.D(_04055_),
    .Q(\design_top.core0.REG1[11][18] ),
    .CLK(clknet_leaf_155_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18478_ (.D(_04056_),
    .Q(\design_top.core0.REG1[11][19] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18479_ (.D(_04057_),
    .Q(\design_top.core0.REG1[11][20] ),
    .CLK(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18480_ (.D(_04058_),
    .Q(\design_top.core0.REG1[11][21] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18481_ (.D(_04059_),
    .Q(\design_top.core0.REG1[11][22] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18482_ (.D(_04060_),
    .Q(\design_top.core0.REG1[11][23] ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18483_ (.D(_04061_),
    .Q(\design_top.core0.REG1[11][24] ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18484_ (.D(_04062_),
    .Q(\design_top.core0.REG1[11][25] ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18485_ (.D(_04063_),
    .Q(\design_top.core0.REG1[11][26] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18486_ (.D(_04064_),
    .Q(\design_top.core0.REG1[11][27] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18487_ (.D(_04065_),
    .Q(\design_top.core0.REG1[11][28] ),
    .CLK(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18488_ (.D(_04066_),
    .Q(\design_top.core0.REG1[11][29] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18489_ (.D(_04067_),
    .Q(\design_top.core0.REG1[11][30] ),
    .CLK(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18490_ (.D(_04068_),
    .Q(\design_top.core0.REG1[11][31] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18491_ (.D(_04069_),
    .Q(\design_top.core0.REG1[10][0] ),
    .CLK(clknet_leaf_155_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18492_ (.D(_04070_),
    .Q(\design_top.core0.REG1[10][1] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18493_ (.D(_04071_),
    .Q(\design_top.core0.REG1[10][2] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18494_ (.D(_04072_),
    .Q(\design_top.core0.REG1[10][3] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18495_ (.D(_04073_),
    .Q(\design_top.core0.REG1[10][4] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18496_ (.D(_04074_),
    .Q(\design_top.core0.REG1[10][5] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18497_ (.D(_04075_),
    .Q(\design_top.core0.REG1[10][6] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18498_ (.D(_04076_),
    .Q(\design_top.core0.REG1[10][7] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18499_ (.D(_04077_),
    .Q(\design_top.core0.REG1[10][8] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18500_ (.D(_04078_),
    .Q(\design_top.core0.REG1[10][9] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18501_ (.D(_04079_),
    .Q(\design_top.core0.REG1[10][10] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18502_ (.D(_04080_),
    .Q(\design_top.core0.REG1[10][11] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18503_ (.D(_04081_),
    .Q(\design_top.core0.REG1[10][12] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18504_ (.D(_04082_),
    .Q(\design_top.core0.REG1[10][13] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18505_ (.D(_04083_),
    .Q(\design_top.core0.REG1[10][14] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18506_ (.D(_04084_),
    .Q(\design_top.core0.REG1[10][15] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18507_ (.D(_04085_),
    .Q(\design_top.core0.REG1[10][16] ),
    .CLK(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18508_ (.D(_04086_),
    .Q(\design_top.core0.REG1[10][17] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18509_ (.D(_04087_),
    .Q(\design_top.core0.REG1[10][18] ),
    .CLK(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18510_ (.D(_04088_),
    .Q(\design_top.core0.REG1[10][19] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18511_ (.D(_04089_),
    .Q(\design_top.core0.REG1[10][20] ),
    .CLK(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18512_ (.D(_04090_),
    .Q(\design_top.core0.REG1[10][21] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18513_ (.D(_04091_),
    .Q(\design_top.core0.REG1[10][22] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18514_ (.D(_04092_),
    .Q(\design_top.core0.REG1[10][23] ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18515_ (.D(_04093_),
    .Q(\design_top.core0.REG1[10][24] ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18516_ (.D(_04094_),
    .Q(\design_top.core0.REG1[10][25] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18517_ (.D(_04095_),
    .Q(\design_top.core0.REG1[10][26] ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18518_ (.D(_04096_),
    .Q(\design_top.core0.REG1[10][27] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18519_ (.D(_04097_),
    .Q(\design_top.core0.REG1[10][28] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18520_ (.D(_04098_),
    .Q(\design_top.core0.REG1[10][29] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18521_ (.D(_04099_),
    .Q(\design_top.core0.REG1[10][30] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18522_ (.D(_04100_),
    .Q(\design_top.core0.REG1[10][31] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18523_ (.D(_04101_),
    .Q(\design_top.core0.REG1[0][0] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18524_ (.D(_04102_),
    .Q(\design_top.core0.REG1[0][1] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18525_ (.D(_04103_),
    .Q(\design_top.core0.REG1[0][2] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18526_ (.D(_04104_),
    .Q(\design_top.core0.REG1[0][3] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18527_ (.D(_04105_),
    .Q(\design_top.core0.REG1[0][4] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18528_ (.D(_04106_),
    .Q(\design_top.core0.REG1[0][5] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18529_ (.D(_04107_),
    .Q(\design_top.core0.REG1[0][6] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18530_ (.D(_04108_),
    .Q(\design_top.core0.REG1[0][7] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18531_ (.D(_04109_),
    .Q(\design_top.core0.REG1[0][8] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18532_ (.D(_04110_),
    .Q(\design_top.core0.REG1[0][9] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18533_ (.D(_04111_),
    .Q(\design_top.core0.REG1[0][10] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18534_ (.D(_04112_),
    .Q(\design_top.core0.REG1[0][11] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18535_ (.D(_04113_),
    .Q(\design_top.core0.REG1[0][12] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18536_ (.D(_04114_),
    .Q(\design_top.core0.REG1[0][13] ),
    .CLK(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18537_ (.D(_04115_),
    .Q(\design_top.core0.REG1[0][14] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18538_ (.D(_04116_),
    .Q(\design_top.core0.REG1[0][15] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18539_ (.D(_04117_),
    .Q(\design_top.core0.REG1[0][16] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18540_ (.D(_04118_),
    .Q(\design_top.core0.REG1[0][17] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18541_ (.D(_04119_),
    .Q(\design_top.core0.REG1[0][18] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18542_ (.D(_04120_),
    .Q(\design_top.core0.REG1[0][19] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18543_ (.D(_04121_),
    .Q(\design_top.core0.REG1[0][20] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18544_ (.D(_04122_),
    .Q(\design_top.core0.REG1[0][21] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18545_ (.D(_04123_),
    .Q(\design_top.core0.REG1[0][22] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18546_ (.D(_04124_),
    .Q(\design_top.core0.REG1[0][23] ),
    .CLK(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18547_ (.D(_04125_),
    .Q(\design_top.core0.REG1[0][24] ),
    .CLK(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18548_ (.D(_04126_),
    .Q(\design_top.core0.REG1[0][25] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18549_ (.D(_04127_),
    .Q(\design_top.core0.REG1[0][26] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18550_ (.D(_04128_),
    .Q(\design_top.core0.REG1[0][27] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18551_ (.D(_04129_),
    .Q(\design_top.core0.REG1[0][28] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18552_ (.D(_04130_),
    .Q(\design_top.core0.REG1[0][29] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18553_ (.D(_04131_),
    .Q(\design_top.core0.REG1[0][30] ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18554_ (.D(_04132_),
    .Q(\design_top.core0.REG1[0][31] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18555_ (.D(_04133_),
    .Q(\design_top.core0.REG1[8][0] ),
    .CLK(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18556_ (.D(_04134_),
    .Q(\design_top.core0.REG1[8][1] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18557_ (.D(_04135_),
    .Q(\design_top.core0.REG1[8][2] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18558_ (.D(_04136_),
    .Q(\design_top.core0.REG1[8][3] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18559_ (.D(_04137_),
    .Q(\design_top.core0.REG1[8][4] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18560_ (.D(_04138_),
    .Q(\design_top.core0.REG1[8][5] ),
    .CLK(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18561_ (.D(_04139_),
    .Q(\design_top.core0.REG1[8][6] ),
    .CLK(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18562_ (.D(_04140_),
    .Q(\design_top.core0.REG1[8][7] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18563_ (.D(_04141_),
    .Q(\design_top.core0.REG1[8][8] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18564_ (.D(_04142_),
    .Q(\design_top.core0.REG1[8][9] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18565_ (.D(_04143_),
    .Q(\design_top.core0.REG1[8][10] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18566_ (.D(_04144_),
    .Q(\design_top.core0.REG1[8][11] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18567_ (.D(_04145_),
    .Q(\design_top.core0.REG1[8][12] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18568_ (.D(_04146_),
    .Q(\design_top.core0.REG1[8][13] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18569_ (.D(_04147_),
    .Q(\design_top.core0.REG1[8][14] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18570_ (.D(_04148_),
    .Q(\design_top.core0.REG1[8][15] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18571_ (.D(_04149_),
    .Q(\design_top.core0.REG1[8][16] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18572_ (.D(_04150_),
    .Q(\design_top.core0.REG1[8][17] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18573_ (.D(_04151_),
    .Q(\design_top.core0.REG1[8][18] ),
    .CLK(clknet_leaf_155_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18574_ (.D(_04152_),
    .Q(\design_top.core0.REG1[8][19] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18575_ (.D(_04153_),
    .Q(\design_top.core0.REG1[8][20] ),
    .CLK(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18576_ (.D(_04154_),
    .Q(\design_top.core0.REG1[8][21] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18577_ (.D(_04155_),
    .Q(\design_top.core0.REG1[8][22] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18578_ (.D(_04156_),
    .Q(\design_top.core0.REG1[8][23] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18579_ (.D(_04157_),
    .Q(\design_top.core0.REG1[8][24] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18580_ (.D(_04158_),
    .Q(\design_top.core0.REG1[8][25] ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18581_ (.D(_04159_),
    .Q(\design_top.core0.REG1[8][26] ),
    .CLK(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18582_ (.D(_04160_),
    .Q(\design_top.core0.REG1[8][27] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18583_ (.D(_04161_),
    .Q(\design_top.core0.REG1[8][28] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18584_ (.D(_04162_),
    .Q(\design_top.core0.REG1[8][29] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18585_ (.D(_04163_),
    .Q(\design_top.core0.REG1[8][30] ),
    .CLK(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18586_ (.D(_04164_),
    .Q(\design_top.core0.REG1[8][31] ),
    .CLK(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18587_ (.D(_04165_),
    .Q(\design_top.MEM[4][0] ),
    .CLK(clknet_leaf_250_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18588_ (.D(_04166_),
    .Q(\design_top.MEM[4][1] ),
    .CLK(clknet_leaf_250_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18589_ (.D(_04167_),
    .Q(\design_top.MEM[4][2] ),
    .CLK(clknet_leaf_249_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18590_ (.D(_04168_),
    .Q(\design_top.MEM[4][3] ),
    .CLK(clknet_leaf_245_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18591_ (.D(_04169_),
    .Q(\design_top.MEM[4][4] ),
    .CLK(clknet_leaf_246_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18592_ (.D(_04170_),
    .Q(\design_top.MEM[4][5] ),
    .CLK(clknet_leaf_245_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18593_ (.D(_04171_),
    .Q(\design_top.MEM[4][6] ),
    .CLK(clknet_leaf_244_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18594_ (.D(_04172_),
    .Q(\design_top.MEM[4][7] ),
    .CLK(clknet_leaf_244_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18595_ (.D(_04173_),
    .Q(\design_top.core0.REG1[7][0] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18596_ (.D(_04174_),
    .Q(\design_top.core0.REG1[7][1] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18597_ (.D(_04175_),
    .Q(\design_top.core0.REG1[7][2] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18598_ (.D(_04176_),
    .Q(\design_top.core0.REG1[7][3] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18599_ (.D(_04177_),
    .Q(\design_top.core0.REG1[7][4] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18600_ (.D(_04178_),
    .Q(\design_top.core0.REG1[7][5] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18601_ (.D(_04179_),
    .Q(\design_top.core0.REG1[7][6] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18602_ (.D(_04180_),
    .Q(\design_top.core0.REG1[7][7] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18603_ (.D(_04181_),
    .Q(\design_top.core0.REG1[7][8] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18604_ (.D(_04182_),
    .Q(\design_top.core0.REG1[7][9] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18605_ (.D(_04183_),
    .Q(\design_top.core0.REG1[7][10] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18606_ (.D(_04184_),
    .Q(\design_top.core0.REG1[7][11] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18607_ (.D(_04185_),
    .Q(\design_top.core0.REG1[7][12] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18608_ (.D(_04186_),
    .Q(\design_top.core0.REG1[7][13] ),
    .CLK(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18609_ (.D(_04187_),
    .Q(\design_top.core0.REG1[7][14] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18610_ (.D(_04188_),
    .Q(\design_top.core0.REG1[7][15] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18611_ (.D(_04189_),
    .Q(\design_top.core0.REG1[7][16] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18612_ (.D(_04190_),
    .Q(\design_top.core0.REG1[7][17] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18613_ (.D(_04191_),
    .Q(\design_top.core0.REG1[7][18] ),
    .CLK(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18614_ (.D(_04192_),
    .Q(\design_top.core0.REG1[7][19] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18615_ (.D(_04193_),
    .Q(\design_top.core0.REG1[7][20] ),
    .CLK(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18616_ (.D(_04194_),
    .Q(\design_top.core0.REG1[7][21] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18617_ (.D(_04195_),
    .Q(\design_top.core0.REG1[7][22] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18618_ (.D(_04196_),
    .Q(\design_top.core0.REG1[7][23] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18619_ (.D(_04197_),
    .Q(\design_top.core0.REG1[7][24] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18620_ (.D(_04198_),
    .Q(\design_top.core0.REG1[7][25] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18621_ (.D(_04199_),
    .Q(\design_top.core0.REG1[7][26] ),
    .CLK(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18622_ (.D(_04200_),
    .Q(\design_top.core0.REG1[7][27] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18623_ (.D(_04201_),
    .Q(\design_top.core0.REG1[7][28] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18624_ (.D(_04202_),
    .Q(\design_top.core0.REG1[7][29] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18625_ (.D(_04203_),
    .Q(\design_top.core0.REG1[7][30] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18626_ (.D(_04204_),
    .Q(\design_top.core0.REG1[7][31] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18627_ (.D(_04205_),
    .Q(\design_top.core0.REG1[6][0] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18628_ (.D(_04206_),
    .Q(\design_top.core0.REG1[6][1] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18629_ (.D(_04207_),
    .Q(\design_top.core0.REG1[6][2] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18630_ (.D(_04208_),
    .Q(\design_top.core0.REG1[6][3] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18631_ (.D(_04209_),
    .Q(\design_top.core0.REG1[6][4] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18632_ (.D(_04210_),
    .Q(\design_top.core0.REG1[6][5] ),
    .CLK(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18633_ (.D(_04211_),
    .Q(\design_top.core0.REG1[6][6] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18634_ (.D(_04212_),
    .Q(\design_top.core0.REG1[6][7] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18635_ (.D(_04213_),
    .Q(\design_top.core0.REG1[6][8] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18636_ (.D(_04214_),
    .Q(\design_top.core0.REG1[6][9] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18637_ (.D(_04215_),
    .Q(\design_top.core0.REG1[6][10] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18638_ (.D(_04216_),
    .Q(\design_top.core0.REG1[6][11] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18639_ (.D(_04217_),
    .Q(\design_top.core0.REG1[6][12] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18640_ (.D(_04218_),
    .Q(\design_top.core0.REG1[6][13] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18641_ (.D(_04219_),
    .Q(\design_top.core0.REG1[6][14] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18642_ (.D(_04220_),
    .Q(\design_top.core0.REG1[6][15] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18643_ (.D(_04221_),
    .Q(\design_top.core0.REG1[6][16] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18644_ (.D(_04222_),
    .Q(\design_top.core0.REG1[6][17] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18645_ (.D(_04223_),
    .Q(\design_top.core0.REG1[6][18] ),
    .CLK(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18646_ (.D(_04224_),
    .Q(\design_top.core0.REG1[6][19] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18647_ (.D(_04225_),
    .Q(\design_top.core0.REG1[6][20] ),
    .CLK(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18648_ (.D(_04226_),
    .Q(\design_top.core0.REG1[6][21] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18649_ (.D(_04227_),
    .Q(\design_top.core0.REG1[6][22] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18650_ (.D(_04228_),
    .Q(\design_top.core0.REG1[6][23] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18651_ (.D(_04229_),
    .Q(\design_top.core0.REG1[6][24] ),
    .CLK(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18652_ (.D(_04230_),
    .Q(\design_top.core0.REG1[6][25] ),
    .CLK(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18653_ (.D(_04231_),
    .Q(\design_top.core0.REG1[6][26] ),
    .CLK(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18654_ (.D(_04232_),
    .Q(\design_top.core0.REG1[6][27] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18655_ (.D(_04233_),
    .Q(\design_top.core0.REG1[6][28] ),
    .CLK(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18656_ (.D(_04234_),
    .Q(\design_top.core0.REG1[6][29] ),
    .CLK(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18657_ (.D(_04235_),
    .Q(\design_top.core0.REG1[6][30] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18658_ (.D(_04236_),
    .Q(\design_top.core0.REG1[6][31] ),
    .CLK(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18659_ (.D(_04237_),
    .Q(\design_top.core0.REG1[5][0] ),
    .CLK(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18660_ (.D(_04238_),
    .Q(\design_top.core0.REG1[5][1] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18661_ (.D(_04239_),
    .Q(\design_top.core0.REG1[5][2] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18662_ (.D(_04240_),
    .Q(\design_top.core0.REG1[5][3] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18663_ (.D(_04241_),
    .Q(\design_top.core0.REG1[5][4] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18664_ (.D(_04242_),
    .Q(\design_top.core0.REG1[5][5] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18665_ (.D(_04243_),
    .Q(\design_top.core0.REG1[5][6] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18666_ (.D(_04244_),
    .Q(\design_top.core0.REG1[5][7] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18667_ (.D(_04245_),
    .Q(\design_top.core0.REG1[5][8] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18668_ (.D(_04246_),
    .Q(\design_top.core0.REG1[5][9] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18669_ (.D(_04247_),
    .Q(\design_top.core0.REG1[5][10] ),
    .CLK(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18670_ (.D(_04248_),
    .Q(\design_top.core0.REG1[5][11] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18671_ (.D(_04249_),
    .Q(\design_top.core0.REG1[5][12] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18672_ (.D(_04250_),
    .Q(\design_top.core0.REG1[5][13] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18673_ (.D(_04251_),
    .Q(\design_top.core0.REG1[5][14] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18674_ (.D(_04252_),
    .Q(\design_top.core0.REG1[5][15] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18675_ (.D(_04253_),
    .Q(\design_top.core0.REG1[5][16] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18676_ (.D(_04254_),
    .Q(\design_top.core0.REG1[5][17] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18677_ (.D(_04255_),
    .Q(\design_top.core0.REG1[5][18] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18678_ (.D(_04256_),
    .Q(\design_top.core0.REG1[5][19] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18679_ (.D(_04257_),
    .Q(\design_top.core0.REG1[5][20] ),
    .CLK(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18680_ (.D(_04258_),
    .Q(\design_top.core0.REG1[5][21] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18681_ (.D(_04259_),
    .Q(\design_top.core0.REG1[5][22] ),
    .CLK(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18682_ (.D(_04260_),
    .Q(\design_top.core0.REG1[5][23] ),
    .CLK(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18683_ (.D(_04261_),
    .Q(\design_top.core0.REG1[5][24] ),
    .CLK(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18684_ (.D(_04262_),
    .Q(\design_top.core0.REG1[5][25] ),
    .CLK(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18685_ (.D(_04263_),
    .Q(\design_top.core0.REG1[5][26] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18686_ (.D(_04264_),
    .Q(\design_top.core0.REG1[5][27] ),
    .CLK(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18687_ (.D(_04265_),
    .Q(\design_top.core0.REG1[5][28] ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18688_ (.D(_04266_),
    .Q(\design_top.core0.REG1[5][29] ),
    .CLK(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18689_ (.D(_04267_),
    .Q(\design_top.core0.REG1[5][30] ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18690_ (.D(_04268_),
    .Q(\design_top.core0.REG1[5][31] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18691_ (.D(_04269_),
    .Q(\design_top.core0.REG1[4][0] ),
    .CLK(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18692_ (.D(_04270_),
    .Q(\design_top.core0.REG1[4][1] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18693_ (.D(_04271_),
    .Q(\design_top.core0.REG1[4][2] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18694_ (.D(_04272_),
    .Q(\design_top.core0.REG1[4][3] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18695_ (.D(_04273_),
    .Q(\design_top.core0.REG1[4][4] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18696_ (.D(_04274_),
    .Q(\design_top.core0.REG1[4][5] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18697_ (.D(_04275_),
    .Q(\design_top.core0.REG1[4][6] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18698_ (.D(_04276_),
    .Q(\design_top.core0.REG1[4][7] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18699_ (.D(_04277_),
    .Q(\design_top.core0.REG1[4][8] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18700_ (.D(_04278_),
    .Q(\design_top.core0.REG1[4][9] ),
    .CLK(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18701_ (.D(_04279_),
    .Q(\design_top.core0.REG1[4][10] ),
    .CLK(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18702_ (.D(_04280_),
    .Q(\design_top.core0.REG1[4][11] ),
    .CLK(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18703_ (.D(_04281_),
    .Q(\design_top.core0.REG1[4][12] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18704_ (.D(_04282_),
    .Q(\design_top.core0.REG1[4][13] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18705_ (.D(_04283_),
    .Q(\design_top.core0.REG1[4][14] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18706_ (.D(_04284_),
    .Q(\design_top.core0.REG1[4][15] ),
    .CLK(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18707_ (.D(_04285_),
    .Q(\design_top.core0.REG1[4][16] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18708_ (.D(_04286_),
    .Q(\design_top.core0.REG1[4][17] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18709_ (.D(_04287_),
    .Q(\design_top.core0.REG1[4][18] ),
    .CLK(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18710_ (.D(_04288_),
    .Q(\design_top.core0.REG1[4][19] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18711_ (.D(_04289_),
    .Q(\design_top.core0.REG1[4][20] ),
    .CLK(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18712_ (.D(_04290_),
    .Q(\design_top.core0.REG1[4][21] ),
    .CLK(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18713_ (.D(_04291_),
    .Q(\design_top.core0.REG1[4][22] ),
    .CLK(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18714_ (.D(_04292_),
    .Q(\design_top.core0.REG1[4][23] ),
    .CLK(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18715_ (.D(_04293_),
    .Q(\design_top.core0.REG1[4][24] ),
    .CLK(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18716_ (.D(_04294_),
    .Q(\design_top.core0.REG1[4][25] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18717_ (.D(_04295_),
    .Q(\design_top.core0.REG1[4][26] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18718_ (.D(_04296_),
    .Q(\design_top.core0.REG1[4][27] ),
    .CLK(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18719_ (.D(_04297_),
    .Q(\design_top.core0.REG1[4][28] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18720_ (.D(_04298_),
    .Q(\design_top.core0.REG1[4][29] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18721_ (.D(_04299_),
    .Q(\design_top.core0.REG1[4][30] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18722_ (.D(_04300_),
    .Q(\design_top.core0.REG1[4][31] ),
    .CLK(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18723_ (.D(_04301_),
    .Q(\design_top.core0.REG1[3][0] ),
    .CLK(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18724_ (.D(_04302_),
    .Q(\design_top.core0.REG1[3][1] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18725_ (.D(_04303_),
    .Q(\design_top.core0.REG1[3][2] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18726_ (.D(_04304_),
    .Q(\design_top.core0.REG1[3][3] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18727_ (.D(_04305_),
    .Q(\design_top.core0.REG1[3][4] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18728_ (.D(_04306_),
    .Q(\design_top.core0.REG1[3][5] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18729_ (.D(_04307_),
    .Q(\design_top.core0.REG1[3][6] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18730_ (.D(_04308_),
    .Q(\design_top.core0.REG1[3][7] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18731_ (.D(_04309_),
    .Q(\design_top.core0.REG1[3][8] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18732_ (.D(_04310_),
    .Q(\design_top.core0.REG1[3][9] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18733_ (.D(_04311_),
    .Q(\design_top.core0.REG1[3][10] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18734_ (.D(_04312_),
    .Q(\design_top.core0.REG1[3][11] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18735_ (.D(_04313_),
    .Q(\design_top.core0.REG1[3][12] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18736_ (.D(_04314_),
    .Q(\design_top.core0.REG1[3][13] ),
    .CLK(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18737_ (.D(_04315_),
    .Q(\design_top.core0.REG1[3][14] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18738_ (.D(_04316_),
    .Q(\design_top.core0.REG1[3][15] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18739_ (.D(_04317_),
    .Q(\design_top.core0.REG1[3][16] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18740_ (.D(_04318_),
    .Q(\design_top.core0.REG1[3][17] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18741_ (.D(_04319_),
    .Q(\design_top.core0.REG1[3][18] ),
    .CLK(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18742_ (.D(_04320_),
    .Q(\design_top.core0.REG1[3][19] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18743_ (.D(_04321_),
    .Q(\design_top.core0.REG1[3][20] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18744_ (.D(_04322_),
    .Q(\design_top.core0.REG1[3][21] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18745_ (.D(_04323_),
    .Q(\design_top.core0.REG1[3][22] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18746_ (.D(_04324_),
    .Q(\design_top.core0.REG1[3][23] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18747_ (.D(_04325_),
    .Q(\design_top.core0.REG1[3][24] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18748_ (.D(_04326_),
    .Q(\design_top.core0.REG1[3][25] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18749_ (.D(_04327_),
    .Q(\design_top.core0.REG1[3][26] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18750_ (.D(_04328_),
    .Q(\design_top.core0.REG1[3][27] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18751_ (.D(_04329_),
    .Q(\design_top.core0.REG1[3][28] ),
    .CLK(clknet_leaf_172_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18752_ (.D(_04330_),
    .Q(\design_top.core0.REG1[3][29] ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18753_ (.D(_04331_),
    .Q(\design_top.core0.REG1[3][30] ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18754_ (.D(_04332_),
    .Q(\design_top.core0.REG1[3][31] ),
    .CLK(clknet_leaf_172_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18755_ (.D(_04333_),
    .Q(\design_top.core0.REG1[2][0] ),
    .CLK(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18756_ (.D(_04334_),
    .Q(\design_top.core0.REG1[2][1] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18757_ (.D(_04335_),
    .Q(\design_top.core0.REG1[2][2] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18758_ (.D(_04336_),
    .Q(\design_top.core0.REG1[2][3] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18759_ (.D(_04337_),
    .Q(\design_top.core0.REG1[2][4] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18760_ (.D(_04338_),
    .Q(\design_top.core0.REG1[2][5] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18761_ (.D(_04339_),
    .Q(\design_top.core0.REG1[2][6] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18762_ (.D(_04340_),
    .Q(\design_top.core0.REG1[2][7] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18763_ (.D(_04341_),
    .Q(\design_top.core0.REG1[2][8] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18764_ (.D(_04342_),
    .Q(\design_top.core0.REG1[2][9] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18765_ (.D(_04343_),
    .Q(\design_top.core0.REG1[2][10] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18766_ (.D(_04344_),
    .Q(\design_top.core0.REG1[2][11] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18767_ (.D(_04345_),
    .Q(\design_top.core0.REG1[2][12] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18768_ (.D(_04346_),
    .Q(\design_top.core0.REG1[2][13] ),
    .CLK(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18769_ (.D(_04347_),
    .Q(\design_top.core0.REG1[2][14] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18770_ (.D(_04348_),
    .Q(\design_top.core0.REG1[2][15] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18771_ (.D(_04349_),
    .Q(\design_top.core0.REG1[2][16] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18772_ (.D(_04350_),
    .Q(\design_top.core0.REG1[2][17] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18773_ (.D(_04351_),
    .Q(\design_top.core0.REG1[2][18] ),
    .CLK(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18774_ (.D(_04352_),
    .Q(\design_top.core0.REG1[2][19] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18775_ (.D(_04353_),
    .Q(\design_top.core0.REG1[2][20] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18776_ (.D(_04354_),
    .Q(\design_top.core0.REG1[2][21] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18777_ (.D(_04355_),
    .Q(\design_top.core0.REG1[2][22] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18778_ (.D(_04356_),
    .Q(\design_top.core0.REG1[2][23] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18779_ (.D(_04357_),
    .Q(\design_top.core0.REG1[2][24] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18780_ (.D(_04358_),
    .Q(\design_top.core0.REG1[2][25] ),
    .CLK(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18781_ (.D(_04359_),
    .Q(\design_top.core0.REG1[2][26] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18782_ (.D(_04360_),
    .Q(\design_top.core0.REG1[2][27] ),
    .CLK(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18783_ (.D(_04361_),
    .Q(\design_top.core0.REG1[2][28] ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18784_ (.D(_04362_),
    .Q(\design_top.core0.REG1[2][29] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18785_ (.D(_04363_),
    .Q(\design_top.core0.REG1[2][30] ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18786_ (.D(_04364_),
    .Q(\design_top.core0.REG1[2][31] ),
    .CLK(clknet_leaf_172_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18787_ (.D(_04365_),
    .Q(\design_top.core0.REG1[1][0] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18788_ (.D(_04366_),
    .Q(\design_top.core0.REG1[1][1] ),
    .CLK(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18789_ (.D(_04367_),
    .Q(\design_top.core0.REG1[1][2] ),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18790_ (.D(_04368_),
    .Q(\design_top.core0.REG1[1][3] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18791_ (.D(_04369_),
    .Q(\design_top.core0.REG1[1][4] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18792_ (.D(_04370_),
    .Q(\design_top.core0.REG1[1][5] ),
    .CLK(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18793_ (.D(_04371_),
    .Q(\design_top.core0.REG1[1][6] ),
    .CLK(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18794_ (.D(_04372_),
    .Q(\design_top.core0.REG1[1][7] ),
    .CLK(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18795_ (.D(_04373_),
    .Q(\design_top.core0.REG1[1][8] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18796_ (.D(_04374_),
    .Q(\design_top.core0.REG1[1][9] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18797_ (.D(_04375_),
    .Q(\design_top.core0.REG1[1][10] ),
    .CLK(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18798_ (.D(_04376_),
    .Q(\design_top.core0.REG1[1][11] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18799_ (.D(_04377_),
    .Q(\design_top.core0.REG1[1][12] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18800_ (.D(_04378_),
    .Q(\design_top.core0.REG1[1][13] ),
    .CLK(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18801_ (.D(_04379_),
    .Q(\design_top.core0.REG1[1][14] ),
    .CLK(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18802_ (.D(_04380_),
    .Q(\design_top.core0.REG1[1][15] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18803_ (.D(_04381_),
    .Q(\design_top.core0.REG1[1][16] ),
    .CLK(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18804_ (.D(_04382_),
    .Q(\design_top.core0.REG1[1][17] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18805_ (.D(_04383_),
    .Q(\design_top.core0.REG1[1][18] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18806_ (.D(_04384_),
    .Q(\design_top.core0.REG1[1][19] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18807_ (.D(_04385_),
    .Q(\design_top.core0.REG1[1][20] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18808_ (.D(_04386_),
    .Q(\design_top.core0.REG1[1][21] ),
    .CLK(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18809_ (.D(_04387_),
    .Q(\design_top.core0.REG1[1][22] ),
    .CLK(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18810_ (.D(_04388_),
    .Q(\design_top.core0.REG1[1][23] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18811_ (.D(_04389_),
    .Q(\design_top.core0.REG1[1][24] ),
    .CLK(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18812_ (.D(_04390_),
    .Q(\design_top.core0.REG1[1][25] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18813_ (.D(_04391_),
    .Q(\design_top.core0.REG1[1][26] ),
    .CLK(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18814_ (.D(_04392_),
    .Q(\design_top.core0.REG1[1][27] ),
    .CLK(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18815_ (.D(_04393_),
    .Q(\design_top.core0.REG1[1][28] ),
    .CLK(clknet_leaf_172_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18816_ (.D(_04394_),
    .Q(\design_top.core0.REG1[1][29] ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18817_ (.D(_04395_),
    .Q(\design_top.core0.REG1[1][30] ),
    .CLK(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18818_ (.D(_04396_),
    .Q(\design_top.core0.REG1[1][31] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18819_ (.D(_04397_),
    .Q(\design_top.core0.REG1[15][0] ),
    .CLK(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18820_ (.D(_04398_),
    .Q(\design_top.core0.REG1[15][1] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18821_ (.D(_04399_),
    .Q(\design_top.core0.REG1[15][2] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18822_ (.D(_04400_),
    .Q(\design_top.core0.REG1[15][3] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18823_ (.D(_04401_),
    .Q(\design_top.core0.REG1[15][4] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18824_ (.D(_04402_),
    .Q(\design_top.core0.REG1[15][5] ),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18825_ (.D(_04403_),
    .Q(\design_top.core0.REG1[15][6] ),
    .CLK(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18826_ (.D(_04404_),
    .Q(\design_top.core0.REG1[15][7] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18827_ (.D(_04405_),
    .Q(\design_top.core0.REG1[15][8] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18828_ (.D(_04406_),
    .Q(\design_top.core0.REG1[15][9] ),
    .CLK(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18829_ (.D(_04407_),
    .Q(\design_top.core0.REG1[15][10] ),
    .CLK(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18830_ (.D(_04408_),
    .Q(\design_top.core0.REG1[15][11] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18831_ (.D(_04409_),
    .Q(\design_top.core0.REG1[15][12] ),
    .CLK(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18832_ (.D(_04410_),
    .Q(\design_top.core0.REG1[15][13] ),
    .CLK(clknet_leaf_155_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18833_ (.D(_04411_),
    .Q(\design_top.core0.REG1[15][14] ),
    .CLK(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18834_ (.D(_04412_),
    .Q(\design_top.core0.REG1[15][15] ),
    .CLK(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18835_ (.D(_04413_),
    .Q(\design_top.core0.REG1[15][16] ),
    .CLK(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18836_ (.D(_04414_),
    .Q(\design_top.core0.REG1[15][17] ),
    .CLK(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18837_ (.D(_04415_),
    .Q(\design_top.core0.REG1[15][18] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18838_ (.D(_04416_),
    .Q(\design_top.core0.REG1[15][19] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18839_ (.D(_04417_),
    .Q(\design_top.core0.REG1[15][20] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18840_ (.D(_04418_),
    .Q(\design_top.core0.REG1[15][21] ),
    .CLK(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18841_ (.D(_04419_),
    .Q(\design_top.core0.REG1[15][22] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18842_ (.D(_04420_),
    .Q(\design_top.core0.REG1[15][23] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18843_ (.D(_04421_),
    .Q(\design_top.core0.REG1[15][24] ),
    .CLK(clknet_leaf_155_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18844_ (.D(_04422_),
    .Q(\design_top.core0.REG1[15][25] ),
    .CLK(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18845_ (.D(_04423_),
    .Q(\design_top.core0.REG1[15][26] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18846_ (.D(_04424_),
    .Q(\design_top.core0.REG1[15][27] ),
    .CLK(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18847_ (.D(_04425_),
    .Q(\design_top.core0.REG1[15][28] ),
    .CLK(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18848_ (.D(_04426_),
    .Q(\design_top.core0.REG1[15][29] ),
    .CLK(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18849_ (.D(_04427_),
    .Q(\design_top.core0.REG1[15][30] ),
    .CLK(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18850_ (.D(_04428_),
    .Q(\design_top.core0.REG1[15][31] ),
    .CLK(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18851_ (.D(_04429_),
    .Q(\design_top.MEM[3][0] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18852_ (.D(_04430_),
    .Q(\design_top.MEM[3][1] ),
    .CLK(clknet_leaf_251_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18853_ (.D(_04431_),
    .Q(\design_top.MEM[3][2] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18854_ (.D(_04432_),
    .Q(\design_top.MEM[3][3] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18855_ (.D(_04433_),
    .Q(\design_top.MEM[3][4] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18856_ (.D(_04434_),
    .Q(\design_top.MEM[3][5] ),
    .CLK(clknet_leaf_247_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18857_ (.D(_04435_),
    .Q(\design_top.MEM[3][6] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18858_ (.D(_04436_),
    .Q(\design_top.MEM[3][7] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18859_ (.D(_04437_),
    .Q(\design_top.MEM[31][0] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18860_ (.D(_04438_),
    .Q(\design_top.MEM[31][1] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18861_ (.D(_04439_),
    .Q(\design_top.MEM[31][2] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18862_ (.D(_04440_),
    .Q(\design_top.MEM[31][3] ),
    .CLK(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18863_ (.D(_04441_),
    .Q(\design_top.MEM[31][4] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18864_ (.D(_04442_),
    .Q(\design_top.MEM[31][5] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18865_ (.D(_04443_),
    .Q(\design_top.MEM[31][6] ),
    .CLK(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18866_ (.D(_04444_),
    .Q(\design_top.MEM[31][7] ),
    .CLK(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18867_ (.D(_04445_),
    .Q(\design_top.MEM[30][0] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18868_ (.D(_04446_),
    .Q(\design_top.MEM[30][1] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18869_ (.D(_04447_),
    .Q(\design_top.MEM[30][2] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18870_ (.D(_04448_),
    .Q(\design_top.MEM[30][3] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18871_ (.D(_04449_),
    .Q(\design_top.MEM[30][4] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18872_ (.D(_04450_),
    .Q(\design_top.MEM[30][5] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18873_ (.D(_04451_),
    .Q(\design_top.MEM[30][6] ),
    .CLK(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18874_ (.D(_04452_),
    .Q(\design_top.MEM[30][7] ),
    .CLK(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18875_ (.D(_04453_),
    .Q(io_out[14]),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18876_ (.D(_04454_),
    .Q(\design_top.MEM[11][0] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18877_ (.D(_04455_),
    .Q(\design_top.MEM[11][1] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18878_ (.D(_04456_),
    .Q(\design_top.MEM[11][2] ),
    .CLK(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18879_ (.D(_04457_),
    .Q(\design_top.MEM[11][3] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18880_ (.D(_04458_),
    .Q(\design_top.MEM[11][4] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18881_ (.D(_04459_),
    .Q(\design_top.MEM[11][5] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18882_ (.D(_04460_),
    .Q(\design_top.MEM[11][6] ),
    .CLK(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18883_ (.D(_04461_),
    .Q(\design_top.MEM[11][7] ),
    .CLK(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18884_ (.D(_04462_),
    .Q(\design_top.TIMER[0] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18885_ (.D(_04463_),
    .Q(\design_top.TIMER[1] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18886_ (.D(_04464_),
    .Q(\design_top.TIMER[2] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18887_ (.D(_04465_),
    .Q(\design_top.TIMER[3] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18888_ (.D(_04466_),
    .Q(\design_top.TIMER[4] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18889_ (.D(_04467_),
    .Q(\design_top.TIMER[5] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18890_ (.D(_04468_),
    .Q(\design_top.TIMER[6] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18891_ (.D(_04469_),
    .Q(\design_top.TIMER[7] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18892_ (.D(_04470_),
    .Q(\design_top.TIMER[8] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18893_ (.D(_04471_),
    .Q(\design_top.TIMER[9] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18894_ (.D(_04472_),
    .Q(\design_top.TIMER[10] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18895_ (.D(_04473_),
    .Q(\design_top.TIMER[11] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18896_ (.D(_04474_),
    .Q(\design_top.TIMER[12] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18897_ (.D(_04475_),
    .Q(\design_top.TIMER[13] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18898_ (.D(_04476_),
    .Q(\design_top.TIMER[14] ),
    .CLK(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18899_ (.D(_04477_),
    .Q(\design_top.TIMER[15] ),
    .CLK(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18900_ (.D(_04478_),
    .Q(\design_top.TIMER[16] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18901_ (.D(_04479_),
    .Q(\design_top.TIMER[17] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18902_ (.D(_04480_),
    .Q(\design_top.TIMER[18] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18903_ (.D(_04481_),
    .Q(\design_top.TIMER[19] ),
    .CLK(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18904_ (.D(_04482_),
    .Q(\design_top.TIMER[20] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18905_ (.D(_04483_),
    .Q(\design_top.TIMER[21] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18906_ (.D(_04484_),
    .Q(\design_top.TIMER[22] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18907_ (.D(_04485_),
    .Q(\design_top.TIMER[23] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18908_ (.D(_04486_),
    .Q(\design_top.TIMER[24] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18909_ (.D(_04487_),
    .Q(\design_top.TIMER[25] ),
    .CLK(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18910_ (.D(_04488_),
    .Q(\design_top.TIMER[26] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18911_ (.D(_04489_),
    .Q(\design_top.TIMER[27] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18912_ (.D(_04490_),
    .Q(\design_top.TIMER[28] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18913_ (.D(_04491_),
    .Q(\design_top.TIMER[29] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18914_ (.D(_04492_),
    .Q(\design_top.TIMER[30] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18915_ (.D(_04493_),
    .Q(\design_top.TIMER[31] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18916_ (.D(_04494_),
    .Q(\design_top.MEM[10][0] ),
    .CLK(clknet_leaf_253_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18917_ (.D(_04495_),
    .Q(\design_top.MEM[10][1] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18918_ (.D(_04496_),
    .Q(\design_top.MEM[10][2] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18919_ (.D(_04497_),
    .Q(\design_top.MEM[10][3] ),
    .CLK(clknet_leaf_235_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18920_ (.D(_04498_),
    .Q(\design_top.MEM[10][4] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18921_ (.D(_04499_),
    .Q(\design_top.MEM[10][5] ),
    .CLK(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18922_ (.D(_04500_),
    .Q(\design_top.MEM[10][6] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18923_ (.D(_04501_),
    .Q(\design_top.MEM[10][7] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18924_ (.D(_04502_),
    .Q(\design_top.MEM[0][0] ),
    .CLK(clknet_leaf_251_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18925_ (.D(_04503_),
    .Q(\design_top.MEM[0][1] ),
    .CLK(clknet_leaf_251_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18926_ (.D(_04504_),
    .Q(\design_top.MEM[0][2] ),
    .CLK(clknet_leaf_248_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18927_ (.D(_04505_),
    .Q(\design_top.MEM[0][3] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18928_ (.D(_04506_),
    .Q(\design_top.MEM[0][4] ),
    .CLK(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18929_ (.D(_04507_),
    .Q(\design_top.MEM[0][5] ),
    .CLK(clknet_leaf_248_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18930_ (.D(_04508_),
    .Q(\design_top.MEM[0][6] ),
    .CLK(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18931_ (.D(_04509_),
    .Q(\design_top.MEM[0][7] ),
    .CLK(clknet_leaf_235_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18932_ (.D(_04510_),
    .Q(\design_top.uart0.UART_XFIFO[0] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18933_ (.D(_04511_),
    .Q(\design_top.uart0.UART_XFIFO[1] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18934_ (.D(_04512_),
    .Q(\design_top.uart0.UART_XFIFO[2] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18935_ (.D(_04513_),
    .Q(\design_top.uart0.UART_XFIFO[3] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18936_ (.D(_04514_),
    .Q(\design_top.uart0.UART_XFIFO[4] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18937_ (.D(_04515_),
    .Q(\design_top.uart0.UART_XFIFO[5] ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18938_ (.D(_04516_),
    .Q(\design_top.uart0.UART_XFIFO[6] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18939_ (.D(_04517_),
    .Q(\design_top.uart0.UART_XFIFO[7] ),
    .CLK(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18940_ (.D(_04518_),
    .Q(\design_top.uart0.UART_XREQ ),
    .CLK(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18941_ (.D(_04519_),
    .Q(\design_top.uart0.UART_RACK ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18942_ (.D(_04520_),
    .Q(\design_top.IRES[0] ),
    .CLK(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18943_ (.D(_04521_),
    .Q(\design_top.IRES[1] ),
    .CLK(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18944_ (.D(_04522_),
    .Q(\design_top.IRES[2] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18945_ (.D(_04523_),
    .Q(\design_top.IRES[3] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18946_ (.D(_04524_),
    .Q(\design_top.IRES[4] ),
    .CLK(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18947_ (.D(_04525_),
    .Q(\design_top.IRES[5] ),
    .CLK(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18948_ (.D(_04526_),
    .Q(\design_top.IRES[6] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18949_ (.D(_04527_),
    .Q(\design_top.IRES[7] ),
    .CLK(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18950_ (.D(_04528_),
    .Q(\design_top.core0.RESMODE[0] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18951_ (.D(_04529_),
    .Q(\design_top.core0.RESMODE[1] ),
    .CLK(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18952_ (.D(_04530_),
    .Q(\design_top.core0.RESMODE[2] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18953_ (.D(_04531_),
    .Q(\design_top.core0.RESMODE[3] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18954_ (.D(_04532_),
    .Q(_00429_),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18955_ (.D(_04533_),
    .Q(_00430_),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18956_ (.D(_04534_),
    .Q(_00431_),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18957_ (.D(_04535_),
    .Q(_00432_),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18958_ (.D(_04536_),
    .Q(\design_top.uart0.UART_RBAUD[1] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18959_ (.D(_04537_),
    .Q(\design_top.uart0.UART_RBAUD[2] ),
    .CLK(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18960_ (.D(_04538_),
    .Q(\design_top.uart0.UART_RBAUD[4] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18961_ (.D(_04539_),
    .Q(\design_top.uart0.UART_RBAUD[6] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18962_ (.D(_04540_),
    .Q(\design_top.uart0.UART_RBAUD[7] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18963_ (.D(_04541_),
    .Q(\design_top.uart0.UART_RBAUD[9] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18964_ (.D(_04542_),
    .Q(\design_top.uart0.UART_RSTATE[0] ),
    .CLK(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18965_ (.D(_04543_),
    .Q(\design_top.uart0.UART_RSTATE[1] ),
    .CLK(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18966_ (.D(_04544_),
    .Q(\design_top.uart0.UART_RSTATE[2] ),
    .CLK(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18967_ (.D(_04545_),
    .Q(\design_top.uart0.UART_RSTATE[3] ),
    .CLK(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18968_ (.D(_04546_),
    .Q(\design_top.uart0.UART_XSTATE[0] ),
    .CLK(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18969_ (.D(_04547_),
    .Q(\design_top.uart0.UART_XSTATE[1] ),
    .CLK(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18970_ (.D(_04548_),
    .Q(\design_top.uart0.UART_XSTATE[2] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18971_ (.D(_04549_),
    .Q(\design_top.uart0.UART_XSTATE[3] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18972_ (.D(_04550_),
    .Q(\design_top.DACK[0] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18973_ (.D(_04551_),
    .Q(\design_top.DACK[1] ),
    .CLK(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18974_ (.D(_04552_),
    .Q(_00433_),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18975_ (.D(_04553_),
    .Q(_00434_),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18976_ (.D(_04554_),
    .Q(_00435_),
    .CLK(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18977_ (.D(_04555_),
    .Q(_00436_),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18978_ (.D(_04556_),
    .Q(\design_top.uart0.UART_XBAUD[0] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18979_ (.D(_04557_),
    .Q(\design_top.uart0.UART_XBAUD[1] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18980_ (.D(_04558_),
    .Q(\design_top.uart0.UART_XBAUD[2] ),
    .CLK(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18981_ (.D(_04559_),
    .Q(\design_top.uart0.UART_XBAUD[3] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18982_ (.D(_04560_),
    .Q(\design_top.uart0.UART_XBAUD[4] ),
    .CLK(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18983_ (.D(_04561_),
    .Q(\design_top.uart0.UART_XBAUD[5] ),
    .CLK(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18984_ (.D(_04562_),
    .Q(\design_top.uart0.UART_XBAUD[6] ),
    .CLK(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18985_ (.D(_04563_),
    .Q(\design_top.uart0.UART_XBAUD[7] ),
    .CLK(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18986_ (.D(_04564_),
    .Q(\design_top.uart0.UART_XBAUD[8] ),
    .CLK(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18987_ (.D(_04565_),
    .Q(\design_top.uart0.UART_XBAUD[9] ),
    .CLK(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18988_ (.D(_04566_),
    .Q(\design_top.uart0.UART_XBAUD[10] ),
    .CLK(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18989_ (.D(_04567_),
    .Q(\design_top.uart0.UART_XBAUD[11] ),
    .CLK(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18990_ (.D(_04568_),
    .Q(\design_top.uart0.UART_XBAUD[12] ),
    .CLK(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18991_ (.D(_04569_),
    .Q(\design_top.uart0.UART_XBAUD[13] ),
    .CLK(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18992_ (.D(_04570_),
    .Q(\design_top.uart0.UART_XBAUD[14] ),
    .CLK(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18993_ (.D(_04571_),
    .Q(\design_top.uart0.UART_XBAUD[15] ),
    .CLK(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18994_ (.D(_04572_),
    .Q(\design_top.uart0.UART_RBAUD[0] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18995_ (.D(_04573_),
    .Q(\design_top.uart0.UART_RBAUD[3] ),
    .CLK(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18996_ (.D(_04574_),
    .Q(\design_top.uart0.UART_RBAUD[5] ),
    .CLK(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18997_ (.D(_04575_),
    .Q(\design_top.uart0.UART_RBAUD[8] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18998_ (.D(_04576_),
    .Q(\design_top.uart0.UART_RBAUD[10] ),
    .CLK(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _18999_ (.D(_04577_),
    .Q(\design_top.uart0.UART_RBAUD[11] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19000_ (.D(_04578_),
    .Q(\design_top.uart0.UART_RBAUD[12] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19001_ (.D(_04579_),
    .Q(\design_top.uart0.UART_RBAUD[13] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19002_ (.D(_04580_),
    .Q(\design_top.uart0.UART_RBAUD[14] ),
    .CLK(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19003_ (.D(_04581_),
    .Q(\design_top.uart0.UART_RBAUD[15] ),
    .CLK(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19004_ (.D(_04582_),
    .Q(io_out[16]),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19005_ (.D(_04583_),
    .Q(io_out[17]),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19006_ (.D(_04584_),
    .Q(\design_top.MEM[12][16] ),
    .CLK(clknet_leaf_269_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19007_ (.D(_04585_),
    .Q(\design_top.MEM[12][17] ),
    .CLK(clknet_leaf_267_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19008_ (.D(_04586_),
    .Q(\design_top.MEM[12][18] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19009_ (.D(_04587_),
    .Q(\design_top.MEM[12][19] ),
    .CLK(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19010_ (.D(_04588_),
    .Q(\design_top.MEM[12][20] ),
    .CLK(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19011_ (.D(_04589_),
    .Q(\design_top.MEM[12][21] ),
    .CLK(clknet_leaf_269_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19012_ (.D(_04590_),
    .Q(\design_top.MEM[12][22] ),
    .CLK(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19013_ (.D(_04591_),
    .Q(\design_top.MEM[12][23] ),
    .CLK(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19014_ (.D(_04592_),
    .Q(\design_top.core0.FLUSH[0] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19015_ (.D(_04593_),
    .Q(\design_top.core0.FLUSH[1] ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19016_ (.D(_04594_),
    .Q(io_out[18]),
    .CLK(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19017_ (.D(_04595_),
    .Q(io_out[19]),
    .CLK(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19018_ (.D(_04596_),
    .Q(\design_top.IADDR[4] ),
    .CLK(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19019_ (.D(_04597_),
    .Q(\design_top.IADDR[5] ),
    .CLK(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19020_ (.D(_04598_),
    .Q(\design_top.IADDR[6] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19021_ (.D(_04599_),
    .Q(\design_top.IADDR[7] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19022_ (.D(_04600_),
    .Q(\design_top.IADDR[8] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19023_ (.D(_04601_),
    .Q(\design_top.IADDR[9] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19024_ (.D(_04602_),
    .Q(\design_top.IADDR[10] ),
    .CLK(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19025_ (.D(_04603_),
    .Q(\design_top.IADDR[11] ),
    .CLK(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19026_ (.D(_04604_),
    .Q(\design_top.IADDR[12] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19027_ (.D(_04605_),
    .Q(\design_top.IADDR[13] ),
    .CLK(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19028_ (.D(_04606_),
    .Q(\design_top.IADDR[14] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19029_ (.D(_04607_),
    .Q(\design_top.IADDR[15] ),
    .CLK(clknet_leaf_172_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19030_ (.D(_04608_),
    .Q(\design_top.IADDR[16] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19031_ (.D(_04609_),
    .Q(\design_top.IADDR[17] ),
    .CLK(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19032_ (.D(_04610_),
    .Q(\design_top.IADDR[18] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19033_ (.D(_04611_),
    .Q(\design_top.IADDR[19] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19034_ (.D(_04612_),
    .Q(\design_top.IADDR[20] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19035_ (.D(_04613_),
    .Q(\design_top.IADDR[21] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19036_ (.D(_04614_),
    .Q(\design_top.IADDR[22] ),
    .CLK(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19037_ (.D(_04615_),
    .Q(\design_top.IADDR[23] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19038_ (.D(_04616_),
    .Q(\design_top.IADDR[24] ),
    .CLK(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19039_ (.D(_04617_),
    .Q(\design_top.IADDR[25] ),
    .CLK(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19040_ (.D(_04618_),
    .Q(\design_top.IADDR[26] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19041_ (.D(_04619_),
    .Q(\design_top.IADDR[27] ),
    .CLK(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19042_ (.D(_04620_),
    .Q(\design_top.IADDR[28] ),
    .CLK(clknet_leaf_172_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19043_ (.D(_04621_),
    .Q(\design_top.IADDR[29] ),
    .CLK(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19044_ (.D(_04622_),
    .Q(\design_top.IADDR[30] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19045_ (.D(_04623_),
    .Q(\design_top.IADDR[31] ),
    .CLK(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19046_ (.D(_04624_),
    .Q(\design_top.core0.XIDATA[7] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19047_ (.D(_04625_),
    .Q(\design_top.core0.XIDATA[8] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19048_ (.D(_04626_),
    .Q(\design_top.core0.XIDATA[9] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19049_ (.D(_04627_),
    .Q(\design_top.core0.XIDATA[10] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19050_ (.D(_04628_),
    .Q(\design_top.core0.FCT3[0] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19051_ (.D(_04629_),
    .Q(\design_top.core0.FCT3[1] ),
    .CLK(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19052_ (.D(_04630_),
    .Q(\design_top.core0.FCT3[2] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19053_ (.D(_04631_),
    .Q(\design_top.core0.S1PTR[0] ),
    .CLK(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19054_ (.D(_04632_),
    .Q(\design_top.core0.S1PTR[1] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19055_ (.D(_04633_),
    .Q(\design_top.core0.S1PTR[2] ),
    .CLK(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19056_ (.D(_04634_),
    .Q(\design_top.core0.S1PTR[3] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19057_ (.D(_04635_),
    .Q(\design_top.core0.S2PTR[0] ),
    .CLK(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19058_ (.D(_04636_),
    .Q(\design_top.core0.S2PTR[1] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19059_ (.D(_04637_),
    .Q(\design_top.core0.S2PTR[2] ),
    .CLK(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19060_ (.D(_04638_),
    .Q(\design_top.core0.S2PTR[3] ),
    .CLK(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19061_ (.D(_04639_),
    .Q(\design_top.core0.FCT7[5] ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19062_ (.D(_04640_),
    .Q(\design_top.core0.XLUI ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19063_ (.D(_04641_),
    .Q(\design_top.core0.XAUIPC ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19064_ (.D(_04642_),
    .Q(\design_top.core0.XJAL ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19065_ (.D(_04643_),
    .Q(\design_top.core0.XJALR ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19066_ (.D(_04644_),
    .Q(\design_top.core0.XBCC ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19067_ (.D(_04645_),
    .Q(\design_top.core0.XLCC ),
    .CLK(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19068_ (.D(_04646_),
    .Q(\design_top.core0.XSCC ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19069_ (.D(_04647_),
    .Q(\design_top.core0.XMCC ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19070_ (.D(_04648_),
    .Q(\design_top.core0.XRCC ),
    .CLK(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19071_ (.D(_04649_),
    .Q(\design_top.core0.SIMM[12] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19072_ (.D(_04650_),
    .Q(\design_top.core0.SIMM[13] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19073_ (.D(_04651_),
    .Q(\design_top.core0.SIMM[14] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19074_ (.D(_04652_),
    .Q(\design_top.core0.SIMM[15] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19075_ (.D(_04653_),
    .Q(\design_top.core0.SIMM[16] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19076_ (.D(_04654_),
    .Q(\design_top.core0.SIMM[17] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19077_ (.D(_04655_),
    .Q(\design_top.core0.SIMM[18] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19078_ (.D(_04656_),
    .Q(\design_top.core0.SIMM[19] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19079_ (.D(_04657_),
    .Q(\design_top.core0.SIMM[20] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19080_ (.D(_04658_),
    .Q(\design_top.core0.SIMM[21] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19081_ (.D(_04659_),
    .Q(\design_top.core0.SIMM[22] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19082_ (.D(_04660_),
    .Q(\design_top.core0.SIMM[23] ),
    .CLK(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19083_ (.D(_04661_),
    .Q(\design_top.core0.SIMM[24] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19084_ (.D(_04662_),
    .Q(\design_top.core0.SIMM[25] ),
    .CLK(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19085_ (.D(_04663_),
    .Q(\design_top.core0.SIMM[26] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19086_ (.D(_04664_),
    .Q(\design_top.core0.SIMM[27] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19087_ (.D(_04665_),
    .Q(\design_top.core0.SIMM[28] ),
    .CLK(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19088_ (.D(_04666_),
    .Q(\design_top.core0.SIMM[29] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19089_ (.D(_04667_),
    .Q(\design_top.core0.SIMM[30] ),
    .CLK(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19090_ (.D(_04668_),
    .Q(\design_top.core0.SIMM[31] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19091_ (.D(_04669_),
    .Q(\design_top.core0.SIMM[0] ),
    .CLK(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19092_ (.D(_04670_),
    .Q(\design_top.core0.SIMM[1] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19093_ (.D(_04671_),
    .Q(\design_top.core0.SIMM[2] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19094_ (.D(_04672_),
    .Q(\design_top.core0.SIMM[3] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19095_ (.D(_04673_),
    .Q(\design_top.core0.SIMM[4] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19096_ (.D(_04674_),
    .Q(\design_top.core0.SIMM[5] ),
    .CLK(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19097_ (.D(_04675_),
    .Q(\design_top.core0.SIMM[6] ),
    .CLK(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19098_ (.D(_04676_),
    .Q(\design_top.core0.SIMM[7] ),
    .CLK(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19099_ (.D(_04677_),
    .Q(\design_top.core0.SIMM[8] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19100_ (.D(_04678_),
    .Q(\design_top.core0.SIMM[9] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19101_ (.D(_04679_),
    .Q(\design_top.core0.SIMM[10] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19102_ (.D(_04680_),
    .Q(\design_top.core0.SIMM[11] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19103_ (.D(_04681_),
    .Q(\design_top.core0.UIMM[12] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19104_ (.D(_04682_),
    .Q(\design_top.core0.UIMM[13] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19105_ (.D(_04683_),
    .Q(\design_top.core0.UIMM[14] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19106_ (.D(_04684_),
    .Q(\design_top.core0.UIMM[15] ),
    .CLK(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19107_ (.D(_04685_),
    .Q(\design_top.core0.UIMM[16] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19108_ (.D(_04686_),
    .Q(\design_top.core0.UIMM[17] ),
    .CLK(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19109_ (.D(_04687_),
    .Q(\design_top.core0.UIMM[18] ),
    .CLK(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19110_ (.D(_04688_),
    .Q(\design_top.core0.UIMM[19] ),
    .CLK(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19111_ (.D(_04689_),
    .Q(\design_top.core0.UIMM[20] ),
    .CLK(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19112_ (.D(_04690_),
    .Q(\design_top.core0.UIMM[21] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19113_ (.D(_04691_),
    .Q(\design_top.core0.UIMM[22] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19114_ (.D(_04692_),
    .Q(\design_top.core0.UIMM[23] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19115_ (.D(_04693_),
    .Q(\design_top.core0.UIMM[24] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19116_ (.D(_04694_),
    .Q(\design_top.core0.UIMM[25] ),
    .CLK(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19117_ (.D(_04695_),
    .Q(\design_top.core0.UIMM[26] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19118_ (.D(_04696_),
    .Q(\design_top.core0.UIMM[27] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19119_ (.D(_04697_),
    .Q(\design_top.core0.UIMM[28] ),
    .CLK(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19120_ (.D(_04698_),
    .Q(\design_top.core0.UIMM[29] ),
    .CLK(clknet_5_26_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19121_ (.D(_04699_),
    .Q(\design_top.core0.UIMM[30] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19122_ (.D(_04700_),
    .Q(\design_top.core0.UIMM[31] ),
    .CLK(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19123_ (.D(_04701_),
    .Q(\design_top.MEM[12][24] ),
    .CLK(clknet_leaf_29_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19124_ (.D(_04702_),
    .Q(\design_top.MEM[12][25] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19125_ (.D(_04703_),
    .Q(\design_top.MEM[12][26] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19126_ (.D(_04704_),
    .Q(\design_top.MEM[12][27] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19127_ (.D(_04705_),
    .Q(\design_top.MEM[12][28] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19128_ (.D(_04706_),
    .Q(\design_top.MEM[12][29] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19129_ (.D(_04707_),
    .Q(\design_top.MEM[12][30] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19130_ (.D(_04708_),
    .Q(\design_top.MEM[12][31] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19131_ (.D(_04709_),
    .Q(\design_top.MEM[12][8] ),
    .CLK(clknet_leaf_289_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19132_ (.D(_04710_),
    .Q(\design_top.MEM[12][9] ),
    .CLK(clknet_leaf_295_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19133_ (.D(_04711_),
    .Q(\design_top.MEM[12][10] ),
    .CLK(clknet_leaf_290_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19134_ (.D(_04712_),
    .Q(\design_top.MEM[12][11] ),
    .CLK(clknet_leaf_300_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19135_ (.D(_04713_),
    .Q(\design_top.MEM[12][12] ),
    .CLK(clknet_leaf_300_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19136_ (.D(_04714_),
    .Q(\design_top.MEM[12][13] ),
    .CLK(clknet_leaf_295_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19137_ (.D(_04715_),
    .Q(\design_top.MEM[12][14] ),
    .CLK(clknet_leaf_300_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19138_ (.D(_04716_),
    .Q(\design_top.MEM[12][15] ),
    .CLK(clknet_leaf_301_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19139_ (.D(_04717_),
    .Q(\design_top.MEM[11][24] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19140_ (.D(_04718_),
    .Q(\design_top.MEM[11][25] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19141_ (.D(_04719_),
    .Q(\design_top.MEM[11][26] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19142_ (.D(_04720_),
    .Q(\design_top.MEM[11][27] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19143_ (.D(_04721_),
    .Q(\design_top.MEM[11][28] ),
    .CLK(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19144_ (.D(_04722_),
    .Q(\design_top.MEM[11][29] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19145_ (.D(_04723_),
    .Q(\design_top.MEM[11][30] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19146_ (.D(_04724_),
    .Q(\design_top.MEM[11][31] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19147_ (.D(_04725_),
    .Q(\design_top.IOMUX[3][0] ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19148_ (.D(_04726_),
    .Q(\design_top.IOMUX[3][1] ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19149_ (.D(_04727_),
    .Q(\design_top.IOMUX[3][2] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19150_ (.D(_04728_),
    .Q(\design_top.IOMUX[3][3] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19151_ (.D(_04729_),
    .Q(\design_top.IOMUX[3][4] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19152_ (.D(_04730_),
    .Q(\design_top.IOMUX[3][5] ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19153_ (.D(_04731_),
    .Q(\design_top.IOMUX[3][6] ),
    .CLK(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19154_ (.D(_04732_),
    .Q(\design_top.IOMUX[3][7] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19155_ (.D(_04733_),
    .Q(\design_top.IOMUX[3][8] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19156_ (.D(_04734_),
    .Q(\design_top.IOMUX[3][9] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19157_ (.D(_04735_),
    .Q(\design_top.IOMUX[3][10] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19158_ (.D(_04736_),
    .Q(\design_top.IOMUX[3][11] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19159_ (.D(_04737_),
    .Q(\design_top.IOMUX[3][12] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19160_ (.D(_04738_),
    .Q(\design_top.IOMUX[3][13] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19161_ (.D(_04739_),
    .Q(\design_top.IOMUX[3][14] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19162_ (.D(_04740_),
    .Q(\design_top.IOMUX[3][15] ),
    .CLK(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19163_ (.D(_04741_),
    .Q(\design_top.IOMUX[3][16] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19164_ (.D(_04742_),
    .Q(\design_top.IOMUX[3][17] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19165_ (.D(_04743_),
    .Q(\design_top.IOMUX[3][18] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19166_ (.D(_04744_),
    .Q(\design_top.IOMUX[3][19] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19167_ (.D(_04745_),
    .Q(\design_top.IOMUX[3][20] ),
    .CLK(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19168_ (.D(_04746_),
    .Q(\design_top.IOMUX[3][21] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19169_ (.D(_04747_),
    .Q(\design_top.IOMUX[3][22] ),
    .CLK(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19170_ (.D(_04748_),
    .Q(\design_top.IOMUX[3][23] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19171_ (.D(_04749_),
    .Q(\design_top.IOMUX[3][24] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19172_ (.D(_04750_),
    .Q(\design_top.IOMUX[3][25] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19173_ (.D(_04751_),
    .Q(\design_top.IOMUX[3][26] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19174_ (.D(_04752_),
    .Q(\design_top.IOMUX[3][27] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19175_ (.D(_04753_),
    .Q(\design_top.IOMUX[3][28] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19176_ (.D(_04754_),
    .Q(\design_top.IOMUX[3][29] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19177_ (.D(_04755_),
    .Q(\design_top.IOMUX[3][30] ),
    .CLK(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19178_ (.D(_04756_),
    .Q(\design_top.IOMUX[3][31] ),
    .CLK(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19179_ (.D(_04757_),
    .Q(\design_top.MEM[11][16] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19180_ (.D(_04758_),
    .Q(\design_top.MEM[11][17] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19181_ (.D(_04759_),
    .Q(\design_top.MEM[11][18] ),
    .CLK(clknet_leaf_292_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19182_ (.D(_04760_),
    .Q(\design_top.MEM[11][19] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19183_ (.D(_04761_),
    .Q(\design_top.MEM[11][20] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19184_ (.D(_04762_),
    .Q(\design_top.MEM[11][21] ),
    .CLK(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19185_ (.D(_04763_),
    .Q(\design_top.MEM[11][22] ),
    .CLK(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19186_ (.D(_04764_),
    .Q(\design_top.MEM[11][23] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19187_ (.D(_04765_),
    .Q(\design_top.MEM[13][8] ),
    .CLK(clknet_leaf_289_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19188_ (.D(_04766_),
    .Q(\design_top.MEM[13][9] ),
    .CLK(clknet_leaf_295_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19189_ (.D(_04767_),
    .Q(\design_top.MEM[13][10] ),
    .CLK(clknet_leaf_290_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19190_ (.D(_04768_),
    .Q(\design_top.MEM[13][11] ),
    .CLK(clknet_leaf_301_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19191_ (.D(_04769_),
    .Q(\design_top.MEM[13][12] ),
    .CLK(clknet_leaf_300_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19192_ (.D(_04770_),
    .Q(\design_top.MEM[13][13] ),
    .CLK(clknet_leaf_295_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19193_ (.D(_04771_),
    .Q(\design_top.MEM[13][14] ),
    .CLK(clknet_leaf_300_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19194_ (.D(_04772_),
    .Q(\design_top.MEM[13][15] ),
    .CLK(clknet_leaf_301_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19195_ (.D(_04773_),
    .Q(\design_top.MEM[2][16] ),
    .CLK(clknet_leaf_278_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19196_ (.D(_04774_),
    .Q(\design_top.MEM[2][17] ),
    .CLK(clknet_leaf_283_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19197_ (.D(_04775_),
    .Q(\design_top.MEM[2][18] ),
    .CLK(clknet_leaf_291_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19198_ (.D(_04776_),
    .Q(\design_top.MEM[2][19] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19199_ (.D(_04777_),
    .Q(\design_top.MEM[2][20] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19200_ (.D(_04778_),
    .Q(\design_top.MEM[2][21] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19201_ (.D(_04779_),
    .Q(\design_top.MEM[2][22] ),
    .CLK(clknet_leaf_277_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19202_ (.D(_04780_),
    .Q(\design_top.MEM[2][23] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19203_ (.D(_04781_),
    .Q(\design_top.MEM[2][8] ),
    .CLK(clknet_leaf_307_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19204_ (.D(_04782_),
    .Q(\design_top.MEM[2][9] ),
    .CLK(clknet_leaf_307_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19205_ (.D(_04783_),
    .Q(\design_top.MEM[2][10] ),
    .CLK(clknet_leaf_288_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19206_ (.D(_04784_),
    .Q(\design_top.MEM[2][11] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19207_ (.D(_04785_),
    .Q(\design_top.MEM[2][12] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19208_ (.D(_04786_),
    .Q(\design_top.MEM[2][13] ),
    .CLK(clknet_leaf_307_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19209_ (.D(_04787_),
    .Q(\design_top.MEM[2][14] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19210_ (.D(_04788_),
    .Q(\design_top.MEM[2][15] ),
    .CLK(clknet_leaf_302_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19211_ (.D(_04789_),
    .Q(\design_top.MEM[29][24] ),
    .CLK(clknet_leaf_310_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19212_ (.D(_04790_),
    .Q(\design_top.MEM[29][25] ),
    .CLK(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19213_ (.D(_04791_),
    .Q(\design_top.MEM[29][26] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19214_ (.D(_04792_),
    .Q(\design_top.MEM[29][27] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19215_ (.D(_04793_),
    .Q(\design_top.MEM[29][28] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19216_ (.D(_04794_),
    .Q(\design_top.MEM[29][29] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19217_ (.D(_04795_),
    .Q(\design_top.MEM[29][30] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19218_ (.D(_04796_),
    .Q(\design_top.MEM[29][31] ),
    .CLK(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19219_ (.D(_04797_),
    .Q(\design_top.MEM[29][16] ),
    .CLK(clknet_leaf_283_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19220_ (.D(_04798_),
    .Q(\design_top.MEM[29][17] ),
    .CLK(clknet_leaf_282_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19221_ (.D(_04799_),
    .Q(\design_top.MEM[29][18] ),
    .CLK(clknet_leaf_291_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19222_ (.D(_04800_),
    .Q(\design_top.MEM[29][19] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19223_ (.D(_04801_),
    .Q(\design_top.MEM[29][20] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19224_ (.D(_04802_),
    .Q(\design_top.MEM[29][21] ),
    .CLK(clknet_leaf_278_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19225_ (.D(_04803_),
    .Q(\design_top.MEM[29][22] ),
    .CLK(clknet_leaf_39_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19226_ (.D(_04804_),
    .Q(\design_top.MEM[29][23] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19227_ (.D(_04805_),
    .Q(\design_top.MEM[23][8] ),
    .CLK(clknet_leaf_312_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19228_ (.D(_04806_),
    .Q(\design_top.MEM[23][9] ),
    .CLK(clknet_leaf_312_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19229_ (.D(_04807_),
    .Q(\design_top.MEM[23][10] ),
    .CLK(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19230_ (.D(_04808_),
    .Q(\design_top.MEM[23][11] ),
    .CLK(clknet_leaf_319_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19231_ (.D(_04809_),
    .Q(\design_top.MEM[23][12] ),
    .CLK(clknet_leaf_318_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19232_ (.D(_04810_),
    .Q(\design_top.MEM[23][13] ),
    .CLK(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19233_ (.D(_04811_),
    .Q(\design_top.MEM[23][14] ),
    .CLK(clknet_leaf_318_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19234_ (.D(_04812_),
    .Q(\design_top.MEM[23][15] ),
    .CLK(clknet_leaf_314_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19235_ (.D(_04813_),
    .Q(\design_top.MEM[29][8] ),
    .CLK(clknet_leaf_309_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19236_ (.D(_04814_),
    .Q(\design_top.MEM[29][9] ),
    .CLK(clknet_leaf_309_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19237_ (.D(_04815_),
    .Q(\design_top.MEM[29][10] ),
    .CLK(clknet_leaf_310_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19238_ (.D(_04816_),
    .Q(\design_top.MEM[29][11] ),
    .CLK(clknet_leaf_316_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19239_ (.D(_04817_),
    .Q(\design_top.MEM[29][12] ),
    .CLK(clknet_leaf_316_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19240_ (.D(_04818_),
    .Q(\design_top.MEM[29][13] ),
    .CLK(clknet_leaf_315_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19241_ (.D(_04819_),
    .Q(\design_top.MEM[29][14] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19242_ (.D(_04820_),
    .Q(\design_top.MEM[29][15] ),
    .CLK(clknet_leaf_315_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19243_ (.D(_04821_),
    .Q(\design_top.MEM[28][24] ),
    .CLK(clknet_leaf_286_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19244_ (.D(_04822_),
    .Q(\design_top.MEM[28][25] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19245_ (.D(_04823_),
    .Q(\design_top.MEM[28][26] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19246_ (.D(_04824_),
    .Q(\design_top.MEM[28][27] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19247_ (.D(_04825_),
    .Q(\design_top.MEM[28][28] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19248_ (.D(_04826_),
    .Q(\design_top.MEM[28][29] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19249_ (.D(_04827_),
    .Q(\design_top.MEM[28][30] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19250_ (.D(_04828_),
    .Q(\design_top.MEM[28][31] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19251_ (.D(_04829_),
    .Q(\design_top.MEM[28][16] ),
    .CLK(clknet_leaf_283_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19252_ (.D(_04830_),
    .Q(\design_top.MEM[28][17] ),
    .CLK(clknet_leaf_282_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19253_ (.D(_04831_),
    .Q(\design_top.MEM[28][18] ),
    .CLK(clknet_leaf_282_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19254_ (.D(_04832_),
    .Q(\design_top.MEM[28][19] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19255_ (.D(_04833_),
    .Q(\design_top.MEM[28][20] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19256_ (.D(_04834_),
    .Q(\design_top.MEM[28][21] ),
    .CLK(clknet_leaf_278_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19257_ (.D(_04835_),
    .Q(\design_top.MEM[28][22] ),
    .CLK(clknet_leaf_39_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19258_ (.D(_04836_),
    .Q(\design_top.MEM[28][23] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19259_ (.D(_04837_),
    .Q(\design_top.MEM[28][8] ),
    .CLK(clknet_leaf_309_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19260_ (.D(_04838_),
    .Q(\design_top.MEM[28][9] ),
    .CLK(clknet_leaf_309_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19261_ (.D(_04839_),
    .Q(\design_top.MEM[28][10] ),
    .CLK(clknet_leaf_310_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19262_ (.D(_04840_),
    .Q(\design_top.MEM[28][11] ),
    .CLK(clknet_leaf_315_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19263_ (.D(_04841_),
    .Q(\design_top.MEM[28][12] ),
    .CLK(clknet_leaf_316_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19264_ (.D(_04842_),
    .Q(\design_top.MEM[28][13] ),
    .CLK(clknet_leaf_315_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19265_ (.D(_04843_),
    .Q(\design_top.MEM[28][14] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19266_ (.D(_04844_),
    .Q(\design_top.MEM[28][15] ),
    .CLK(clknet_leaf_315_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19267_ (.D(_04845_),
    .Q(\design_top.MEM[27][24] ),
    .CLK(clknet_leaf_311_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19268_ (.D(_04846_),
    .Q(\design_top.MEM[27][25] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19269_ (.D(_04847_),
    .Q(\design_top.MEM[27][26] ),
    .CLK(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19270_ (.D(_04848_),
    .Q(\design_top.MEM[27][27] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19271_ (.D(_04849_),
    .Q(\design_top.MEM[27][28] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19272_ (.D(_04850_),
    .Q(\design_top.MEM[27][29] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19273_ (.D(_04851_),
    .Q(\design_top.MEM[27][30] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19274_ (.D(_04852_),
    .Q(\design_top.MEM[27][31] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19275_ (.D(_04853_),
    .Q(\design_top.MEM[27][16] ),
    .CLK(clknet_leaf_284_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19276_ (.D(_04854_),
    .Q(\design_top.MEM[27][17] ),
    .CLK(clknet_leaf_282_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19277_ (.D(_04855_),
    .Q(\design_top.MEM[27][18] ),
    .CLK(clknet_leaf_290_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19278_ (.D(_04856_),
    .Q(\design_top.MEM[27][19] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19279_ (.D(_04857_),
    .Q(\design_top.MEM[27][20] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19280_ (.D(_04858_),
    .Q(\design_top.MEM[27][21] ),
    .CLK(clknet_leaf_284_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19281_ (.D(_04859_),
    .Q(\design_top.MEM[27][22] ),
    .CLK(clknet_leaf_39_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19282_ (.D(_04860_),
    .Q(\design_top.MEM[27][23] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19283_ (.D(_04861_),
    .Q(\design_top.MEM[27][8] ),
    .CLK(clknet_leaf_312_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19284_ (.D(_04862_),
    .Q(\design_top.MEM[27][9] ),
    .CLK(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19285_ (.D(_04863_),
    .Q(\design_top.MEM[27][10] ),
    .CLK(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19286_ (.D(_04864_),
    .Q(\design_top.MEM[27][11] ),
    .CLK(clknet_leaf_319_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19287_ (.D(_04865_),
    .Q(\design_top.MEM[27][12] ),
    .CLK(clknet_leaf_318_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19288_ (.D(_04866_),
    .Q(\design_top.MEM[27][13] ),
    .CLK(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19289_ (.D(_04867_),
    .Q(\design_top.MEM[27][14] ),
    .CLK(clknet_leaf_318_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19290_ (.D(_04868_),
    .Q(\design_top.MEM[27][15] ),
    .CLK(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19291_ (.D(_04869_),
    .Q(\design_top.MEM[26][24] ),
    .CLK(clknet_leaf_311_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19292_ (.D(_04870_),
    .Q(\design_top.MEM[26][25] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19293_ (.D(_04871_),
    .Q(\design_top.MEM[26][26] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19294_ (.D(_04872_),
    .Q(\design_top.MEM[26][27] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19295_ (.D(_04873_),
    .Q(\design_top.MEM[26][28] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19296_ (.D(_04874_),
    .Q(\design_top.MEM[26][29] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19297_ (.D(_04875_),
    .Q(\design_top.MEM[26][30] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19298_ (.D(_04876_),
    .Q(\design_top.MEM[26][31] ),
    .CLK(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19299_ (.D(_04877_),
    .Q(\design_top.MEM[26][16] ),
    .CLK(clknet_leaf_283_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19300_ (.D(_04878_),
    .Q(\design_top.MEM[26][17] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19301_ (.D(_04879_),
    .Q(\design_top.MEM[26][18] ),
    .CLK(clknet_leaf_291_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19302_ (.D(_04880_),
    .Q(\design_top.MEM[26][19] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19303_ (.D(_04881_),
    .Q(\design_top.MEM[26][20] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19304_ (.D(_04882_),
    .Q(\design_top.MEM[26][21] ),
    .CLK(clknet_leaf_284_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19305_ (.D(_04883_),
    .Q(\design_top.MEM[26][22] ),
    .CLK(clknet_leaf_39_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19306_ (.D(_04884_),
    .Q(\design_top.MEM[26][23] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19307_ (.D(_04885_),
    .Q(\design_top.MEM[22][24] ),
    .CLK(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19308_ (.D(_04886_),
    .Q(\design_top.MEM[22][25] ),
    .CLK(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19309_ (.D(_04887_),
    .Q(\design_top.MEM[22][26] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19310_ (.D(_04888_),
    .Q(\design_top.MEM[22][27] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19311_ (.D(_04889_),
    .Q(\design_top.MEM[22][28] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19312_ (.D(_04890_),
    .Q(\design_top.MEM[22][29] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19313_ (.D(_04891_),
    .Q(\design_top.MEM[22][30] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19314_ (.D(_04892_),
    .Q(\design_top.MEM[22][31] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19315_ (.D(_04893_),
    .Q(\design_top.MEM[22][16] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19316_ (.D(_04894_),
    .Q(\design_top.MEM[22][17] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19317_ (.D(_04895_),
    .Q(\design_top.MEM[22][18] ),
    .CLK(clknet_leaf_288_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19318_ (.D(_04896_),
    .Q(\design_top.MEM[22][19] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19319_ (.D(_04897_),
    .Q(\design_top.MEM[22][20] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19320_ (.D(_04898_),
    .Q(\design_top.MEM[22][21] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19321_ (.D(_04899_),
    .Q(\design_top.MEM[22][22] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19322_ (.D(_04900_),
    .Q(\design_top.MEM[22][23] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19323_ (.D(_04901_),
    .Q(\design_top.MEM[26][8] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19324_ (.D(_04902_),
    .Q(\design_top.MEM[26][9] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19325_ (.D(_04903_),
    .Q(\design_top.MEM[26][10] ),
    .CLK(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19326_ (.D(_04904_),
    .Q(\design_top.MEM[26][11] ),
    .CLK(clknet_leaf_318_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19327_ (.D(_04905_),
    .Q(\design_top.MEM[26][12] ),
    .CLK(clknet_leaf_321_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19328_ (.D(_04906_),
    .Q(\design_top.MEM[26][13] ),
    .CLK(clknet_leaf_320_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19329_ (.D(_04907_),
    .Q(\design_top.MEM[26][14] ),
    .CLK(clknet_leaf_322_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19330_ (.D(_04908_),
    .Q(\design_top.MEM[26][15] ),
    .CLK(clknet_leaf_320_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19331_ (.D(_04909_),
    .Q(\design_top.MEM[25][24] ),
    .CLK(clknet_leaf_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19332_ (.D(_04910_),
    .Q(\design_top.MEM[25][25] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19333_ (.D(_04911_),
    .Q(\design_top.MEM[25][26] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19334_ (.D(_04912_),
    .Q(\design_top.MEM[25][27] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19335_ (.D(_04913_),
    .Q(\design_top.MEM[25][28] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19336_ (.D(_04914_),
    .Q(\design_top.MEM[25][29] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19337_ (.D(_04915_),
    .Q(\design_top.MEM[25][30] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19338_ (.D(_04916_),
    .Q(\design_top.MEM[25][31] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19339_ (.D(_04917_),
    .Q(\design_top.MEM[25][16] ),
    .CLK(clknet_leaf_284_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19340_ (.D(_04918_),
    .Q(\design_top.MEM[25][17] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19341_ (.D(_04919_),
    .Q(\design_top.MEM[25][18] ),
    .CLK(clknet_leaf_288_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19342_ (.D(_04920_),
    .Q(\design_top.MEM[25][19] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19343_ (.D(_04921_),
    .Q(\design_top.MEM[25][20] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19344_ (.D(_04922_),
    .Q(\design_top.MEM[25][21] ),
    .CLK(clknet_leaf_39_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19345_ (.D(_04923_),
    .Q(\design_top.MEM[25][22] ),
    .CLK(clknet_leaf_39_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19346_ (.D(_04924_),
    .Q(\design_top.MEM[25][23] ),
    .CLK(clknet_leaf_39_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19347_ (.D(_04925_),
    .Q(\design_top.MEM[25][8] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19348_ (.D(_04926_),
    .Q(\design_top.MEM[25][9] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19349_ (.D(_04927_),
    .Q(\design_top.MEM[25][10] ),
    .CLK(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19350_ (.D(_04928_),
    .Q(\design_top.MEM[25][11] ),
    .CLK(clknet_leaf_319_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19351_ (.D(_04929_),
    .Q(\design_top.MEM[25][12] ),
    .CLK(clknet_leaf_321_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19352_ (.D(_04930_),
    .Q(\design_top.MEM[25][13] ),
    .CLK(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19353_ (.D(_04931_),
    .Q(\design_top.MEM[25][14] ),
    .CLK(clknet_leaf_322_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19354_ (.D(_04932_),
    .Q(\design_top.MEM[25][15] ),
    .CLK(clknet_leaf_320_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19355_ (.D(_04933_),
    .Q(\design_top.MEM[24][24] ),
    .CLK(clknet_leaf_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19356_ (.D(_04934_),
    .Q(\design_top.MEM[24][25] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19357_ (.D(_04935_),
    .Q(\design_top.MEM[24][26] ),
    .CLK(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19358_ (.D(_04936_),
    .Q(\design_top.MEM[24][27] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19359_ (.D(_04937_),
    .Q(\design_top.MEM[24][28] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19360_ (.D(_04938_),
    .Q(\design_top.MEM[24][29] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19361_ (.D(_04939_),
    .Q(\design_top.MEM[24][30] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19362_ (.D(_04940_),
    .Q(\design_top.MEM[24][31] ),
    .CLK(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19363_ (.D(_04941_),
    .Q(\design_top.MEM[24][16] ),
    .CLK(clknet_leaf_284_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19364_ (.D(_04942_),
    .Q(\design_top.MEM[24][17] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19365_ (.D(_04943_),
    .Q(\design_top.MEM[24][18] ),
    .CLK(clknet_leaf_287_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19366_ (.D(_04944_),
    .Q(\design_top.MEM[24][19] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19367_ (.D(_04945_),
    .Q(\design_top.MEM[24][20] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19368_ (.D(_04946_),
    .Q(\design_top.MEM[24][21] ),
    .CLK(clknet_leaf_39_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19369_ (.D(_04947_),
    .Q(\design_top.MEM[24][22] ),
    .CLK(clknet_leaf_39_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19370_ (.D(_04948_),
    .Q(\design_top.MEM[24][23] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19371_ (.D(_04949_),
    .Q(\design_top.MEM[9][16] ),
    .CLK(clknet_leaf_278_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19372_ (.D(_04950_),
    .Q(\design_top.MEM[9][17] ),
    .CLK(clknet_leaf_283_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19373_ (.D(_04951_),
    .Q(\design_top.MEM[9][18] ),
    .CLK(clknet_leaf_291_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19374_ (.D(_04952_),
    .Q(\design_top.MEM[9][19] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19375_ (.D(_04953_),
    .Q(\design_top.MEM[9][20] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19376_ (.D(_04954_),
    .Q(\design_top.MEM[9][21] ),
    .CLK(clknet_leaf_277_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19377_ (.D(_04955_),
    .Q(\design_top.MEM[9][22] ),
    .CLK(clknet_leaf_277_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19378_ (.D(_04956_),
    .Q(\design_top.MEM[9][23] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19379_ (.D(_04957_),
    .Q(\design_top.MEM[24][8] ),
    .CLK(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19380_ (.D(_04958_),
    .Q(\design_top.MEM[24][9] ),
    .CLK(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19381_ (.D(_04959_),
    .Q(\design_top.MEM[24][10] ),
    .CLK(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19382_ (.D(_04960_),
    .Q(\design_top.MEM[24][11] ),
    .CLK(clknet_leaf_318_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19383_ (.D(_04961_),
    .Q(\design_top.MEM[24][12] ),
    .CLK(clknet_leaf_318_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19384_ (.D(_04962_),
    .Q(\design_top.MEM[24][13] ),
    .CLK(clknet_leaf_320_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19385_ (.D(_04963_),
    .Q(\design_top.MEM[24][14] ),
    .CLK(clknet_leaf_318_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19386_ (.D(_04964_),
    .Q(\design_top.MEM[24][15] ),
    .CLK(clknet_leaf_319_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19387_ (.D(_04965_),
    .Q(\design_top.MEM[23][24] ),
    .CLK(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19388_ (.D(_04966_),
    .Q(\design_top.MEM[23][25] ),
    .CLK(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19389_ (.D(_04967_),
    .Q(\design_top.MEM[23][26] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19390_ (.D(_04968_),
    .Q(\design_top.MEM[23][27] ),
    .CLK(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19391_ (.D(_04969_),
    .Q(\design_top.MEM[23][28] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19392_ (.D(_04970_),
    .Q(\design_top.MEM[23][29] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19393_ (.D(_04971_),
    .Q(\design_top.MEM[23][30] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19394_ (.D(_04972_),
    .Q(\design_top.MEM[23][31] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19395_ (.D(_04973_),
    .Q(\design_top.MEM[9][8] ),
    .CLK(clknet_leaf_308_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19396_ (.D(_04974_),
    .Q(\design_top.MEM[9][9] ),
    .CLK(clknet_leaf_307_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19397_ (.D(_04975_),
    .Q(\design_top.MEM[9][10] ),
    .CLK(clknet_leaf_287_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19398_ (.D(_04976_),
    .Q(\design_top.MEM[9][11] ),
    .CLK(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19399_ (.D(_04977_),
    .Q(\design_top.MEM[9][12] ),
    .CLK(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19400_ (.D(_04978_),
    .Q(\design_top.MEM[9][13] ),
    .CLK(clknet_leaf_307_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19401_ (.D(_04979_),
    .Q(\design_top.MEM[9][14] ),
    .CLK(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19402_ (.D(_04980_),
    .Q(\design_top.MEM[9][15] ),
    .CLK(clknet_leaf_306_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19403_ (.D(_04981_),
    .Q(\design_top.MEM[23][16] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19404_ (.D(_04982_),
    .Q(\design_top.MEM[23][17] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19405_ (.D(_04983_),
    .Q(\design_top.MEM[23][18] ),
    .CLK(clknet_leaf_287_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19406_ (.D(_04984_),
    .Q(\design_top.MEM[23][19] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19407_ (.D(_04985_),
    .Q(\design_top.MEM[23][20] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19408_ (.D(_04986_),
    .Q(\design_top.MEM[23][21] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19409_ (.D(_04987_),
    .Q(\design_top.MEM[23][22] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19410_ (.D(_04988_),
    .Q(\design_top.MEM[23][23] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19411_ (.D(_04989_),
    .Q(\design_top.MEM[8][24] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19412_ (.D(_04990_),
    .Q(\design_top.MEM[8][25] ),
    .CLK(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19413_ (.D(_04991_),
    .Q(\design_top.MEM[8][26] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19414_ (.D(_04992_),
    .Q(\design_top.MEM[8][27] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19415_ (.D(_04993_),
    .Q(\design_top.MEM[8][28] ),
    .CLK(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19416_ (.D(_04994_),
    .Q(\design_top.MEM[8][29] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19417_ (.D(_04995_),
    .Q(\design_top.MEM[8][30] ),
    .CLK(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19418_ (.D(_04996_),
    .Q(\design_top.MEM[8][31] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19419_ (.D(_04997_),
    .Q(\design_top.MEM[8][16] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19420_ (.D(_04998_),
    .Q(\design_top.MEM[8][17] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19421_ (.D(_04999_),
    .Q(\design_top.MEM[8][18] ),
    .CLK(clknet_leaf_292_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19422_ (.D(_05000_),
    .Q(\design_top.MEM[8][19] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19423_ (.D(_05001_),
    .Q(\design_top.MEM[8][20] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19424_ (.D(_05002_),
    .Q(\design_top.MEM[8][21] ),
    .CLK(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19425_ (.D(_05003_),
    .Q(\design_top.MEM[8][22] ),
    .CLK(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19426_ (.D(_05004_),
    .Q(\design_top.MEM[8][23] ),
    .CLK(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19427_ (.D(_05005_),
    .Q(\design_top.MEM[8][8] ),
    .CLK(clknet_leaf_308_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19428_ (.D(_05006_),
    .Q(\design_top.MEM[8][9] ),
    .CLK(clknet_leaf_308_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19429_ (.D(_05007_),
    .Q(\design_top.MEM[8][10] ),
    .CLK(clknet_leaf_287_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19430_ (.D(_05008_),
    .Q(\design_top.MEM[8][11] ),
    .CLK(clknet_leaf_306_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19431_ (.D(_05009_),
    .Q(\design_top.MEM[8][12] ),
    .CLK(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19432_ (.D(_05010_),
    .Q(\design_top.MEM[8][13] ),
    .CLK(clknet_leaf_306_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19433_ (.D(_05011_),
    .Q(\design_top.MEM[8][14] ),
    .CLK(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19434_ (.D(_05012_),
    .Q(\design_top.MEM[8][15] ),
    .CLK(clknet_leaf_306_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19435_ (.D(_05013_),
    .Q(\design_top.MEM[7][16] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19436_ (.D(_05014_),
    .Q(\design_top.MEM[7][17] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19437_ (.D(_05015_),
    .Q(\design_top.MEM[7][18] ),
    .CLK(clknet_leaf_292_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19438_ (.D(_05016_),
    .Q(\design_top.MEM[7][19] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19439_ (.D(_05017_),
    .Q(\design_top.MEM[7][20] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19440_ (.D(_05018_),
    .Q(\design_top.MEM[7][21] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19441_ (.D(_05019_),
    .Q(\design_top.MEM[7][22] ),
    .CLK(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19442_ (.D(_05020_),
    .Q(\design_top.MEM[7][23] ),
    .CLK(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19443_ (.D(_05021_),
    .Q(\design_top.MEM[22][8] ),
    .CLK(clknet_leaf_312_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19444_ (.D(_05022_),
    .Q(\design_top.MEM[22][9] ),
    .CLK(clknet_leaf_312_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19445_ (.D(_05023_),
    .Q(\design_top.MEM[22][10] ),
    .CLK(clknet_leaf_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19446_ (.D(_05024_),
    .Q(\design_top.MEM[22][11] ),
    .CLK(clknet_leaf_316_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19447_ (.D(_05025_),
    .Q(\design_top.MEM[22][12] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19448_ (.D(_05026_),
    .Q(\design_top.MEM[22][13] ),
    .CLK(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19449_ (.D(_05027_),
    .Q(\design_top.MEM[22][14] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19450_ (.D(_05028_),
    .Q(\design_top.MEM[22][15] ),
    .CLK(clknet_leaf_314_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19451_ (.D(_05029_),
    .Q(\design_top.MEM[21][24] ),
    .CLK(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19452_ (.D(_05030_),
    .Q(\design_top.MEM[21][25] ),
    .CLK(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19453_ (.D(_05031_),
    .Q(\design_top.MEM[21][26] ),
    .CLK(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19454_ (.D(_05032_),
    .Q(\design_top.MEM[21][27] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19455_ (.D(_05033_),
    .Q(\design_top.MEM[21][28] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19456_ (.D(_05034_),
    .Q(\design_top.MEM[21][29] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19457_ (.D(_05035_),
    .Q(\design_top.MEM[21][30] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19458_ (.D(_05036_),
    .Q(\design_top.MEM[21][31] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19459_ (.D(_05037_),
    .Q(\design_top.MEM[21][16] ),
    .CLK(clknet_leaf_284_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19460_ (.D(_05038_),
    .Q(\design_top.MEM[21][17] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19461_ (.D(_05039_),
    .Q(\design_top.MEM[21][18] ),
    .CLK(clknet_leaf_287_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19462_ (.D(_05040_),
    .Q(\design_top.MEM[21][19] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19463_ (.D(_05041_),
    .Q(\design_top.MEM[21][20] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19464_ (.D(_05042_),
    .Q(\design_top.MEM[21][21] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19465_ (.D(_05043_),
    .Q(\design_top.MEM[21][22] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19466_ (.D(_05044_),
    .Q(\design_top.MEM[21][23] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19467_ (.D(_05045_),
    .Q(\design_top.MEM[21][8] ),
    .CLK(clknet_leaf_312_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19468_ (.D(_05046_),
    .Q(\design_top.MEM[21][9] ),
    .CLK(clknet_leaf_312_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19469_ (.D(_05047_),
    .Q(\design_top.MEM[21][10] ),
    .CLK(clknet_leaf_311_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19470_ (.D(_05048_),
    .Q(\design_top.MEM[21][11] ),
    .CLK(clknet_leaf_316_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19471_ (.D(_05049_),
    .Q(\design_top.MEM[21][12] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19472_ (.D(_05050_),
    .Q(\design_top.MEM[21][13] ),
    .CLK(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19473_ (.D(_05051_),
    .Q(\design_top.MEM[21][14] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19474_ (.D(_05052_),
    .Q(\design_top.MEM[21][15] ),
    .CLK(clknet_leaf_314_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19475_ (.D(_05053_),
    .Q(\design_top.MEM[20][24] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19476_ (.D(_05054_),
    .Q(\design_top.MEM[20][25] ),
    .CLK(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19477_ (.D(_05055_),
    .Q(\design_top.MEM[20][26] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19478_ (.D(_05056_),
    .Q(\design_top.MEM[20][27] ),
    .CLK(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19479_ (.D(_05057_),
    .Q(\design_top.MEM[20][28] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19480_ (.D(_05058_),
    .Q(\design_top.MEM[20][29] ),
    .CLK(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19481_ (.D(_05059_),
    .Q(\design_top.MEM[20][30] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19482_ (.D(_05060_),
    .Q(\design_top.MEM[20][31] ),
    .CLK(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19483_ (.D(_05061_),
    .Q(\design_top.MEM[20][16] ),
    .CLK(clknet_leaf_284_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19484_ (.D(_05062_),
    .Q(\design_top.MEM[20][17] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19485_ (.D(_05063_),
    .Q(\design_top.MEM[20][18] ),
    .CLK(clknet_leaf_287_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19486_ (.D(_05064_),
    .Q(\design_top.MEM[20][19] ),
    .CLK(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19487_ (.D(_05065_),
    .Q(\design_top.MEM[20][20] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19488_ (.D(_05066_),
    .Q(\design_top.MEM[20][21] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19489_ (.D(_05067_),
    .Q(\design_top.MEM[20][22] ),
    .CLK(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19490_ (.D(_05068_),
    .Q(\design_top.MEM[20][23] ),
    .CLK(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19491_ (.D(_05069_),
    .Q(\design_top.MEM[20][8] ),
    .CLK(clknet_leaf_311_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19492_ (.D(_05070_),
    .Q(\design_top.MEM[20][9] ),
    .CLK(clknet_leaf_312_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19493_ (.D(_05071_),
    .Q(\design_top.MEM[20][10] ),
    .CLK(clknet_leaf_311_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19494_ (.D(_05072_),
    .Q(\design_top.MEM[20][11] ),
    .CLK(clknet_leaf_316_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19495_ (.D(_05073_),
    .Q(\design_top.MEM[20][12] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19496_ (.D(_05074_),
    .Q(\design_top.MEM[20][13] ),
    .CLK(clknet_leaf_314_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19497_ (.D(_05075_),
    .Q(\design_top.MEM[20][14] ),
    .CLK(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19498_ (.D(_05076_),
    .Q(\design_top.MEM[20][15] ),
    .CLK(clknet_leaf_314_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19499_ (.D(_05077_),
    .Q(\design_top.MEM[7][24] ),
    .CLK(clknet_leaf_31_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19500_ (.D(_05078_),
    .Q(\design_top.MEM[7][25] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19501_ (.D(_05079_),
    .Q(\design_top.MEM[7][26] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19502_ (.D(_05080_),
    .Q(\design_top.MEM[7][27] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19503_ (.D(_05081_),
    .Q(\design_top.MEM[7][28] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19504_ (.D(_05082_),
    .Q(\design_top.MEM[7][29] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19505_ (.D(_05083_),
    .Q(\design_top.MEM[7][30] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19506_ (.D(_05084_),
    .Q(\design_top.MEM[7][31] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19507_ (.D(_05085_),
    .Q(\design_top.MEM[7][8] ),
    .CLK(clknet_leaf_294_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19508_ (.D(_05086_),
    .Q(\design_top.MEM[7][9] ),
    .CLK(clknet_leaf_294_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19509_ (.D(_05087_),
    .Q(\design_top.MEM[7][10] ),
    .CLK(clknet_leaf_290_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19510_ (.D(_05088_),
    .Q(\design_top.MEM[7][11] ),
    .CLK(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19511_ (.D(_05089_),
    .Q(\design_top.MEM[7][12] ),
    .CLK(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19512_ (.D(_05090_),
    .Q(\design_top.MEM[7][13] ),
    .CLK(clknet_leaf_296_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19513_ (.D(_05091_),
    .Q(\design_top.MEM[7][14] ),
    .CLK(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19514_ (.D(_05092_),
    .Q(\design_top.MEM[7][15] ),
    .CLK(clknet_leaf_296_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19515_ (.D(_05093_),
    .Q(\design_top.MEM[6][24] ),
    .CLK(clknet_leaf_31_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19516_ (.D(_05094_),
    .Q(\design_top.MEM[6][25] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19517_ (.D(_05095_),
    .Q(\design_top.MEM[6][26] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19518_ (.D(_05096_),
    .Q(\design_top.MEM[6][27] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19519_ (.D(_05097_),
    .Q(\design_top.MEM[6][28] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19520_ (.D(_05098_),
    .Q(\design_top.MEM[6][29] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19521_ (.D(_05099_),
    .Q(\design_top.MEM[6][30] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19522_ (.D(_05100_),
    .Q(\design_top.MEM[6][31] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19523_ (.D(_05101_),
    .Q(\design_top.MEM[1][24] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19524_ (.D(_05102_),
    .Q(\design_top.MEM[1][25] ),
    .CLK(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19525_ (.D(_05103_),
    .Q(\design_top.MEM[1][26] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19526_ (.D(_05104_),
    .Q(\design_top.MEM[1][27] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19527_ (.D(_05105_),
    .Q(\design_top.MEM[1][28] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19528_ (.D(_05106_),
    .Q(\design_top.MEM[1][29] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19529_ (.D(_05107_),
    .Q(\design_top.MEM[1][30] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19530_ (.D(_05108_),
    .Q(\design_top.MEM[1][31] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19531_ (.D(_05109_),
    .Q(\design_top.MEM[1][16] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19532_ (.D(_05110_),
    .Q(\design_top.MEM[1][17] ),
    .CLK(clknet_leaf_281_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19533_ (.D(_05111_),
    .Q(\design_top.MEM[1][18] ),
    .CLK(clknet_leaf_291_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19534_ (.D(_05112_),
    .Q(\design_top.MEM[1][19] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19535_ (.D(_05113_),
    .Q(\design_top.MEM[1][20] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19536_ (.D(_05114_),
    .Q(\design_top.MEM[1][21] ),
    .CLK(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19537_ (.D(_05115_),
    .Q(\design_top.MEM[1][22] ),
    .CLK(clknet_leaf_277_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19538_ (.D(_05116_),
    .Q(\design_top.MEM[1][23] ),
    .CLK(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19539_ (.D(_05117_),
    .Q(\design_top.MEM[1][8] ),
    .CLK(clknet_leaf_289_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19540_ (.D(_05118_),
    .Q(\design_top.MEM[1][9] ),
    .CLK(clknet_leaf_307_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19541_ (.D(_05119_),
    .Q(\design_top.MEM[1][10] ),
    .CLK(clknet_leaf_288_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19542_ (.D(_05120_),
    .Q(\design_top.MEM[1][11] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19543_ (.D(_05121_),
    .Q(\design_top.MEM[1][12] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19544_ (.D(_05122_),
    .Q(\design_top.MEM[1][13] ),
    .CLK(clknet_leaf_302_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19545_ (.D(_05123_),
    .Q(\design_top.MEM[1][14] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19546_ (.D(_05124_),
    .Q(\design_top.MEM[1][15] ),
    .CLK(clknet_leaf_302_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19547_ (.D(_05125_),
    .Q(\design_top.MEM[19][24] ),
    .CLK(clknet_leaf_29_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19548_ (.D(_05126_),
    .Q(\design_top.MEM[19][25] ),
    .CLK(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19549_ (.D(_05127_),
    .Q(\design_top.MEM[19][26] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19550_ (.D(_05128_),
    .Q(\design_top.MEM[19][27] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19551_ (.D(_05129_),
    .Q(\design_top.MEM[19][28] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19552_ (.D(_05130_),
    .Q(\design_top.MEM[19][29] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19553_ (.D(_05131_),
    .Q(\design_top.MEM[19][30] ),
    .CLK(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19554_ (.D(_05132_),
    .Q(\design_top.MEM[19][31] ),
    .CLK(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19555_ (.D(_05133_),
    .Q(\design_top.MEM[19][16] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19556_ (.D(_05134_),
    .Q(\design_top.MEM[19][17] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19557_ (.D(_05135_),
    .Q(\design_top.MEM[19][18] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19558_ (.D(_05136_),
    .Q(\design_top.MEM[19][19] ),
    .CLK(clknet_leaf_37_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19559_ (.D(_05137_),
    .Q(\design_top.MEM[19][20] ),
    .CLK(clknet_leaf_37_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19560_ (.D(_05138_),
    .Q(\design_top.MEM[19][21] ),
    .CLK(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19561_ (.D(_05139_),
    .Q(\design_top.MEM[19][22] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19562_ (.D(_05140_),
    .Q(\design_top.MEM[19][23] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19563_ (.D(_05141_),
    .Q(\design_top.MEM[19][8] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19564_ (.D(_05142_),
    .Q(\design_top.MEM[19][9] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19565_ (.D(_05143_),
    .Q(\design_top.MEM[19][10] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19566_ (.D(_05144_),
    .Q(\design_top.MEM[19][11] ),
    .CLK(clknet_leaf_321_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19567_ (.D(_05145_),
    .Q(\design_top.MEM[19][12] ),
    .CLK(clknet_leaf_323_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19568_ (.D(_05146_),
    .Q(\design_top.MEM[19][13] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19569_ (.D(_05147_),
    .Q(\design_top.MEM[19][14] ),
    .CLK(clknet_leaf_321_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19570_ (.D(_05148_),
    .Q(\design_top.MEM[19][15] ),
    .CLK(clknet_leaf_323_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19571_ (.D(_05149_),
    .Q(\design_top.MEM[18][24] ),
    .CLK(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19572_ (.D(_05150_),
    .Q(\design_top.MEM[18][25] ),
    .CLK(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19573_ (.D(_05151_),
    .Q(\design_top.MEM[18][26] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19574_ (.D(_05152_),
    .Q(\design_top.MEM[18][27] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19575_ (.D(_05153_),
    .Q(\design_top.MEM[18][28] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19576_ (.D(_05154_),
    .Q(\design_top.MEM[18][29] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19577_ (.D(_05155_),
    .Q(\design_top.MEM[18][30] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19578_ (.D(_05156_),
    .Q(\design_top.MEM[18][31] ),
    .CLK(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19579_ (.D(_05157_),
    .Q(\design_top.MEM[18][16] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19580_ (.D(_05158_),
    .Q(\design_top.MEM[18][17] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19581_ (.D(_05159_),
    .Q(\design_top.MEM[18][18] ),
    .CLK(clknet_leaf_31_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19582_ (.D(_05160_),
    .Q(\design_top.MEM[18][19] ),
    .CLK(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19583_ (.D(_05161_),
    .Q(\design_top.MEM[18][20] ),
    .CLK(clknet_leaf_48_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19584_ (.D(_05162_),
    .Q(\design_top.MEM[18][21] ),
    .CLK(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19585_ (.D(_05163_),
    .Q(\design_top.MEM[18][22] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19586_ (.D(_05164_),
    .Q(\design_top.MEM[18][23] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19587_ (.D(_05165_),
    .Q(\design_top.MEM[18][8] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19588_ (.D(_05166_),
    .Q(\design_top.MEM[18][9] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19589_ (.D(_05167_),
    .Q(\design_top.MEM[18][10] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19590_ (.D(_05168_),
    .Q(\design_top.MEM[18][11] ),
    .CLK(clknet_leaf_321_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19591_ (.D(_05169_),
    .Q(\design_top.MEM[18][12] ),
    .CLK(clknet_leaf_323_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19592_ (.D(_05170_),
    .Q(\design_top.MEM[18][13] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19593_ (.D(_05171_),
    .Q(\design_top.MEM[18][14] ),
    .CLK(clknet_leaf_321_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19594_ (.D(_05172_),
    .Q(\design_top.MEM[18][15] ),
    .CLK(clknet_leaf_323_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19595_ (.D(_05173_),
    .Q(\design_top.MEM[17][24] ),
    .CLK(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19596_ (.D(_05174_),
    .Q(\design_top.MEM[17][25] ),
    .CLK(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19597_ (.D(_05175_),
    .Q(\design_top.MEM[17][26] ),
    .CLK(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19598_ (.D(_05176_),
    .Q(\design_top.MEM[17][27] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19599_ (.D(_05177_),
    .Q(\design_top.MEM[17][28] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19600_ (.D(_05178_),
    .Q(\design_top.MEM[17][29] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19601_ (.D(_05179_),
    .Q(\design_top.MEM[17][30] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19602_ (.D(_05180_),
    .Q(\design_top.MEM[17][31] ),
    .CLK(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19603_ (.D(_05181_),
    .Q(\design_top.MEM[17][16] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19604_ (.D(_05182_),
    .Q(\design_top.MEM[17][17] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19605_ (.D(_05183_),
    .Q(\design_top.MEM[17][18] ),
    .CLK(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19606_ (.D(_05184_),
    .Q(\design_top.MEM[17][19] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19607_ (.D(_05185_),
    .Q(\design_top.MEM[17][20] ),
    .CLK(clknet_leaf_48_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19608_ (.D(_05186_),
    .Q(\design_top.MEM[17][21] ),
    .CLK(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19609_ (.D(_05187_),
    .Q(\design_top.MEM[17][22] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19610_ (.D(_05188_),
    .Q(\design_top.MEM[17][23] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19611_ (.D(_05189_),
    .Q(\design_top.MEM[17][8] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19612_ (.D(_05190_),
    .Q(\design_top.MEM[17][9] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19613_ (.D(_05191_),
    .Q(\design_top.MEM[17][10] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19614_ (.D(_05192_),
    .Q(\design_top.MEM[17][11] ),
    .CLK(clknet_leaf_320_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19615_ (.D(_05193_),
    .Q(\design_top.MEM[17][12] ),
    .CLK(clknet_leaf_322_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19616_ (.D(_05194_),
    .Q(\design_top.MEM[17][13] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19617_ (.D(_05195_),
    .Q(\design_top.MEM[17][14] ),
    .CLK(clknet_leaf_322_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19618_ (.D(_05196_),
    .Q(\design_top.MEM[17][15] ),
    .CLK(clknet_leaf_323_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19619_ (.D(_05197_),
    .Q(\design_top.MEM[16][16] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19620_ (.D(_05198_),
    .Q(\design_top.MEM[16][17] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19621_ (.D(_05199_),
    .Q(\design_top.MEM[16][18] ),
    .CLK(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19622_ (.D(_05200_),
    .Q(\design_top.MEM[16][19] ),
    .CLK(clknet_leaf_37_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19623_ (.D(_05201_),
    .Q(\design_top.MEM[16][20] ),
    .CLK(clknet_leaf_37_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19624_ (.D(_05202_),
    .Q(\design_top.MEM[16][21] ),
    .CLK(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19625_ (.D(_05203_),
    .Q(\design_top.MEM[16][22] ),
    .CLK(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19626_ (.D(_05204_),
    .Q(\design_top.MEM[16][23] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19627_ (.D(_05205_),
    .Q(\design_top.MEM[16][24] ),
    .CLK(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19628_ (.D(_05206_),
    .Q(\design_top.MEM[16][25] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19629_ (.D(_05207_),
    .Q(\design_top.MEM[16][26] ),
    .CLK(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19630_ (.D(_05208_),
    .Q(\design_top.MEM[16][27] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19631_ (.D(_05209_),
    .Q(\design_top.MEM[16][28] ),
    .CLK(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19632_ (.D(_05210_),
    .Q(\design_top.MEM[16][29] ),
    .CLK(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19633_ (.D(_05211_),
    .Q(\design_top.MEM[16][30] ),
    .CLK(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19634_ (.D(_05212_),
    .Q(\design_top.MEM[16][31] ),
    .CLK(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19635_ (.D(_05213_),
    .Q(\design_top.MEM[16][8] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19636_ (.D(_05214_),
    .Q(\design_top.MEM[16][9] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19637_ (.D(_05215_),
    .Q(\design_top.MEM[16][10] ),
    .CLK(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19638_ (.D(_05216_),
    .Q(\design_top.MEM[16][11] ),
    .CLK(clknet_leaf_321_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19639_ (.D(_05217_),
    .Q(\design_top.MEM[16][12] ),
    .CLK(clknet_leaf_323_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19640_ (.D(_05218_),
    .Q(\design_top.MEM[16][13] ),
    .CLK(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19641_ (.D(_05219_),
    .Q(\design_top.MEM[16][14] ),
    .CLK(clknet_leaf_322_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19642_ (.D(_05220_),
    .Q(\design_top.MEM[16][15] ),
    .CLK(clknet_leaf_323_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19643_ (.D(_05221_),
    .Q(\design_top.MEM[15][24] ),
    .CLK(clknet_leaf_29_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19644_ (.D(_05222_),
    .Q(\design_top.MEM[15][25] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19645_ (.D(_05223_),
    .Q(\design_top.MEM[15][26] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19646_ (.D(_05224_),
    .Q(\design_top.MEM[15][27] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19647_ (.D(_05225_),
    .Q(\design_top.MEM[15][28] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19648_ (.D(_05226_),
    .Q(\design_top.MEM[15][29] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19649_ (.D(_05227_),
    .Q(\design_top.MEM[15][30] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19650_ (.D(_05228_),
    .Q(\design_top.MEM[15][31] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19651_ (.D(_05229_),
    .Q(\design_top.MEM[15][16] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19652_ (.D(_05230_),
    .Q(\design_top.MEM[15][17] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19653_ (.D(_05231_),
    .Q(\design_top.MEM[15][18] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19654_ (.D(_05232_),
    .Q(\design_top.MEM[15][19] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19655_ (.D(_05233_),
    .Q(\design_top.MEM[15][20] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19656_ (.D(_05234_),
    .Q(\design_top.MEM[15][21] ),
    .CLK(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19657_ (.D(_05235_),
    .Q(\design_top.MEM[15][22] ),
    .CLK(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19658_ (.D(_05236_),
    .Q(\design_top.MEM[15][23] ),
    .CLK(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19659_ (.D(_05237_),
    .Q(\design_top.MEM[15][8] ),
    .CLK(clknet_leaf_289_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19660_ (.D(_05238_),
    .Q(\design_top.MEM[15][9] ),
    .CLK(clknet_leaf_307_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19661_ (.D(_05239_),
    .Q(\design_top.MEM[15][10] ),
    .CLK(clknet_leaf_288_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19662_ (.D(_05240_),
    .Q(\design_top.MEM[15][11] ),
    .CLK(clknet_leaf_302_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19663_ (.D(_05241_),
    .Q(\design_top.MEM[15][12] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19664_ (.D(_05242_),
    .Q(\design_top.MEM[15][13] ),
    .CLK(clknet_leaf_307_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19665_ (.D(_05243_),
    .Q(\design_top.MEM[15][14] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19666_ (.D(_05244_),
    .Q(\design_top.MEM[15][15] ),
    .CLK(clknet_leaf_302_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19667_ (.D(_05245_),
    .Q(\design_top.MEM[14][24] ),
    .CLK(clknet_leaf_29_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19668_ (.D(_05246_),
    .Q(\design_top.MEM[14][25] ),
    .CLK(clknet_leaf_29_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19669_ (.D(_05247_),
    .Q(\design_top.MEM[14][26] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19670_ (.D(_05248_),
    .Q(\design_top.MEM[14][27] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19671_ (.D(_05249_),
    .Q(\design_top.MEM[14][28] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19672_ (.D(_05250_),
    .Q(\design_top.MEM[14][29] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19673_ (.D(_05251_),
    .Q(\design_top.MEM[14][30] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19674_ (.D(_05252_),
    .Q(\design_top.MEM[14][31] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19675_ (.D(_05253_),
    .Q(\design_top.MEM[14][16] ),
    .CLK(clknet_leaf_268_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19676_ (.D(_05254_),
    .Q(\design_top.MEM[14][17] ),
    .CLK(clknet_leaf_267_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19677_ (.D(_05255_),
    .Q(\design_top.MEM[14][18] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19678_ (.D(_05256_),
    .Q(\design_top.MEM[14][19] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19679_ (.D(_05257_),
    .Q(\design_top.MEM[14][20] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19680_ (.D(_05258_),
    .Q(\design_top.MEM[14][21] ),
    .CLK(clknet_leaf_269_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19681_ (.D(_05259_),
    .Q(\design_top.MEM[14][22] ),
    .CLK(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19682_ (.D(_05260_),
    .Q(\design_top.MEM[14][23] ),
    .CLK(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19683_ (.D(_05261_),
    .Q(\design_top.MEM[14][8] ),
    .CLK(clknet_leaf_289_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19684_ (.D(_05262_),
    .Q(\design_top.MEM[14][9] ),
    .CLK(clknet_leaf_294_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19685_ (.D(_05263_),
    .Q(\design_top.MEM[14][10] ),
    .CLK(clknet_leaf_290_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19686_ (.D(_05264_),
    .Q(\design_top.MEM[14][11] ),
    .CLK(clknet_leaf_300_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19687_ (.D(_05265_),
    .Q(\design_top.MEM[14][12] ),
    .CLK(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19688_ (.D(_05266_),
    .Q(\design_top.MEM[14][13] ),
    .CLK(clknet_leaf_295_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19689_ (.D(_05267_),
    .Q(\design_top.MEM[14][14] ),
    .CLK(clknet_leaf_301_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19690_ (.D(_05268_),
    .Q(\design_top.MEM[14][15] ),
    .CLK(clknet_leaf_301_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19691_ (.D(_05269_),
    .Q(\design_top.MEM[13][24] ),
    .CLK(clknet_leaf_31_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19692_ (.D(_05270_),
    .Q(\design_top.MEM[13][25] ),
    .CLK(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19693_ (.D(_05271_),
    .Q(\design_top.MEM[13][26] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19694_ (.D(_05272_),
    .Q(\design_top.MEM[13][27] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19695_ (.D(_05273_),
    .Q(\design_top.MEM[13][28] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19696_ (.D(_05274_),
    .Q(\design_top.MEM[13][29] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19697_ (.D(_05275_),
    .Q(\design_top.MEM[13][30] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19698_ (.D(_05276_),
    .Q(\design_top.MEM[13][31] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19699_ (.D(_05277_),
    .Q(\design_top.MEM[13][16] ),
    .CLK(clknet_leaf_268_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19700_ (.D(_05278_),
    .Q(\design_top.MEM[13][17] ),
    .CLK(clknet_leaf_267_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19701_ (.D(_05279_),
    .Q(\design_top.MEM[13][18] ),
    .CLK(clknet_leaf_267_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19702_ (.D(_05280_),
    .Q(\design_top.MEM[13][19] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19703_ (.D(_05281_),
    .Q(\design_top.MEM[13][20] ),
    .CLK(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19704_ (.D(_05282_),
    .Q(\design_top.MEM[13][21] ),
    .CLK(clknet_leaf_269_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19705_ (.D(_05283_),
    .Q(\design_top.MEM[13][22] ),
    .CLK(clknet_leaf_272_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19706_ (.D(_05284_),
    .Q(\design_top.MEM[13][23] ),
    .CLK(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19707_ (.D(_05285_),
    .Q(\design_top.MEM[6][16] ),
    .CLK(clknet_leaf_270_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19708_ (.D(_05286_),
    .Q(\design_top.MEM[6][17] ),
    .CLK(clknet_leaf_267_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19709_ (.D(_05287_),
    .Q(\design_top.MEM[6][18] ),
    .CLK(clknet_leaf_254_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19710_ (.D(_05288_),
    .Q(\design_top.MEM[6][19] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19711_ (.D(_05289_),
    .Q(\design_top.MEM[6][20] ),
    .CLK(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19712_ (.D(_05290_),
    .Q(\design_top.MEM[6][21] ),
    .CLK(clknet_leaf_269_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19713_ (.D(_05291_),
    .Q(\design_top.MEM[6][22] ),
    .CLK(clknet_leaf_271_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19714_ (.D(_05292_),
    .Q(\design_top.MEM[6][23] ),
    .CLK(clknet_leaf_272_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19715_ (.D(_05293_),
    .Q(\design_top.MEM[6][8] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19716_ (.D(_05294_),
    .Q(\design_top.MEM[6][9] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19717_ (.D(_05295_),
    .Q(\design_top.MEM[6][10] ),
    .CLK(clknet_leaf_292_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19718_ (.D(_05296_),
    .Q(\design_top.MEM[6][11] ),
    .CLK(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19719_ (.D(_05297_),
    .Q(\design_top.MEM[6][12] ),
    .CLK(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19720_ (.D(_05298_),
    .Q(\design_top.MEM[6][13] ),
    .CLK(clknet_leaf_296_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19721_ (.D(_05299_),
    .Q(\design_top.MEM[6][14] ),
    .CLK(clknet_leaf_298_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19722_ (.D(_05300_),
    .Q(\design_top.MEM[6][15] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19723_ (.D(_05301_),
    .Q(\design_top.MEM[5][24] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19724_ (.D(_05302_),
    .Q(\design_top.MEM[5][25] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19725_ (.D(_05303_),
    .Q(\design_top.MEM[5][26] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19726_ (.D(_05304_),
    .Q(\design_top.MEM[5][27] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19727_ (.D(_05305_),
    .Q(\design_top.MEM[5][28] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19728_ (.D(_05306_),
    .Q(\design_top.MEM[5][29] ),
    .CLK(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19729_ (.D(_05307_),
    .Q(\design_top.MEM[5][30] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19730_ (.D(_05308_),
    .Q(\design_top.MEM[5][31] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19731_ (.D(_05309_),
    .Q(\design_top.MEM[5][16] ),
    .CLK(clknet_leaf_268_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19732_ (.D(_05310_),
    .Q(\design_top.MEM[5][17] ),
    .CLK(clknet_leaf_267_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19733_ (.D(_05311_),
    .Q(\design_top.MEM[5][18] ),
    .CLK(clknet_leaf_267_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19734_ (.D(_05312_),
    .Q(\design_top.MEM[5][19] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19735_ (.D(_05313_),
    .Q(\design_top.MEM[5][20] ),
    .CLK(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19736_ (.D(_05314_),
    .Q(\design_top.MEM[5][21] ),
    .CLK(clknet_leaf_270_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19737_ (.D(_05315_),
    .Q(\design_top.MEM[5][22] ),
    .CLK(clknet_leaf_272_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19738_ (.D(_05316_),
    .Q(\design_top.MEM[5][23] ),
    .CLK(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19739_ (.D(_05317_),
    .Q(\design_top.MEM[5][8] ),
    .CLK(clknet_leaf_294_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19740_ (.D(_05318_),
    .Q(\design_top.MEM[5][9] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19741_ (.D(_05319_),
    .Q(\design_top.MEM[5][10] ),
    .CLK(clknet_leaf_292_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19742_ (.D(_05320_),
    .Q(\design_top.MEM[5][11] ),
    .CLK(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19743_ (.D(_05321_),
    .Q(\design_top.MEM[5][12] ),
    .CLK(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19744_ (.D(_05322_),
    .Q(\design_top.MEM[5][13] ),
    .CLK(clknet_leaf_296_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19745_ (.D(_05323_),
    .Q(\design_top.MEM[5][14] ),
    .CLK(clknet_leaf_298_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19746_ (.D(_05324_),
    .Q(\design_top.MEM[5][15] ),
    .CLK(clknet_leaf_298_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19747_ (.D(_05325_),
    .Q(\design_top.MEM[4][24] ),
    .CLK(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19748_ (.D(_05326_),
    .Q(\design_top.MEM[4][25] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19749_ (.D(_05327_),
    .Q(\design_top.MEM[4][26] ),
    .CLK(clknet_leaf_37_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19750_ (.D(_05328_),
    .Q(\design_top.MEM[4][27] ),
    .CLK(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19751_ (.D(_05329_),
    .Q(\design_top.MEM[4][28] ),
    .CLK(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19752_ (.D(_05330_),
    .Q(\design_top.MEM[4][29] ),
    .CLK(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19753_ (.D(_05331_),
    .Q(\design_top.MEM[4][30] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19754_ (.D(_05332_),
    .Q(\design_top.MEM[4][31] ),
    .CLK(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19755_ (.D(_05333_),
    .Q(\design_top.MEM[4][16] ),
    .CLK(clknet_leaf_268_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19756_ (.D(_05334_),
    .Q(\design_top.MEM[4][17] ),
    .CLK(clknet_leaf_267_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19757_ (.D(_05335_),
    .Q(\design_top.MEM[4][18] ),
    .CLK(clknet_leaf_254_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19758_ (.D(_05336_),
    .Q(\design_top.MEM[4][19] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19759_ (.D(_05337_),
    .Q(\design_top.MEM[4][20] ),
    .CLK(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19760_ (.D(_05338_),
    .Q(\design_top.MEM[4][21] ),
    .CLK(clknet_leaf_270_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19761_ (.D(_05339_),
    .Q(\design_top.MEM[4][22] ),
    .CLK(clknet_leaf_272_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19762_ (.D(_05340_),
    .Q(\design_top.MEM[4][23] ),
    .CLK(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19763_ (.D(_05341_),
    .Q(\design_top.MEM[4][8] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19764_ (.D(_05342_),
    .Q(\design_top.MEM[4][9] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19765_ (.D(_05343_),
    .Q(\design_top.MEM[4][10] ),
    .CLK(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19766_ (.D(_05344_),
    .Q(\design_top.MEM[4][11] ),
    .CLK(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19767_ (.D(_05345_),
    .Q(\design_top.MEM[4][12] ),
    .CLK(clknet_leaf_298_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19768_ (.D(_05346_),
    .Q(\design_top.MEM[4][13] ),
    .CLK(clknet_leaf_296_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19769_ (.D(_05347_),
    .Q(\design_top.MEM[4][14] ),
    .CLK(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19770_ (.D(_05348_),
    .Q(\design_top.MEM[4][15] ),
    .CLK(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19771_ (.D(_05349_),
    .Q(\design_top.MEM[3][24] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19772_ (.D(_05350_),
    .Q(\design_top.MEM[3][25] ),
    .CLK(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19773_ (.D(_05351_),
    .Q(\design_top.MEM[3][26] ),
    .CLK(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19774_ (.D(_05352_),
    .Q(\design_top.MEM[3][27] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19775_ (.D(_05353_),
    .Q(\design_top.MEM[3][28] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19776_ (.D(_05354_),
    .Q(\design_top.MEM[3][29] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19777_ (.D(_05355_),
    .Q(\design_top.MEM[3][30] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19778_ (.D(_05356_),
    .Q(\design_top.MEM[3][31] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19779_ (.D(_05357_),
    .Q(\design_top.MEM[3][16] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19780_ (.D(_05358_),
    .Q(\design_top.MEM[3][17] ),
    .CLK(clknet_leaf_281_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19781_ (.D(_05359_),
    .Q(\design_top.MEM[3][18] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19782_ (.D(_05360_),
    .Q(\design_top.MEM[3][19] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19783_ (.D(_05361_),
    .Q(\design_top.MEM[3][20] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19784_ (.D(_05362_),
    .Q(\design_top.MEM[3][21] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19785_ (.D(_05363_),
    .Q(\design_top.MEM[3][22] ),
    .CLK(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19786_ (.D(_05364_),
    .Q(\design_top.MEM[3][23] ),
    .CLK(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19787_ (.D(_05365_),
    .Q(\design_top.MEM[3][8] ),
    .CLK(clknet_leaf_289_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19788_ (.D(_05366_),
    .Q(\design_top.MEM[3][9] ),
    .CLK(clknet_leaf_289_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19789_ (.D(_05367_),
    .Q(\design_top.MEM[3][10] ),
    .CLK(clknet_leaf_290_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19790_ (.D(_05368_),
    .Q(\design_top.MEM[3][11] ),
    .CLK(clknet_leaf_300_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19791_ (.D(_05369_),
    .Q(\design_top.MEM[3][12] ),
    .CLK(clknet_leaf_300_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19792_ (.D(_05370_),
    .Q(\design_top.MEM[3][13] ),
    .CLK(clknet_leaf_302_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19793_ (.D(_05371_),
    .Q(\design_top.MEM[3][14] ),
    .CLK(clknet_leaf_300_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19794_ (.D(_05372_),
    .Q(\design_top.MEM[3][15] ),
    .CLK(clknet_leaf_301_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19795_ (.D(_05373_),
    .Q(\design_top.MEM[31][24] ),
    .CLK(clknet_leaf_286_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19796_ (.D(_05374_),
    .Q(\design_top.MEM[31][25] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19797_ (.D(_05375_),
    .Q(\design_top.MEM[31][26] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19798_ (.D(_05376_),
    .Q(\design_top.MEM[31][27] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19799_ (.D(_05377_),
    .Q(\design_top.MEM[31][28] ),
    .CLK(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19800_ (.D(_05378_),
    .Q(\design_top.MEM[31][29] ),
    .CLK(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19801_ (.D(_05379_),
    .Q(\design_top.MEM[31][30] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19802_ (.D(_05380_),
    .Q(\design_top.MEM[31][31] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19803_ (.D(_05381_),
    .Q(\design_top.MEM[31][16] ),
    .CLK(clknet_leaf_283_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19804_ (.D(_05382_),
    .Q(\design_top.MEM[31][17] ),
    .CLK(clknet_leaf_281_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19805_ (.D(_05383_),
    .Q(\design_top.MEM[31][18] ),
    .CLK(clknet_leaf_281_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19806_ (.D(_05384_),
    .Q(\design_top.MEM[31][19] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19807_ (.D(_05385_),
    .Q(\design_top.MEM[31][20] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19808_ (.D(_05386_),
    .Q(\design_top.MEM[31][21] ),
    .CLK(clknet_leaf_278_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19809_ (.D(_05387_),
    .Q(\design_top.MEM[31][22] ),
    .CLK(clknet_leaf_277_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19810_ (.D(_05388_),
    .Q(\design_top.MEM[31][23] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19811_ (.D(_05389_),
    .Q(\design_top.MEM[31][8] ),
    .CLK(clknet_leaf_309_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19812_ (.D(_05390_),
    .Q(\design_top.MEM[31][9] ),
    .CLK(clknet_leaf_308_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19813_ (.D(_05391_),
    .Q(\design_top.MEM[31][10] ),
    .CLK(clknet_leaf_310_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19814_ (.D(_05392_),
    .Q(\design_top.MEM[31][11] ),
    .CLK(clknet_leaf_305_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19815_ (.D(_05393_),
    .Q(\design_top.MEM[31][12] ),
    .CLK(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19816_ (.D(_05394_),
    .Q(\design_top.MEM[31][13] ),
    .CLK(clknet_leaf_306_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19817_ (.D(_05395_),
    .Q(\design_top.MEM[31][14] ),
    .CLK(clknet_leaf_305_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19818_ (.D(_05396_),
    .Q(\design_top.MEM[31][15] ),
    .CLK(clknet_leaf_306_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19819_ (.D(_05397_),
    .Q(\design_top.MEM[30][24] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19820_ (.D(_05398_),
    .Q(\design_top.MEM[30][25] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19821_ (.D(_05399_),
    .Q(\design_top.MEM[30][26] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19822_ (.D(_05400_),
    .Q(\design_top.MEM[30][27] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19823_ (.D(_05401_),
    .Q(\design_top.MEM[30][28] ),
    .CLK(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19824_ (.D(_05402_),
    .Q(\design_top.MEM[30][29] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19825_ (.D(_05403_),
    .Q(\design_top.MEM[30][30] ),
    .CLK(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19826_ (.D(_05404_),
    .Q(\design_top.MEM[30][31] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19827_ (.D(_05405_),
    .Q(\design_top.MEM[30][16] ),
    .CLK(clknet_leaf_278_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19828_ (.D(_05406_),
    .Q(\design_top.MEM[30][17] ),
    .CLK(clknet_leaf_281_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19829_ (.D(_05407_),
    .Q(\design_top.MEM[30][18] ),
    .CLK(clknet_leaf_281_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19830_ (.D(_05408_),
    .Q(\design_top.MEM[30][19] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19831_ (.D(_05409_),
    .Q(\design_top.MEM[30][20] ),
    .CLK(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19832_ (.D(_05410_),
    .Q(\design_top.MEM[30][21] ),
    .CLK(clknet_leaf_277_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19833_ (.D(_05411_),
    .Q(\design_top.MEM[30][22] ),
    .CLK(clknet_leaf_277_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19834_ (.D(_05412_),
    .Q(\design_top.MEM[30][23] ),
    .CLK(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19835_ (.D(_05413_),
    .Q(\design_top.MEM[30][8] ),
    .CLK(clknet_leaf_309_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19836_ (.D(_05414_),
    .Q(\design_top.MEM[30][9] ),
    .CLK(clknet_leaf_308_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19837_ (.D(_05415_),
    .Q(\design_top.MEM[30][10] ),
    .CLK(clknet_leaf_310_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19838_ (.D(_05416_),
    .Q(\design_top.MEM[30][11] ),
    .CLK(clknet_leaf_306_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19839_ (.D(_05417_),
    .Q(\design_top.MEM[30][12] ),
    .CLK(clknet_leaf_305_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19840_ (.D(_05418_),
    .Q(\design_top.MEM[30][13] ),
    .CLK(clknet_leaf_306_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19841_ (.D(_05419_),
    .Q(\design_top.MEM[30][14] ),
    .CLK(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19842_ (.D(_05420_),
    .Q(\design_top.MEM[30][15] ),
    .CLK(clknet_leaf_306_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19843_ (.D(_05421_),
    .Q(\design_top.MEM[2][24] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19844_ (.D(_05422_),
    .Q(\design_top.MEM[2][25] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19845_ (.D(_05423_),
    .Q(\design_top.MEM[2][26] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19846_ (.D(_05424_),
    .Q(\design_top.MEM[2][27] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19847_ (.D(_05425_),
    .Q(\design_top.MEM[2][28] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19848_ (.D(_05426_),
    .Q(\design_top.MEM[2][29] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19849_ (.D(_05427_),
    .Q(\design_top.MEM[2][30] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19850_ (.D(_05428_),
    .Q(\design_top.MEM[2][31] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19851_ (.D(_05429_),
    .Q(\design_top.MEM[11][8] ),
    .CLK(clknet_leaf_308_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19852_ (.D(_05430_),
    .Q(\design_top.MEM[11][9] ),
    .CLK(clknet_leaf_308_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19853_ (.D(_05431_),
    .Q(\design_top.MEM[11][10] ),
    .CLK(clknet_leaf_286_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19854_ (.D(_05432_),
    .Q(\design_top.MEM[11][11] ),
    .CLK(clknet_leaf_305_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19855_ (.D(_05433_),
    .Q(\design_top.MEM[11][12] ),
    .CLK(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19856_ (.D(_05434_),
    .Q(\design_top.MEM[11][13] ),
    .CLK(clknet_leaf_306_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19857_ (.D(_05435_),
    .Q(\design_top.MEM[11][14] ),
    .CLK(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19858_ (.D(_05436_),
    .Q(\design_top.MEM[11][15] ),
    .CLK(clknet_leaf_306_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19859_ (.D(_05437_),
    .Q(\design_top.MEM[10][24] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19860_ (.D(_05438_),
    .Q(\design_top.MEM[10][25] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19861_ (.D(_05439_),
    .Q(\design_top.MEM[10][26] ),
    .CLK(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19862_ (.D(_05440_),
    .Q(\design_top.MEM[10][27] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19863_ (.D(_05441_),
    .Q(\design_top.MEM[10][28] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19864_ (.D(_05442_),
    .Q(\design_top.MEM[10][29] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19865_ (.D(_05443_),
    .Q(\design_top.MEM[10][30] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19866_ (.D(_05444_),
    .Q(\design_top.MEM[10][31] ),
    .CLK(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19867_ (.D(_05445_),
    .Q(\design_top.MEM[10][16] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19868_ (.D(_05446_),
    .Q(\design_top.MEM[10][17] ),
    .CLK(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19869_ (.D(_05447_),
    .Q(\design_top.MEM[10][18] ),
    .CLK(clknet_leaf_292_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19870_ (.D(_05448_),
    .Q(\design_top.MEM[10][19] ),
    .CLK(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19871_ (.D(_05449_),
    .Q(\design_top.MEM[10][20] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19872_ (.D(_05450_),
    .Q(\design_top.MEM[10][21] ),
    .CLK(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19873_ (.D(_05451_),
    .Q(\design_top.MEM[10][22] ),
    .CLK(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19874_ (.D(_05452_),
    .Q(\design_top.MEM[10][23] ),
    .CLK(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19875_ (.D(_05453_),
    .Q(\design_top.IREQ[7] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19876_ (.D(_05454_),
    .Q(\design_top.IACK[7] ),
    .CLK(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19877_ (.D(_05455_),
    .Q(\design_top.MEM[10][8] ),
    .CLK(clknet_leaf_308_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19878_ (.D(_05456_),
    .Q(\design_top.MEM[10][9] ),
    .CLK(clknet_leaf_308_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19879_ (.D(_05457_),
    .Q(\design_top.MEM[10][10] ),
    .CLK(clknet_leaf_286_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19880_ (.D(_05458_),
    .Q(\design_top.MEM[10][11] ),
    .CLK(clknet_leaf_305_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19881_ (.D(_05459_),
    .Q(\design_top.MEM[10][12] ),
    .CLK(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19882_ (.D(_05460_),
    .Q(\design_top.MEM[10][13] ),
    .CLK(clknet_leaf_306_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19883_ (.D(_05461_),
    .Q(\design_top.MEM[10][14] ),
    .CLK(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19884_ (.D(_05462_),
    .Q(\design_top.MEM[10][15] ),
    .CLK(clknet_leaf_306_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19885_ (.D(_05463_),
    .Q(\design_top.MEM[0][16] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19886_ (.D(_05464_),
    .Q(\design_top.MEM[0][17] ),
    .CLK(clknet_leaf_281_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19887_ (.D(_05465_),
    .Q(\design_top.MEM[0][18] ),
    .CLK(clknet_leaf_292_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19888_ (.D(_05466_),
    .Q(\design_top.MEM[0][19] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19889_ (.D(_05467_),
    .Q(\design_top.MEM[0][20] ),
    .CLK(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19890_ (.D(_05468_),
    .Q(\design_top.MEM[0][21] ),
    .CLK(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19891_ (.D(_05469_),
    .Q(\design_top.MEM[0][22] ),
    .CLK(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19892_ (.D(_05470_),
    .Q(\design_top.MEM[0][23] ),
    .CLK(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19893_ (.D(_05471_),
    .Q(\design_top.MEM[0][8] ),
    .CLK(clknet_leaf_289_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19894_ (.D(_05472_),
    .Q(\design_top.MEM[0][9] ),
    .CLK(clknet_leaf_307_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19895_ (.D(_05473_),
    .Q(\design_top.MEM[0][10] ),
    .CLK(clknet_leaf_288_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19896_ (.D(_05474_),
    .Q(\design_top.MEM[0][11] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19897_ (.D(_05475_),
    .Q(\design_top.MEM[0][12] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19898_ (.D(_05476_),
    .Q(\design_top.MEM[0][13] ),
    .CLK(clknet_leaf_307_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19899_ (.D(_05477_),
    .Q(\design_top.MEM[0][14] ),
    .CLK(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19900_ (.D(_05478_),
    .Q(\design_top.MEM[0][15] ),
    .CLK(clknet_leaf_302_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19901_ (.D(_05479_),
    .Q(\design_top.MEM[0][24] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19902_ (.D(_05480_),
    .Q(\design_top.MEM[0][25] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19903_ (.D(_05481_),
    .Q(\design_top.MEM[0][26] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19904_ (.D(_05482_),
    .Q(\design_top.MEM[0][27] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19905_ (.D(_05483_),
    .Q(\design_top.MEM[0][28] ),
    .CLK(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19906_ (.D(_05484_),
    .Q(\design_top.MEM[0][29] ),
    .CLK(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19907_ (.D(_05485_),
    .Q(\design_top.MEM[0][30] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19908_ (.D(_05486_),
    .Q(\design_top.MEM[0][31] ),
    .CLK(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19909_ (.D(_05487_),
    .Q(\design_top.MEM[9][24] ),
    .CLK(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19910_ (.D(_05488_),
    .Q(\design_top.MEM[9][25] ),
    .CLK(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19911_ (.D(_05489_),
    .Q(\design_top.MEM[9][26] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19912_ (.D(_05490_),
    .Q(\design_top.MEM[9][27] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19913_ (.D(_05491_),
    .Q(\design_top.MEM[9][28] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19914_ (.D(_05492_),
    .Q(\design_top.MEM[9][29] ),
    .CLK(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19915_ (.D(_05493_),
    .Q(\design_top.MEM[9][30] ),
    .CLK(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__dfxtp_2 _19916_ (.D(_05494_),
    .Q(\design_top.MEM[9][31] ),
    .CLK(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_user_clock2 (.A(clknet_opt_0_user_clock2),
    .X(clknet_leaf_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_9_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_10_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_11_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_12_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_13_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_14_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_15_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_16_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_17_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_18_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_19_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_20_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_21_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_22_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_23_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_24_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_25_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_26_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_27_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_28_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_user_clock2 (.A(clknet_5_5_0_user_clock2),
    .X(clknet_leaf_29_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_user_clock2 (.A(clknet_5_4_0_user_clock2),
    .X(clknet_leaf_30_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_31_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_32_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_33_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_34_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_35_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_36_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_37_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_38_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_39_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_40_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_41_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_42_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_43_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_44_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_45_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_46_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_47_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_48_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_49_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_user_clock2 (.A(clknet_5_18_0_user_clock2),
    .X(clknet_leaf_50_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_51_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_52_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_53_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_54_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_55_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_56_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_user_clock2 (.A(clknet_opt_2_user_clock2),
    .X(clknet_leaf_57_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_58_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_59_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_60_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_61_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_62_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_63_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_64_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_65_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_66_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_67_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_68_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_user_clock2 (.A(clknet_5_16_0_user_clock2),
    .X(clknet_leaf_69_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_70_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_71_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_72_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_73_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_74_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_75_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_leaf_76_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_77_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_78_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_79_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_80_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_81_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_82_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_83_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_user_clock2 (.A(clknet_5_20_0_user_clock2),
    .X(clknet_leaf_84_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_85_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_86_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_87_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_88_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_user_clock2 (.A(clknet_opt_3_user_clock2),
    .X(clknet_leaf_89_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_90_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_91_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_92_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_leaf_93_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_94_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_95_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_96_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_97_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_98_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_99_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_100_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_101_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_102_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_103_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_user_clock2 (.A(clknet_5_23_0_user_clock2),
    .X(clknet_leaf_104_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_105_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_106_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_107_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_108_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_109_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_110_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_111_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_112_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_113_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_114_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_115_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_116_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_117_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_118_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_119_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_leaf_121_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_122_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_123_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_user_clock2 (.A(clknet_opt_4_user_clock2),
    .X(clknet_leaf_124_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_125_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_126_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_127_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_128_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_129_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_user_clock2 (.A(clknet_5_19_0_user_clock2),
    .X(clknet_leaf_130_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_131_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_132_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_133_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_134_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_135_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_136_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_137_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_138_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_139_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_140_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_141_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_142_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_144_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_145_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_user_clock2 (.A(clknet_opt_7_user_clock2),
    .X(clknet_leaf_146_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_147_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_148_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_149_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_user_clock2 (.A(clknet_5_25_0_user_clock2),
    .X(clknet_leaf_150_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_151_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_152_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_153_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_user_clock2 (.A(clknet_5_28_0_user_clock2),
    .X(clknet_leaf_154_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_155_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_156_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_157_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_158_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_159_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_160_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_user_clock2 (.A(clknet_5_29_0_user_clock2),
    .X(clknet_leaf_161_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_162_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_163_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_164_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_165_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_166_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_167_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_168_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_169_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_170_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_171_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_172_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_173_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_174_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_175_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_176_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_177_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_user_clock2 (.A(clknet_5_31_0_user_clock2),
    .X(clknet_leaf_178_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_179_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_180_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_user_clock2 (.A(clknet_opt_8_user_clock2),
    .X(clknet_leaf_181_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_182_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_leaf_183_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_184_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_user_clock2 (.A(clknet_opt_5_user_clock2),
    .X(clknet_leaf_185_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_user_clock2 (.A(clknet_opt_6_user_clock2),
    .X(clknet_leaf_186_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_leaf_188_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_189_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_190_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_191_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_192_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_193_user_clock2 (.A(clknet_5_26_0_user_clock2),
    .X(clknet_leaf_193_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_194_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_194_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_195_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_195_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_196_user_clock2 (.A(clknet_5_24_0_user_clock2),
    .X(clknet_leaf_196_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_197_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_197_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_198_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_198_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_199_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_199_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_200_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_200_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_201_user_clock2 (.A(clknet_opt_1_user_clock2),
    .X(clknet_leaf_201_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_202_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_202_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_203_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_203_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_204_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_204_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_205_user_clock2 (.A(clknet_5_14_0_user_clock2),
    .X(clknet_leaf_205_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_206_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_206_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_207_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_207_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_208_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_208_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_209_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_209_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_210_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_210_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_211_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_211_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_212_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_212_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_213_user_clock2 (.A(clknet_5_14_0_user_clock2),
    .X(clknet_leaf_213_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_214_user_clock2 (.A(clknet_5_14_0_user_clock2),
    .X(clknet_leaf_214_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_215_user_clock2 (.A(clknet_5_15_0_user_clock2),
    .X(clknet_leaf_215_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_216_user_clock2 (.A(clknet_5_14_0_user_clock2),
    .X(clknet_leaf_216_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_217_user_clock2 (.A(clknet_5_14_0_user_clock2),
    .X(clknet_leaf_217_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_218_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_218_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_219_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_219_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_220_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_220_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_221_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_221_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_222_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_222_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_223_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_223_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_224_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_224_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_225_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_225_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_226_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_226_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_227_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_227_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_228_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_228_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_229_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_229_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_230_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_230_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_231_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_231_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_232_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_232_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_233_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_233_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_234_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_234_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_235_user_clock2 (.A(clknet_5_10_0_user_clock2),
    .X(clknet_leaf_235_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_236_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_236_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_237_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_237_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_238_user_clock2 (.A(clknet_5_11_0_user_clock2),
    .X(clknet_leaf_238_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_239_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_239_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_240_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_240_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_241_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_241_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_242_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_242_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_243_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_243_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_244_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_244_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_245_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_245_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_246_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_246_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_247_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_247_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_248_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_248_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_249_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_249_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_250_user_clock2 (.A(clknet_5_8_0_user_clock2),
    .X(clknet_leaf_250_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_251_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_251_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_252_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_252_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_253_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_253_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_254_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_254_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_255_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_255_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_256_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_256_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_257_user_clock2 (.A(clknet_5_9_0_user_clock2),
    .X(clknet_leaf_257_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_258_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_258_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_259_user_clock2 (.A(clknet_5_14_0_user_clock2),
    .X(clknet_leaf_259_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_260_user_clock2 (.A(clknet_5_14_0_user_clock2),
    .X(clknet_leaf_260_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_261_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_261_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_262_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_262_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_263_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_263_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_264_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_264_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_265_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_265_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_266_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_266_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_267_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_267_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_268_user_clock2 (.A(clknet_5_12_0_user_clock2),
    .X(clknet_leaf_268_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_269_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_269_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_270_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_270_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_271_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_271_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_272_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_272_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_273_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_273_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_274_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_leaf_274_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_275_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_275_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_276_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_276_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_277_user_clock2 (.A(clknet_5_7_0_user_clock2),
    .X(clknet_leaf_277_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_278_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_278_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_279_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_279_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_280_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_280_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_281_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_281_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_282_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_282_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_283_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_283_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_284_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_284_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_285_user_clock2 (.A(clknet_5_6_0_user_clock2),
    .X(clknet_leaf_285_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_286_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_286_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_287_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_287_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_288_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_288_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_289_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_289_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_290_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_290_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_291_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_291_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_292_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_292_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_293_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_293_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_294_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_294_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_295_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_295_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_296_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_296_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_297_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_297_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_298_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_298_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_299_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_299_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_300_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_300_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_301_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_301_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_302_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_302_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_303_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_303_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_304_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_304_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_305_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_305_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_306_user_clock2 (.A(clknet_5_2_0_user_clock2),
    .X(clknet_leaf_306_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_307_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_307_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_308_user_clock2 (.A(clknet_5_3_0_user_clock2),
    .X(clknet_leaf_308_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_309_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_309_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_310_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_310_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_311_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_311_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_312_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_312_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_313_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_leaf_313_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_314_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_314_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_315_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_315_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_316_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_316_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_317_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_317_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_318_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_318_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_319_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_319_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_320_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_320_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_321_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_321_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_322_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_322_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_323_user_clock2 (.A(clknet_5_0_0_user_clock2),
    .X(clknet_leaf_323_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_user_clock2 (.A(user_clock2),
    .X(clknet_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_0_user_clock2 (.A(clknet_0_user_clock2),
    .X(clknet_1_0_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_0_1_user_clock2 (.A(clknet_1_0_0_user_clock2),
    .X(clknet_1_0_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_0_user_clock2 (.A(clknet_0_user_clock2),
    .X(clknet_1_1_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_1_1_1_user_clock2 (.A(clknet_1_1_0_user_clock2),
    .X(clknet_1_1_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_0_0_user_clock2 (.A(clknet_1_0_1_user_clock2),
    .X(clknet_2_0_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_0_1_user_clock2 (.A(clknet_2_0_0_user_clock2),
    .X(clknet_2_0_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_1_0_user_clock2 (.A(clknet_1_0_1_user_clock2),
    .X(clknet_2_1_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_1_1_user_clock2 (.A(clknet_2_1_0_user_clock2),
    .X(clknet_2_1_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_2_0_user_clock2 (.A(clknet_1_1_1_user_clock2),
    .X(clknet_2_2_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_2_1_user_clock2 (.A(clknet_2_2_0_user_clock2),
    .X(clknet_2_2_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_3_0_user_clock2 (.A(clknet_1_1_1_user_clock2),
    .X(clknet_2_3_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_2_3_1_user_clock2 (.A(clknet_2_3_0_user_clock2),
    .X(clknet_2_3_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_0_0_user_clock2 (.A(clknet_2_0_1_user_clock2),
    .X(clknet_3_0_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_1_0_user_clock2 (.A(clknet_2_0_1_user_clock2),
    .X(clknet_3_1_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_2_0_user_clock2 (.A(clknet_2_1_1_user_clock2),
    .X(clknet_3_2_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_3_0_user_clock2 (.A(clknet_2_1_1_user_clock2),
    .X(clknet_3_3_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_4_0_user_clock2 (.A(clknet_2_2_1_user_clock2),
    .X(clknet_3_4_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_5_0_user_clock2 (.A(clknet_2_2_1_user_clock2),
    .X(clknet_3_5_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_6_0_user_clock2 (.A(clknet_2_3_1_user_clock2),
    .X(clknet_3_6_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_3_7_0_user_clock2 (.A(clknet_2_3_1_user_clock2),
    .X(clknet_3_7_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_0_0_user_clock2 (.A(clknet_3_0_0_user_clock2),
    .X(clknet_4_0_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_1_0_user_clock2 (.A(clknet_3_0_0_user_clock2),
    .X(clknet_4_1_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_2_0_user_clock2 (.A(clknet_3_1_0_user_clock2),
    .X(clknet_4_2_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_3_0_user_clock2 (.A(clknet_3_1_0_user_clock2),
    .X(clknet_4_3_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_4_0_user_clock2 (.A(clknet_3_2_0_user_clock2),
    .X(clknet_4_4_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_5_0_user_clock2 (.A(clknet_3_2_0_user_clock2),
    .X(clknet_4_5_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_6_0_user_clock2 (.A(clknet_3_3_0_user_clock2),
    .X(clknet_4_6_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_7_0_user_clock2 (.A(clknet_3_3_0_user_clock2),
    .X(clknet_4_7_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_8_0_user_clock2 (.A(clknet_3_4_0_user_clock2),
    .X(clknet_4_8_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_9_0_user_clock2 (.A(clknet_3_4_0_user_clock2),
    .X(clknet_4_9_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_10_0_user_clock2 (.A(clknet_3_5_0_user_clock2),
    .X(clknet_4_10_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_11_0_user_clock2 (.A(clknet_3_5_0_user_clock2),
    .X(clknet_4_11_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_12_0_user_clock2 (.A(clknet_3_6_0_user_clock2),
    .X(clknet_4_12_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_13_0_user_clock2 (.A(clknet_3_6_0_user_clock2),
    .X(clknet_4_13_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_14_0_user_clock2 (.A(clknet_3_7_0_user_clock2),
    .X(clknet_4_14_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_4_15_0_user_clock2 (.A(clknet_3_7_0_user_clock2),
    .X(clknet_4_15_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_0_0_user_clock2 (.A(clknet_4_0_0_user_clock2),
    .X(clknet_5_0_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_1_0_user_clock2 (.A(clknet_4_0_0_user_clock2),
    .X(clknet_5_1_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_2_0_user_clock2 (.A(clknet_4_1_0_user_clock2),
    .X(clknet_5_2_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_3_0_user_clock2 (.A(clknet_4_1_0_user_clock2),
    .X(clknet_5_3_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_4_0_user_clock2 (.A(clknet_4_2_0_user_clock2),
    .X(clknet_5_4_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_5_0_user_clock2 (.A(clknet_4_2_0_user_clock2),
    .X(clknet_5_5_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_6_0_user_clock2 (.A(clknet_4_3_0_user_clock2),
    .X(clknet_5_6_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_7_0_user_clock2 (.A(clknet_4_3_0_user_clock2),
    .X(clknet_5_7_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_8_0_user_clock2 (.A(clknet_4_4_0_user_clock2),
    .X(clknet_5_8_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_9_0_user_clock2 (.A(clknet_4_4_0_user_clock2),
    .X(clknet_5_9_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_10_0_user_clock2 (.A(clknet_4_5_0_user_clock2),
    .X(clknet_5_10_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_11_0_user_clock2 (.A(clknet_4_5_0_user_clock2),
    .X(clknet_5_11_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_12_0_user_clock2 (.A(clknet_4_6_0_user_clock2),
    .X(clknet_5_12_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_13_0_user_clock2 (.A(clknet_4_6_0_user_clock2),
    .X(clknet_5_13_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_14_0_user_clock2 (.A(clknet_4_7_0_user_clock2),
    .X(clknet_5_14_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_15_0_user_clock2 (.A(clknet_4_7_0_user_clock2),
    .X(clknet_5_15_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_16_0_user_clock2 (.A(clknet_4_8_0_user_clock2),
    .X(clknet_5_16_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_17_0_user_clock2 (.A(clknet_4_8_0_user_clock2),
    .X(clknet_5_17_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_18_0_user_clock2 (.A(clknet_4_9_0_user_clock2),
    .X(clknet_5_18_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_19_0_user_clock2 (.A(clknet_4_9_0_user_clock2),
    .X(clknet_5_19_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_20_0_user_clock2 (.A(clknet_4_10_0_user_clock2),
    .X(clknet_5_20_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_21_0_user_clock2 (.A(clknet_4_10_0_user_clock2),
    .X(clknet_5_21_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_22_0_user_clock2 (.A(clknet_4_11_0_user_clock2),
    .X(clknet_5_22_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_23_0_user_clock2 (.A(clknet_4_11_0_user_clock2),
    .X(clknet_5_23_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_24_0_user_clock2 (.A(clknet_4_12_0_user_clock2),
    .X(clknet_5_24_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_25_0_user_clock2 (.A(clknet_4_12_0_user_clock2),
    .X(clknet_5_25_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_26_0_user_clock2 (.A(clknet_4_13_0_user_clock2),
    .X(clknet_5_26_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_27_0_user_clock2 (.A(clknet_4_13_0_user_clock2),
    .X(clknet_5_27_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_28_0_user_clock2 (.A(clknet_4_14_0_user_clock2),
    .X(clknet_5_28_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_29_0_user_clock2 (.A(clknet_4_14_0_user_clock2),
    .X(clknet_5_29_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_30_0_user_clock2 (.A(clknet_4_15_0_user_clock2),
    .X(clknet_5_30_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 clkbuf_5_31_0_user_clock2 (.A(clknet_4_15_0_user_clock2),
    .X(clknet_5_31_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_0_user_clock2 (.A(clknet_5_1_0_user_clock2),
    .X(clknet_opt_0_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_user_clock2 (.A(clknet_5_13_0_user_clock2),
    .X(clknet_opt_1_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_user_clock2 (.A(clknet_5_17_0_user_clock2),
    .X(clknet_opt_2_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_3_user_clock2 (.A(clknet_5_21_0_user_clock2),
    .X(clknet_opt_3_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_4_user_clock2 (.A(clknet_5_22_0_user_clock2),
    .X(clknet_opt_4_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_5_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_opt_5_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_6_user_clock2 (.A(clknet_5_27_0_user_clock2),
    .X(clknet_opt_6_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_7_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_opt_7_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_8_user_clock2 (.A(clknet_5_30_0_user_clock2),
    .X(clknet_opt_8_user_clock2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
endmodule
