magic
tech sky130A
magscale 1 2
timestamp 1622193948
<< obsli1 >>
rect 2145 2261 107427 107627
<< obsm1 >>
rect 1104 2128 108178 108304
<< metal2 >>
rect 478 110175 534 110975
rect 938 110175 994 110975
rect 1398 110175 1454 110975
rect 1858 110175 1914 110975
rect 2778 110175 2834 110975
rect 3238 110175 3294 110975
rect 3698 110175 3754 110975
rect 4158 110175 4214 110975
rect 5078 110175 5134 110975
rect 5538 110175 5594 110975
rect 5998 110175 6054 110975
rect 6458 110175 6514 110975
rect 6918 110175 6974 110975
rect 7838 110175 7894 110975
rect 8298 110175 8354 110975
rect 8758 110175 8814 110975
rect 9218 110175 9274 110975
rect 10138 110175 10194 110975
rect 10598 110175 10654 110975
rect 11058 110175 11114 110975
rect 11518 110175 11574 110975
rect 12438 110175 12494 110975
rect 12898 110175 12954 110975
rect 13358 110175 13414 110975
rect 13818 110175 13874 110975
rect 14738 110175 14794 110975
rect 15198 110175 15254 110975
rect 15658 110175 15714 110975
rect 16118 110175 16174 110975
rect 17038 110175 17094 110975
rect 17498 110175 17554 110975
rect 17958 110175 18014 110975
rect 18418 110175 18474 110975
rect 19338 110175 19394 110975
rect 19798 110175 19854 110975
rect 20258 110175 20314 110975
rect 20718 110175 20774 110975
rect 21638 110175 21694 110975
rect 22098 110175 22154 110975
rect 22558 110175 22614 110975
rect 23018 110175 23074 110975
rect 23938 110175 23994 110975
rect 24398 110175 24454 110975
rect 24858 110175 24914 110975
rect 25318 110175 25374 110975
rect 26238 110175 26294 110975
rect 26698 110175 26754 110975
rect 27158 110175 27214 110975
rect 27618 110175 27674 110975
rect 28538 110175 28594 110975
rect 28998 110175 29054 110975
rect 29458 110175 29514 110975
rect 29918 110175 29974 110975
rect 30838 110175 30894 110975
rect 31298 110175 31354 110975
rect 31758 110175 31814 110975
rect 32218 110175 32274 110975
rect 33138 110175 33194 110975
rect 33598 110175 33654 110975
rect 34058 110175 34114 110975
rect 34518 110175 34574 110975
rect 35438 110175 35494 110975
rect 35898 110175 35954 110975
rect 36358 110175 36414 110975
rect 36818 110175 36874 110975
rect 37738 110175 37794 110975
rect 38198 110175 38254 110975
rect 38658 110175 38714 110975
rect 39118 110175 39174 110975
rect 40038 110175 40094 110975
rect 40498 110175 40554 110975
rect 40958 110175 41014 110975
rect 41418 110175 41474 110975
rect 42338 110175 42394 110975
rect 42798 110175 42854 110975
rect 43258 110175 43314 110975
rect 43718 110175 43774 110975
rect 44638 110175 44694 110975
rect 45098 110175 45154 110975
rect 45558 110175 45614 110975
rect 46018 110175 46074 110975
rect 46938 110175 46994 110975
rect 47398 110175 47454 110975
rect 47858 110175 47914 110975
rect 48318 110175 48374 110975
rect 48778 110175 48834 110975
rect 49698 110175 49754 110975
rect 50158 110175 50214 110975
rect 50618 110175 50674 110975
rect 51078 110175 51134 110975
rect 51998 110175 52054 110975
rect 52458 110175 52514 110975
rect 52918 110175 52974 110975
rect 53378 110175 53434 110975
rect 54298 110175 54354 110975
rect 54758 110175 54814 110975
rect 55218 110175 55274 110975
rect 55678 110175 55734 110975
rect 56598 110175 56654 110975
rect 57058 110175 57114 110975
rect 57518 110175 57574 110975
rect 57978 110175 58034 110975
rect 58898 110175 58954 110975
rect 59358 110175 59414 110975
rect 59818 110175 59874 110975
rect 60278 110175 60334 110975
rect 61198 110175 61254 110975
rect 61658 110175 61714 110975
rect 62118 110175 62174 110975
rect 62578 110175 62634 110975
rect 63498 110175 63554 110975
rect 63958 110175 64014 110975
rect 64418 110175 64474 110975
rect 64878 110175 64934 110975
rect 65798 110175 65854 110975
rect 66258 110175 66314 110975
rect 66718 110175 66774 110975
rect 67178 110175 67234 110975
rect 68098 110175 68154 110975
rect 68558 110175 68614 110975
rect 69018 110175 69074 110975
rect 69478 110175 69534 110975
rect 70398 110175 70454 110975
rect 70858 110175 70914 110975
rect 71318 110175 71374 110975
rect 71778 110175 71834 110975
rect 72698 110175 72754 110975
rect 73158 110175 73214 110975
rect 73618 110175 73674 110975
rect 74078 110175 74134 110975
rect 74998 110175 75054 110975
rect 75458 110175 75514 110975
rect 75918 110175 75974 110975
rect 76378 110175 76434 110975
rect 77298 110175 77354 110975
rect 77758 110175 77814 110975
rect 78218 110175 78274 110975
rect 78678 110175 78734 110975
rect 79598 110175 79654 110975
rect 80058 110175 80114 110975
rect 80518 110175 80574 110975
rect 80978 110175 81034 110975
rect 81898 110175 81954 110975
rect 82358 110175 82414 110975
rect 82818 110175 82874 110975
rect 83278 110175 83334 110975
rect 84198 110175 84254 110975
rect 84658 110175 84714 110975
rect 85118 110175 85174 110975
rect 85578 110175 85634 110975
rect 86498 110175 86554 110975
rect 86958 110175 87014 110975
rect 87418 110175 87474 110975
rect 87878 110175 87934 110975
rect 88338 110175 88394 110975
rect 89258 110175 89314 110975
rect 89718 110175 89774 110975
rect 90178 110175 90234 110975
rect 90638 110175 90694 110975
rect 91558 110175 91614 110975
rect 92018 110175 92074 110975
rect 92478 110175 92534 110975
rect 92938 110175 92994 110975
rect 93858 110175 93914 110975
rect 94318 110175 94374 110975
rect 94778 110175 94834 110975
rect 95238 110175 95294 110975
rect 96158 110175 96214 110975
rect 96618 110175 96674 110975
rect 97078 110175 97134 110975
rect 97538 110175 97594 110975
rect 98458 110175 98514 110975
rect 98918 110175 98974 110975
rect 99378 110175 99434 110975
rect 99838 110175 99894 110975
rect 100758 110175 100814 110975
rect 101218 110175 101274 110975
rect 101678 110175 101734 110975
rect 102138 110175 102194 110975
rect 103058 110175 103114 110975
rect 103518 110175 103574 110975
rect 103978 110175 104034 110975
rect 104438 110175 104494 110975
rect 105358 110175 105414 110975
rect 105818 110175 105874 110975
rect 106278 110175 106334 110975
rect 106738 110175 106794 110975
rect 107658 110175 107714 110975
rect 108118 110175 108174 110975
rect 478 0 534 800
rect 938 0 994 800
rect 1398 0 1454 800
rect 1858 0 1914 800
rect 2318 0 2374 800
rect 3238 0 3294 800
rect 3698 0 3754 800
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 6918 0 6974 800
rect 7838 0 7894 800
rect 8298 0 8354 800
rect 8758 0 8814 800
rect 9218 0 9274 800
rect 10138 0 10194 800
rect 10598 0 10654 800
rect 11058 0 11114 800
rect 11518 0 11574 800
rect 12438 0 12494 800
rect 12898 0 12954 800
rect 13358 0 13414 800
rect 13818 0 13874 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 17958 0 18014 800
rect 18418 0 18474 800
rect 19338 0 19394 800
rect 19798 0 19854 800
rect 20258 0 20314 800
rect 20718 0 20774 800
rect 21638 0 21694 800
rect 22098 0 22154 800
rect 22558 0 22614 800
rect 23018 0 23074 800
rect 23938 0 23994 800
rect 24398 0 24454 800
rect 24858 0 24914 800
rect 25318 0 25374 800
rect 26238 0 26294 800
rect 26698 0 26754 800
rect 27158 0 27214 800
rect 27618 0 27674 800
rect 28538 0 28594 800
rect 28998 0 29054 800
rect 29458 0 29514 800
rect 29918 0 29974 800
rect 30838 0 30894 800
rect 31298 0 31354 800
rect 31758 0 31814 800
rect 32218 0 32274 800
rect 33138 0 33194 800
rect 33598 0 33654 800
rect 34058 0 34114 800
rect 34518 0 34574 800
rect 35438 0 35494 800
rect 35898 0 35954 800
rect 36358 0 36414 800
rect 36818 0 36874 800
rect 37738 0 37794 800
rect 38198 0 38254 800
rect 38658 0 38714 800
rect 39118 0 39174 800
rect 40038 0 40094 800
rect 40498 0 40554 800
rect 40958 0 41014 800
rect 41418 0 41474 800
rect 41878 0 41934 800
rect 42798 0 42854 800
rect 43258 0 43314 800
rect 43718 0 43774 800
rect 44178 0 44234 800
rect 45098 0 45154 800
rect 45558 0 45614 800
rect 46018 0 46074 800
rect 46478 0 46534 800
rect 47398 0 47454 800
rect 47858 0 47914 800
rect 48318 0 48374 800
rect 48778 0 48834 800
rect 49698 0 49754 800
rect 50158 0 50214 800
rect 50618 0 50674 800
rect 51078 0 51134 800
rect 51998 0 52054 800
rect 52458 0 52514 800
rect 52918 0 52974 800
rect 53378 0 53434 800
rect 54298 0 54354 800
rect 54758 0 54814 800
rect 55218 0 55274 800
rect 55678 0 55734 800
rect 56598 0 56654 800
rect 57058 0 57114 800
rect 57518 0 57574 800
rect 57978 0 58034 800
rect 58898 0 58954 800
rect 59358 0 59414 800
rect 59818 0 59874 800
rect 60278 0 60334 800
rect 61198 0 61254 800
rect 61658 0 61714 800
rect 62118 0 62174 800
rect 62578 0 62634 800
rect 63498 0 63554 800
rect 63958 0 64014 800
rect 64418 0 64474 800
rect 64878 0 64934 800
rect 65798 0 65854 800
rect 66258 0 66314 800
rect 66718 0 66774 800
rect 67178 0 67234 800
rect 68098 0 68154 800
rect 68558 0 68614 800
rect 69018 0 69074 800
rect 69478 0 69534 800
rect 70398 0 70454 800
rect 70858 0 70914 800
rect 71318 0 71374 800
rect 71778 0 71834 800
rect 72698 0 72754 800
rect 73158 0 73214 800
rect 73618 0 73674 800
rect 74078 0 74134 800
rect 74998 0 75054 800
rect 75458 0 75514 800
rect 75918 0 75974 800
rect 76378 0 76434 800
rect 77298 0 77354 800
rect 77758 0 77814 800
rect 78218 0 78274 800
rect 78678 0 78734 800
rect 79598 0 79654 800
rect 80058 0 80114 800
rect 80518 0 80574 800
rect 80978 0 81034 800
rect 81438 0 81494 800
rect 82358 0 82414 800
rect 82818 0 82874 800
rect 83278 0 83334 800
rect 83738 0 83794 800
rect 84658 0 84714 800
rect 85118 0 85174 800
rect 85578 0 85634 800
rect 86038 0 86094 800
rect 86958 0 87014 800
rect 87418 0 87474 800
rect 87878 0 87934 800
rect 88338 0 88394 800
rect 89258 0 89314 800
rect 89718 0 89774 800
rect 90178 0 90234 800
rect 90638 0 90694 800
rect 91558 0 91614 800
rect 92018 0 92074 800
rect 92478 0 92534 800
rect 92938 0 92994 800
rect 93858 0 93914 800
rect 94318 0 94374 800
rect 94778 0 94834 800
rect 95238 0 95294 800
rect 96158 0 96214 800
rect 96618 0 96674 800
rect 97078 0 97134 800
rect 97538 0 97594 800
rect 98458 0 98514 800
rect 98918 0 98974 800
rect 99378 0 99434 800
rect 99838 0 99894 800
rect 100758 0 100814 800
rect 101218 0 101274 800
rect 101678 0 101734 800
rect 102138 0 102194 800
rect 103058 0 103114 800
rect 103518 0 103574 800
rect 103978 0 104034 800
rect 104438 0 104494 800
rect 105358 0 105414 800
rect 105818 0 105874 800
rect 106278 0 106334 800
rect 106738 0 106794 800
rect 107658 0 107714 800
rect 108118 0 108174 800
<< obsm2 >>
rect 1510 110119 1802 110265
rect 1970 110119 2722 110265
rect 2890 110119 3182 110265
rect 3350 110119 3642 110265
rect 3810 110119 4102 110265
rect 4270 110119 5022 110265
rect 5190 110119 5482 110265
rect 5650 110119 5942 110265
rect 6110 110119 6402 110265
rect 6570 110119 6862 110265
rect 7030 110119 7782 110265
rect 7950 110119 8242 110265
rect 8410 110119 8702 110265
rect 8870 110119 9162 110265
rect 9330 110119 10082 110265
rect 10250 110119 10542 110265
rect 10710 110119 11002 110265
rect 11170 110119 11462 110265
rect 11630 110119 12382 110265
rect 12550 110119 12842 110265
rect 13010 110119 13302 110265
rect 13470 110119 13762 110265
rect 13930 110119 14682 110265
rect 14850 110119 15142 110265
rect 15310 110119 15602 110265
rect 15770 110119 16062 110265
rect 16230 110119 16982 110265
rect 17150 110119 17442 110265
rect 17610 110119 17902 110265
rect 18070 110119 18362 110265
rect 18530 110119 19282 110265
rect 19450 110119 19742 110265
rect 19910 110119 20202 110265
rect 20370 110119 20662 110265
rect 20830 110119 21582 110265
rect 21750 110119 22042 110265
rect 22210 110119 22502 110265
rect 22670 110119 22962 110265
rect 23130 110119 23882 110265
rect 24050 110119 24342 110265
rect 24510 110119 24802 110265
rect 24970 110119 25262 110265
rect 25430 110119 26182 110265
rect 26350 110119 26642 110265
rect 26810 110119 27102 110265
rect 27270 110119 27562 110265
rect 27730 110119 28482 110265
rect 28650 110119 28942 110265
rect 29110 110119 29402 110265
rect 29570 110119 29862 110265
rect 30030 110119 30782 110265
rect 30950 110119 31242 110265
rect 31410 110119 31702 110265
rect 31870 110119 32162 110265
rect 32330 110119 33082 110265
rect 33250 110119 33542 110265
rect 33710 110119 34002 110265
rect 34170 110119 34462 110265
rect 34630 110119 35382 110265
rect 35550 110119 35842 110265
rect 36010 110119 36302 110265
rect 36470 110119 36762 110265
rect 36930 110119 37682 110265
rect 37850 110119 38142 110265
rect 38310 110119 38602 110265
rect 38770 110119 39062 110265
rect 39230 110119 39982 110265
rect 40150 110119 40442 110265
rect 40610 110119 40902 110265
rect 41070 110119 41362 110265
rect 41530 110119 42282 110265
rect 42450 110119 42742 110265
rect 42910 110119 43202 110265
rect 43370 110119 43662 110265
rect 43830 110119 44582 110265
rect 44750 110119 45042 110265
rect 45210 110119 45502 110265
rect 45670 110119 45962 110265
rect 46130 110119 46882 110265
rect 47050 110119 47342 110265
rect 47510 110119 47802 110265
rect 47970 110119 48262 110265
rect 48430 110119 48722 110265
rect 48890 110119 49642 110265
rect 49810 110119 50102 110265
rect 50270 110119 50562 110265
rect 50730 110119 51022 110265
rect 51190 110119 51942 110265
rect 52110 110119 52402 110265
rect 52570 110119 52862 110265
rect 53030 110119 53322 110265
rect 53490 110119 54242 110265
rect 54410 110119 54702 110265
rect 54870 110119 55162 110265
rect 55330 110119 55622 110265
rect 55790 110119 56542 110265
rect 56710 110119 57002 110265
rect 57170 110119 57462 110265
rect 57630 110119 57922 110265
rect 58090 110119 58842 110265
rect 59010 110119 59302 110265
rect 59470 110119 59762 110265
rect 59930 110119 60222 110265
rect 60390 110119 61142 110265
rect 61310 110119 61602 110265
rect 61770 110119 62062 110265
rect 62230 110119 62522 110265
rect 62690 110119 63442 110265
rect 63610 110119 63902 110265
rect 64070 110119 64362 110265
rect 64530 110119 64822 110265
rect 64990 110119 65742 110265
rect 65910 110119 66202 110265
rect 66370 110119 66662 110265
rect 66830 110119 67122 110265
rect 67290 110119 68042 110265
rect 68210 110119 68502 110265
rect 68670 110119 68962 110265
rect 69130 110119 69422 110265
rect 69590 110119 70342 110265
rect 70510 110119 70802 110265
rect 70970 110119 71262 110265
rect 71430 110119 71722 110265
rect 71890 110119 72642 110265
rect 72810 110119 73102 110265
rect 73270 110119 73562 110265
rect 73730 110119 74022 110265
rect 74190 110119 74942 110265
rect 75110 110119 75402 110265
rect 75570 110119 75862 110265
rect 76030 110119 76322 110265
rect 76490 110119 77242 110265
rect 77410 110119 77702 110265
rect 77870 110119 78162 110265
rect 78330 110119 78622 110265
rect 78790 110119 79542 110265
rect 79710 110119 80002 110265
rect 80170 110119 80462 110265
rect 80630 110119 80922 110265
rect 81090 110119 81842 110265
rect 82010 110119 82302 110265
rect 82470 110119 82762 110265
rect 82930 110119 83222 110265
rect 83390 110119 84142 110265
rect 84310 110119 84602 110265
rect 84770 110119 85062 110265
rect 85230 110119 85522 110265
rect 85690 110119 86442 110265
rect 86610 110119 86902 110265
rect 87070 110119 87362 110265
rect 87530 110119 87822 110265
rect 87990 110119 88282 110265
rect 88450 110119 89202 110265
rect 89370 110119 89662 110265
rect 89830 110119 90122 110265
rect 90290 110119 90582 110265
rect 90750 110119 91502 110265
rect 91670 110119 91962 110265
rect 92130 110119 92422 110265
rect 92590 110119 92882 110265
rect 93050 110119 93802 110265
rect 93970 110119 94262 110265
rect 94430 110119 94722 110265
rect 94890 110119 95182 110265
rect 95350 110119 96102 110265
rect 96270 110119 96562 110265
rect 96730 110119 97022 110265
rect 97190 110119 97482 110265
rect 97650 110119 98402 110265
rect 98570 110119 98862 110265
rect 99030 110119 99322 110265
rect 99490 110119 99782 110265
rect 99950 110119 100702 110265
rect 100870 110119 101162 110265
rect 101330 110119 101622 110265
rect 101790 110119 102082 110265
rect 102250 110119 103002 110265
rect 103170 110119 103462 110265
rect 103630 110119 103922 110265
rect 104090 110119 104382 110265
rect 104550 110119 105302 110265
rect 105470 110119 105762 110265
rect 105930 110119 106222 110265
rect 106390 110119 106682 110265
rect 106850 110119 107602 110265
rect 107770 110119 108062 110265
rect 1400 856 108172 110119
rect 1510 711 1802 856
rect 1970 711 2262 856
rect 2430 711 3182 856
rect 3350 711 3642 856
rect 3810 711 4102 856
rect 4270 711 4562 856
rect 4730 711 5482 856
rect 5650 711 5942 856
rect 6110 711 6402 856
rect 6570 711 6862 856
rect 7030 711 7782 856
rect 7950 711 8242 856
rect 8410 711 8702 856
rect 8870 711 9162 856
rect 9330 711 10082 856
rect 10250 711 10542 856
rect 10710 711 11002 856
rect 11170 711 11462 856
rect 11630 711 12382 856
rect 12550 711 12842 856
rect 13010 711 13302 856
rect 13470 711 13762 856
rect 13930 711 14682 856
rect 14850 711 15142 856
rect 15310 711 15602 856
rect 15770 711 16062 856
rect 16230 711 16982 856
rect 17150 711 17442 856
rect 17610 711 17902 856
rect 18070 711 18362 856
rect 18530 711 19282 856
rect 19450 711 19742 856
rect 19910 711 20202 856
rect 20370 711 20662 856
rect 20830 711 21582 856
rect 21750 711 22042 856
rect 22210 711 22502 856
rect 22670 711 22962 856
rect 23130 711 23882 856
rect 24050 711 24342 856
rect 24510 711 24802 856
rect 24970 711 25262 856
rect 25430 711 26182 856
rect 26350 711 26642 856
rect 26810 711 27102 856
rect 27270 711 27562 856
rect 27730 711 28482 856
rect 28650 711 28942 856
rect 29110 711 29402 856
rect 29570 711 29862 856
rect 30030 711 30782 856
rect 30950 711 31242 856
rect 31410 711 31702 856
rect 31870 711 32162 856
rect 32330 711 33082 856
rect 33250 711 33542 856
rect 33710 711 34002 856
rect 34170 711 34462 856
rect 34630 711 35382 856
rect 35550 711 35842 856
rect 36010 711 36302 856
rect 36470 711 36762 856
rect 36930 711 37682 856
rect 37850 711 38142 856
rect 38310 711 38602 856
rect 38770 711 39062 856
rect 39230 711 39982 856
rect 40150 711 40442 856
rect 40610 711 40902 856
rect 41070 711 41362 856
rect 41530 711 41822 856
rect 41990 711 42742 856
rect 42910 711 43202 856
rect 43370 711 43662 856
rect 43830 711 44122 856
rect 44290 711 45042 856
rect 45210 711 45502 856
rect 45670 711 45962 856
rect 46130 711 46422 856
rect 46590 711 47342 856
rect 47510 711 47802 856
rect 47970 711 48262 856
rect 48430 711 48722 856
rect 48890 711 49642 856
rect 49810 711 50102 856
rect 50270 711 50562 856
rect 50730 711 51022 856
rect 51190 711 51942 856
rect 52110 711 52402 856
rect 52570 711 52862 856
rect 53030 711 53322 856
rect 53490 711 54242 856
rect 54410 711 54702 856
rect 54870 711 55162 856
rect 55330 711 55622 856
rect 55790 711 56542 856
rect 56710 711 57002 856
rect 57170 711 57462 856
rect 57630 711 57922 856
rect 58090 711 58842 856
rect 59010 711 59302 856
rect 59470 711 59762 856
rect 59930 711 60222 856
rect 60390 711 61142 856
rect 61310 711 61602 856
rect 61770 711 62062 856
rect 62230 711 62522 856
rect 62690 711 63442 856
rect 63610 711 63902 856
rect 64070 711 64362 856
rect 64530 711 64822 856
rect 64990 711 65742 856
rect 65910 711 66202 856
rect 66370 711 66662 856
rect 66830 711 67122 856
rect 67290 711 68042 856
rect 68210 711 68502 856
rect 68670 711 68962 856
rect 69130 711 69422 856
rect 69590 711 70342 856
rect 70510 711 70802 856
rect 70970 711 71262 856
rect 71430 711 71722 856
rect 71890 711 72642 856
rect 72810 711 73102 856
rect 73270 711 73562 856
rect 73730 711 74022 856
rect 74190 711 74942 856
rect 75110 711 75402 856
rect 75570 711 75862 856
rect 76030 711 76322 856
rect 76490 711 77242 856
rect 77410 711 77702 856
rect 77870 711 78162 856
rect 78330 711 78622 856
rect 78790 711 79542 856
rect 79710 711 80002 856
rect 80170 711 80462 856
rect 80630 711 80922 856
rect 81090 711 81382 856
rect 81550 711 82302 856
rect 82470 711 82762 856
rect 82930 711 83222 856
rect 83390 711 83682 856
rect 83850 711 84602 856
rect 84770 711 85062 856
rect 85230 711 85522 856
rect 85690 711 85982 856
rect 86150 711 86902 856
rect 87070 711 87362 856
rect 87530 711 87822 856
rect 87990 711 88282 856
rect 88450 711 89202 856
rect 89370 711 89662 856
rect 89830 711 90122 856
rect 90290 711 90582 856
rect 90750 711 91502 856
rect 91670 711 91962 856
rect 92130 711 92422 856
rect 92590 711 92882 856
rect 93050 711 93802 856
rect 93970 711 94262 856
rect 94430 711 94722 856
rect 94890 711 95182 856
rect 95350 711 96102 856
rect 96270 711 96562 856
rect 96730 711 97022 856
rect 97190 711 97482 856
rect 97650 711 98402 856
rect 98570 711 98862 856
rect 99030 711 99322 856
rect 99490 711 99782 856
rect 99950 711 100702 856
rect 100870 711 101162 856
rect 101330 711 101622 856
rect 101790 711 102082 856
rect 102250 711 103002 856
rect 103170 711 103462 856
rect 103630 711 103922 856
rect 104090 711 104382 856
rect 104550 711 105302 856
rect 105470 711 105762 856
rect 105930 711 106222 856
rect 106390 711 106682 856
rect 106850 711 107602 856
rect 107770 711 108062 856
<< metal3 >>
rect 108031 110168 108831 110288
rect 0 109488 800 109608
rect 108031 109488 108831 109608
rect 0 108808 800 108928
rect 0 108128 800 108248
rect 108031 108128 108831 108248
rect 0 107448 800 107568
rect 108031 107448 108831 107568
rect 108031 106768 108831 106888
rect 0 106088 800 106208
rect 108031 106088 108831 106208
rect 0 105408 800 105528
rect 0 104728 800 104848
rect 108031 104728 108831 104848
rect 0 104048 800 104168
rect 108031 104048 108831 104168
rect 108031 103368 108831 103488
rect 0 102688 800 102808
rect 108031 102688 108831 102808
rect 0 102008 800 102128
rect 0 101328 800 101448
rect 108031 101328 108831 101448
rect 0 100648 800 100768
rect 108031 100648 108831 100768
rect 108031 99968 108831 100088
rect 0 99288 800 99408
rect 108031 99288 108831 99408
rect 0 98608 800 98728
rect 0 97928 800 98048
rect 108031 97928 108831 98048
rect 0 97248 800 97368
rect 108031 97248 108831 97368
rect 108031 96568 108831 96688
rect 0 95888 800 96008
rect 108031 95888 108831 96008
rect 0 95208 800 95328
rect 0 94528 800 94648
rect 108031 94528 108831 94648
rect 0 93848 800 93968
rect 108031 93848 108831 93968
rect 108031 93168 108831 93288
rect 0 92488 800 92608
rect 108031 92488 108831 92608
rect 0 91808 800 91928
rect 0 91128 800 91248
rect 108031 91128 108831 91248
rect 0 90448 800 90568
rect 108031 90448 108831 90568
rect 108031 89768 108831 89888
rect 0 89088 800 89208
rect 108031 89088 108831 89208
rect 0 88408 800 88528
rect 0 87728 800 87848
rect 108031 87728 108831 87848
rect 0 87048 800 87168
rect 108031 87048 108831 87168
rect 108031 86368 108831 86488
rect 0 85688 800 85808
rect 108031 85688 108831 85808
rect 0 85008 800 85128
rect 0 84328 800 84448
rect 108031 84328 108831 84448
rect 0 83648 800 83768
rect 108031 83648 108831 83768
rect 108031 82968 108831 83088
rect 0 82288 800 82408
rect 108031 82288 108831 82408
rect 0 81608 800 81728
rect 0 80928 800 81048
rect 108031 80928 108831 81048
rect 0 80248 800 80368
rect 108031 80248 108831 80368
rect 108031 79568 108831 79688
rect 0 78888 800 79008
rect 108031 78888 108831 79008
rect 0 78208 800 78328
rect 108031 78208 108831 78328
rect 0 77528 800 77648
rect 0 76848 800 76968
rect 108031 76848 108831 76968
rect 108031 76168 108831 76288
rect 0 75488 800 75608
rect 108031 75488 108831 75608
rect 0 74808 800 74928
rect 108031 74808 108831 74928
rect 0 74128 800 74248
rect 0 73448 800 73568
rect 108031 73448 108831 73568
rect 108031 72768 108831 72888
rect 0 72088 800 72208
rect 108031 72088 108831 72208
rect 0 71408 800 71528
rect 108031 71408 108831 71528
rect 0 70728 800 70848
rect 0 70048 800 70168
rect 108031 70048 108831 70168
rect 108031 69368 108831 69488
rect 0 68688 800 68808
rect 108031 68688 108831 68808
rect 0 68008 800 68128
rect 108031 68008 108831 68128
rect 0 67328 800 67448
rect 0 66648 800 66768
rect 108031 66648 108831 66768
rect 108031 65968 108831 66088
rect 0 65288 800 65408
rect 108031 65288 108831 65408
rect 0 64608 800 64728
rect 108031 64608 108831 64728
rect 0 63928 800 64048
rect 0 63248 800 63368
rect 108031 63248 108831 63368
rect 108031 62568 108831 62688
rect 0 61888 800 62008
rect 108031 61888 108831 62008
rect 0 61208 800 61328
rect 108031 61208 108831 61328
rect 0 60528 800 60648
rect 0 59848 800 59968
rect 108031 59848 108831 59968
rect 0 59168 800 59288
rect 108031 59168 108831 59288
rect 108031 58488 108831 58608
rect 0 57808 800 57928
rect 108031 57808 108831 57928
rect 0 57128 800 57248
rect 0 56448 800 56568
rect 108031 56448 108831 56568
rect 0 55768 800 55888
rect 108031 55768 108831 55888
rect 108031 55088 108831 55208
rect 0 54408 800 54528
rect 108031 54408 108831 54528
rect 0 53728 800 53848
rect 0 53048 800 53168
rect 108031 53048 108831 53168
rect 0 52368 800 52488
rect 108031 52368 108831 52488
rect 108031 51688 108831 51808
rect 0 51008 800 51128
rect 108031 51008 108831 51128
rect 0 50328 800 50448
rect 0 49648 800 49768
rect 108031 49648 108831 49768
rect 0 48968 800 49088
rect 108031 48968 108831 49088
rect 108031 48288 108831 48408
rect 0 47608 800 47728
rect 108031 47608 108831 47728
rect 0 46928 800 47048
rect 0 46248 800 46368
rect 108031 46248 108831 46368
rect 0 45568 800 45688
rect 108031 45568 108831 45688
rect 108031 44888 108831 45008
rect 0 44208 800 44328
rect 108031 44208 108831 44328
rect 0 43528 800 43648
rect 0 42848 800 42968
rect 108031 42848 108831 42968
rect 0 42168 800 42288
rect 108031 42168 108831 42288
rect 108031 41488 108831 41608
rect 0 40808 800 40928
rect 108031 40808 108831 40928
rect 0 40128 800 40248
rect 0 39448 800 39568
rect 108031 39448 108831 39568
rect 0 38768 800 38888
rect 108031 38768 108831 38888
rect 108031 38088 108831 38208
rect 0 37408 800 37528
rect 108031 37408 108831 37528
rect 0 36728 800 36848
rect 0 36048 800 36168
rect 108031 36048 108831 36168
rect 0 35368 800 35488
rect 108031 35368 108831 35488
rect 108031 34688 108831 34808
rect 0 34008 800 34128
rect 108031 34008 108831 34128
rect 0 33328 800 33448
rect 0 32648 800 32768
rect 108031 32648 108831 32768
rect 0 31968 800 32088
rect 108031 31968 108831 32088
rect 108031 31288 108831 31408
rect 0 30608 800 30728
rect 108031 30608 108831 30728
rect 0 29928 800 30048
rect 0 29248 800 29368
rect 108031 29248 108831 29368
rect 0 28568 800 28688
rect 108031 28568 108831 28688
rect 108031 27888 108831 28008
rect 0 27208 800 27328
rect 108031 27208 108831 27328
rect 0 26528 800 26648
rect 0 25848 800 25968
rect 108031 25848 108831 25968
rect 0 25168 800 25288
rect 108031 25168 108831 25288
rect 108031 24488 108831 24608
rect 0 23808 800 23928
rect 108031 23808 108831 23928
rect 0 23128 800 23248
rect 0 22448 800 22568
rect 108031 22448 108831 22568
rect 0 21768 800 21888
rect 108031 21768 108831 21888
rect 108031 21088 108831 21208
rect 0 20408 800 20528
rect 108031 20408 108831 20528
rect 0 19728 800 19848
rect 108031 19728 108831 19848
rect 0 19048 800 19168
rect 0 18368 800 18488
rect 108031 18368 108831 18488
rect 108031 17688 108831 17808
rect 0 17008 800 17128
rect 108031 17008 108831 17128
rect 0 16328 800 16448
rect 108031 16328 108831 16448
rect 0 15648 800 15768
rect 0 14968 800 15088
rect 108031 14968 108831 15088
rect 108031 14288 108831 14408
rect 0 13608 800 13728
rect 108031 13608 108831 13728
rect 0 12928 800 13048
rect 108031 12928 108831 13048
rect 0 12248 800 12368
rect 0 11568 800 11688
rect 108031 11568 108831 11688
rect 108031 10888 108831 11008
rect 0 10208 800 10328
rect 108031 10208 108831 10328
rect 0 9528 800 9648
rect 108031 9528 108831 9648
rect 0 8848 800 8968
rect 0 8168 800 8288
rect 108031 8168 108831 8288
rect 108031 7488 108831 7608
rect 0 6808 800 6928
rect 108031 6808 108831 6928
rect 0 6128 800 6248
rect 108031 6128 108831 6248
rect 0 5448 800 5568
rect 0 4768 800 4888
rect 108031 4768 108831 4888
rect 108031 4088 108831 4208
rect 0 3408 800 3528
rect 108031 3408 108831 3528
rect 0 2728 800 2848
rect 108031 2728 108831 2848
rect 0 2048 800 2168
rect 0 1368 800 1488
rect 108031 1368 108831 1488
rect 108031 688 108831 808
<< obsm3 >>
rect 800 110088 107951 110261
rect 800 109688 108031 110088
rect 880 109408 107951 109688
rect 800 109008 108031 109408
rect 880 108728 108031 109008
rect 800 108328 108031 108728
rect 880 108048 107951 108328
rect 800 107648 108031 108048
rect 880 107368 107951 107648
rect 800 106968 108031 107368
rect 800 106688 107951 106968
rect 800 106288 108031 106688
rect 880 106008 107951 106288
rect 800 105608 108031 106008
rect 880 105328 108031 105608
rect 800 104928 108031 105328
rect 880 104648 107951 104928
rect 800 104248 108031 104648
rect 880 103968 107951 104248
rect 800 103568 108031 103968
rect 800 103288 107951 103568
rect 800 102888 108031 103288
rect 880 102608 107951 102888
rect 800 102208 108031 102608
rect 880 101928 108031 102208
rect 800 101528 108031 101928
rect 880 101248 107951 101528
rect 800 100848 108031 101248
rect 880 100568 107951 100848
rect 800 100168 108031 100568
rect 800 99888 107951 100168
rect 800 99488 108031 99888
rect 880 99208 107951 99488
rect 800 98808 108031 99208
rect 880 98528 108031 98808
rect 800 98128 108031 98528
rect 880 97848 107951 98128
rect 800 97448 108031 97848
rect 880 97168 107951 97448
rect 800 96768 108031 97168
rect 800 96488 107951 96768
rect 800 96088 108031 96488
rect 880 95808 107951 96088
rect 800 95408 108031 95808
rect 880 95128 108031 95408
rect 800 94728 108031 95128
rect 880 94448 107951 94728
rect 800 94048 108031 94448
rect 880 93768 107951 94048
rect 800 93368 108031 93768
rect 800 93088 107951 93368
rect 800 92688 108031 93088
rect 880 92408 107951 92688
rect 800 92008 108031 92408
rect 880 91728 108031 92008
rect 800 91328 108031 91728
rect 880 91048 107951 91328
rect 800 90648 108031 91048
rect 880 90368 107951 90648
rect 800 89968 108031 90368
rect 800 89688 107951 89968
rect 800 89288 108031 89688
rect 880 89008 107951 89288
rect 800 88608 108031 89008
rect 880 88328 108031 88608
rect 800 87928 108031 88328
rect 880 87648 107951 87928
rect 800 87248 108031 87648
rect 880 86968 107951 87248
rect 800 86568 108031 86968
rect 800 86288 107951 86568
rect 800 85888 108031 86288
rect 880 85608 107951 85888
rect 800 85208 108031 85608
rect 880 84928 108031 85208
rect 800 84528 108031 84928
rect 880 84248 107951 84528
rect 800 83848 108031 84248
rect 880 83568 107951 83848
rect 800 83168 108031 83568
rect 800 82888 107951 83168
rect 800 82488 108031 82888
rect 880 82208 107951 82488
rect 800 81808 108031 82208
rect 880 81528 108031 81808
rect 800 81128 108031 81528
rect 880 80848 107951 81128
rect 800 80448 108031 80848
rect 880 80168 107951 80448
rect 800 79768 108031 80168
rect 800 79488 107951 79768
rect 800 79088 108031 79488
rect 880 78808 107951 79088
rect 800 78408 108031 78808
rect 880 78128 107951 78408
rect 800 77728 108031 78128
rect 880 77448 108031 77728
rect 800 77048 108031 77448
rect 880 76768 107951 77048
rect 800 76368 108031 76768
rect 800 76088 107951 76368
rect 800 75688 108031 76088
rect 880 75408 107951 75688
rect 800 75008 108031 75408
rect 880 74728 107951 75008
rect 800 74328 108031 74728
rect 880 74048 108031 74328
rect 800 73648 108031 74048
rect 880 73368 107951 73648
rect 800 72968 108031 73368
rect 800 72688 107951 72968
rect 800 72288 108031 72688
rect 880 72008 107951 72288
rect 800 71608 108031 72008
rect 880 71328 107951 71608
rect 800 70928 108031 71328
rect 880 70648 108031 70928
rect 800 70248 108031 70648
rect 880 69968 107951 70248
rect 800 69568 108031 69968
rect 800 69288 107951 69568
rect 800 68888 108031 69288
rect 880 68608 107951 68888
rect 800 68208 108031 68608
rect 880 67928 107951 68208
rect 800 67528 108031 67928
rect 880 67248 108031 67528
rect 800 66848 108031 67248
rect 880 66568 107951 66848
rect 800 66168 108031 66568
rect 800 65888 107951 66168
rect 800 65488 108031 65888
rect 880 65208 107951 65488
rect 800 64808 108031 65208
rect 880 64528 107951 64808
rect 800 64128 108031 64528
rect 880 63848 108031 64128
rect 800 63448 108031 63848
rect 880 63168 107951 63448
rect 800 62768 108031 63168
rect 800 62488 107951 62768
rect 800 62088 108031 62488
rect 880 61808 107951 62088
rect 800 61408 108031 61808
rect 880 61128 107951 61408
rect 800 60728 108031 61128
rect 880 60448 108031 60728
rect 800 60048 108031 60448
rect 880 59768 107951 60048
rect 800 59368 108031 59768
rect 880 59088 107951 59368
rect 800 58688 108031 59088
rect 800 58408 107951 58688
rect 800 58008 108031 58408
rect 880 57728 107951 58008
rect 800 57328 108031 57728
rect 880 57048 108031 57328
rect 800 56648 108031 57048
rect 880 56368 107951 56648
rect 800 55968 108031 56368
rect 880 55688 107951 55968
rect 800 55288 108031 55688
rect 800 55008 107951 55288
rect 800 54608 108031 55008
rect 880 54328 107951 54608
rect 800 53928 108031 54328
rect 880 53648 108031 53928
rect 800 53248 108031 53648
rect 880 52968 107951 53248
rect 800 52568 108031 52968
rect 880 52288 107951 52568
rect 800 51888 108031 52288
rect 800 51608 107951 51888
rect 800 51208 108031 51608
rect 880 50928 107951 51208
rect 800 50528 108031 50928
rect 880 50248 108031 50528
rect 800 49848 108031 50248
rect 880 49568 107951 49848
rect 800 49168 108031 49568
rect 880 48888 107951 49168
rect 800 48488 108031 48888
rect 800 48208 107951 48488
rect 800 47808 108031 48208
rect 880 47528 107951 47808
rect 800 47128 108031 47528
rect 880 46848 108031 47128
rect 800 46448 108031 46848
rect 880 46168 107951 46448
rect 800 45768 108031 46168
rect 880 45488 107951 45768
rect 800 45088 108031 45488
rect 800 44808 107951 45088
rect 800 44408 108031 44808
rect 880 44128 107951 44408
rect 800 43728 108031 44128
rect 880 43448 108031 43728
rect 800 43048 108031 43448
rect 880 42768 107951 43048
rect 800 42368 108031 42768
rect 880 42088 107951 42368
rect 800 41688 108031 42088
rect 800 41408 107951 41688
rect 800 41008 108031 41408
rect 880 40728 107951 41008
rect 800 40328 108031 40728
rect 880 40048 108031 40328
rect 800 39648 108031 40048
rect 880 39368 107951 39648
rect 800 38968 108031 39368
rect 880 38688 107951 38968
rect 800 38288 108031 38688
rect 800 38008 107951 38288
rect 800 37608 108031 38008
rect 880 37328 107951 37608
rect 800 36928 108031 37328
rect 880 36648 108031 36928
rect 800 36248 108031 36648
rect 880 35968 107951 36248
rect 800 35568 108031 35968
rect 880 35288 107951 35568
rect 800 34888 108031 35288
rect 800 34608 107951 34888
rect 800 34208 108031 34608
rect 880 33928 107951 34208
rect 800 33528 108031 33928
rect 880 33248 108031 33528
rect 800 32848 108031 33248
rect 880 32568 107951 32848
rect 800 32168 108031 32568
rect 880 31888 107951 32168
rect 800 31488 108031 31888
rect 800 31208 107951 31488
rect 800 30808 108031 31208
rect 880 30528 107951 30808
rect 800 30128 108031 30528
rect 880 29848 108031 30128
rect 800 29448 108031 29848
rect 880 29168 107951 29448
rect 800 28768 108031 29168
rect 880 28488 107951 28768
rect 800 28088 108031 28488
rect 800 27808 107951 28088
rect 800 27408 108031 27808
rect 880 27128 107951 27408
rect 800 26728 108031 27128
rect 880 26448 108031 26728
rect 800 26048 108031 26448
rect 880 25768 107951 26048
rect 800 25368 108031 25768
rect 880 25088 107951 25368
rect 800 24688 108031 25088
rect 800 24408 107951 24688
rect 800 24008 108031 24408
rect 880 23728 107951 24008
rect 800 23328 108031 23728
rect 880 23048 108031 23328
rect 800 22648 108031 23048
rect 880 22368 107951 22648
rect 800 21968 108031 22368
rect 880 21688 107951 21968
rect 800 21288 108031 21688
rect 800 21008 107951 21288
rect 800 20608 108031 21008
rect 880 20328 107951 20608
rect 800 19928 108031 20328
rect 880 19648 107951 19928
rect 800 19248 108031 19648
rect 880 18968 108031 19248
rect 800 18568 108031 18968
rect 880 18288 107951 18568
rect 800 17888 108031 18288
rect 800 17608 107951 17888
rect 800 17208 108031 17608
rect 880 16928 107951 17208
rect 800 16528 108031 16928
rect 880 16248 107951 16528
rect 800 15848 108031 16248
rect 880 15568 108031 15848
rect 800 15168 108031 15568
rect 880 14888 107951 15168
rect 800 14488 108031 14888
rect 800 14208 107951 14488
rect 800 13808 108031 14208
rect 880 13528 107951 13808
rect 800 13128 108031 13528
rect 880 12848 107951 13128
rect 800 12448 108031 12848
rect 880 12168 108031 12448
rect 800 11768 108031 12168
rect 880 11488 107951 11768
rect 800 11088 108031 11488
rect 800 10808 107951 11088
rect 800 10408 108031 10808
rect 880 10128 107951 10408
rect 800 9728 108031 10128
rect 880 9448 107951 9728
rect 800 9048 108031 9448
rect 880 8768 108031 9048
rect 800 8368 108031 8768
rect 880 8088 107951 8368
rect 800 7688 108031 8088
rect 800 7408 107951 7688
rect 800 7008 108031 7408
rect 880 6728 107951 7008
rect 800 6328 108031 6728
rect 880 6048 107951 6328
rect 800 5648 108031 6048
rect 880 5368 108031 5648
rect 800 4968 108031 5368
rect 880 4688 107951 4968
rect 800 4288 108031 4688
rect 800 4008 107951 4288
rect 800 3608 108031 4008
rect 880 3328 107951 3608
rect 800 2928 108031 3328
rect 880 2648 107951 2928
rect 800 2248 108031 2648
rect 880 1968 108031 2248
rect 800 1568 108031 1968
rect 880 1288 107951 1568
rect 800 888 108031 1288
rect 800 715 107951 888
<< metal4 >>
rect -8576 -7504 -7976 117936
rect -7636 -6564 -7036 116996
rect -6696 -5624 -6096 116056
rect -5756 -4684 -5156 115116
rect -4816 -3744 -4216 114176
rect -3876 -2804 -3276 113236
rect -2936 -1864 -2336 112296
rect -1996 -924 -1396 111356
rect 804 -1864 1404 112296
rect 4404 -3744 5004 114176
rect 8004 -5624 8604 116056
rect 11604 -7504 12204 117936
rect 18804 -1864 19404 112296
rect 22404 -3744 23004 114176
rect 26004 -5624 26604 116056
rect 29604 -7504 30204 117936
rect 36804 -1864 37404 112296
rect 40404 -3744 41004 114176
rect 44004 -5624 44604 116056
rect 47604 -7504 48204 117936
rect 54804 -1864 55404 112296
rect 58404 -3744 59004 114176
rect 62004 -5624 62604 116056
rect 65604 -7504 66204 117936
rect 72804 -1864 73404 112296
rect 76404 -3744 77004 114176
rect 80004 -5624 80604 116056
rect 83604 -7504 84204 117936
rect 90804 -1864 91404 112296
rect 94404 -3744 95004 114176
rect 98004 -5624 98604 116056
rect 101604 -7504 102204 117936
rect 110140 -924 110740 111356
rect 111080 -1864 111680 112296
rect 112020 -2804 112620 113236
rect 112960 -3744 113560 114176
rect 113900 -4684 114500 115116
rect 114840 -5624 115440 116056
rect 115780 -6564 116380 116996
rect 116720 -7504 117320 117936
<< obsm4 >>
rect 27843 12955 29524 93397
rect 30284 12955 36724 93397
rect 37484 12955 40324 93397
rect 41084 12955 43924 93397
rect 44684 12955 47524 93397
rect 48284 12955 54724 93397
rect 55484 12955 58324 93397
rect 59084 12955 61924 93397
rect 62684 12955 65524 93397
rect 66284 12955 72724 93397
rect 73484 12955 76324 93397
rect 77084 12955 79924 93397
rect 80684 12955 83524 93397
rect 84284 12955 90724 93397
rect 91484 12955 93781 93397
<< metal5 >>
rect -8576 117336 117320 117936
rect -7636 116396 116380 116996
rect -6696 115456 115440 116056
rect -5756 114516 114500 115116
rect -4816 113576 113560 114176
rect -3876 112636 112620 113236
rect -2936 111696 111680 112296
rect -1996 110756 110740 111356
rect -8576 102676 117320 103276
rect -6696 99076 115440 99676
rect -4816 95476 113560 96076
rect -2936 91828 111680 92428
rect -8576 84676 117320 85276
rect -6696 81076 115440 81676
rect -4816 77476 113560 78076
rect -2936 73828 111680 74428
rect -8576 66676 117320 67276
rect -6696 63076 115440 63676
rect -4816 59476 113560 60076
rect -2936 55828 111680 56428
rect -8576 48676 117320 49276
rect -6696 45076 115440 45676
rect -4816 41476 113560 42076
rect -2936 37828 111680 38428
rect -8576 30676 117320 31276
rect -6696 27076 115440 27676
rect -4816 23476 113560 24076
rect -2936 19828 111680 20428
rect -8576 12676 117320 13276
rect -6696 9076 115440 9676
rect -4816 5476 113560 6076
rect -2936 1828 111680 2428
rect -1996 -924 110740 -324
rect -2936 -1864 111680 -1264
rect -3876 -2804 112620 -2204
rect -4816 -3744 113560 -3144
rect -5756 -4684 114500 -4084
rect -6696 -5624 115440 -5024
rect -7636 -6564 116380 -5964
rect -8576 -7504 117320 -6904
<< obsm5 >>
rect -8576 117936 -7976 117938
rect 29604 117936 30204 117938
rect 65604 117936 66204 117938
rect 101604 117936 102204 117938
rect 116720 117936 117320 117938
rect -8576 117334 -7976 117336
rect 29604 117334 30204 117336
rect 65604 117334 66204 117336
rect 101604 117334 102204 117336
rect 116720 117334 117320 117336
rect -7636 116996 -7036 116998
rect 11604 116996 12204 116998
rect 47604 116996 48204 116998
rect 83604 116996 84204 116998
rect 115780 116996 116380 116998
rect -7636 116394 -7036 116396
rect 11604 116394 12204 116396
rect 47604 116394 48204 116396
rect 83604 116394 84204 116396
rect 115780 116394 116380 116396
rect -6696 116056 -6096 116058
rect 26004 116056 26604 116058
rect 62004 116056 62604 116058
rect 98004 116056 98604 116058
rect 114840 116056 115440 116058
rect -6696 115454 -6096 115456
rect 26004 115454 26604 115456
rect 62004 115454 62604 115456
rect 98004 115454 98604 115456
rect 114840 115454 115440 115456
rect -5756 115116 -5156 115118
rect 8004 115116 8604 115118
rect 44004 115116 44604 115118
rect 80004 115116 80604 115118
rect 113900 115116 114500 115118
rect -5756 114514 -5156 114516
rect 8004 114514 8604 114516
rect 44004 114514 44604 114516
rect 80004 114514 80604 114516
rect 113900 114514 114500 114516
rect -4816 114176 -4216 114178
rect 22404 114176 23004 114178
rect 58404 114176 59004 114178
rect 94404 114176 95004 114178
rect 112960 114176 113560 114178
rect -4816 113574 -4216 113576
rect 22404 113574 23004 113576
rect 58404 113574 59004 113576
rect 94404 113574 95004 113576
rect 112960 113574 113560 113576
rect -3876 113236 -3276 113238
rect 4404 113236 5004 113238
rect 40404 113236 41004 113238
rect 76404 113236 77004 113238
rect 112020 113236 112620 113238
rect -3876 112634 -3276 112636
rect 4404 112634 5004 112636
rect 40404 112634 41004 112636
rect 76404 112634 77004 112636
rect 112020 112634 112620 112636
rect -2936 112296 -2336 112298
rect 18804 112296 19404 112298
rect 54804 112296 55404 112298
rect 90804 112296 91404 112298
rect 111080 112296 111680 112298
rect -2936 111694 -2336 111696
rect 18804 111694 19404 111696
rect 54804 111694 55404 111696
rect 90804 111694 91404 111696
rect 111080 111694 111680 111696
rect -1996 111356 -1396 111358
rect 804 111356 1404 111358
rect 36804 111356 37404 111358
rect 72804 111356 73404 111358
rect 110140 111356 110740 111358
rect -1996 110754 -1396 110756
rect 110140 110754 110740 110756
rect 0 103596 108831 110436
rect -8576 103276 -7976 103278
rect 116720 103276 117320 103278
rect -8576 102674 -7976 102676
rect 116720 102674 117320 102676
rect 0 99996 108831 102356
rect -6696 99676 -6096 99678
rect 114840 99676 115440 99678
rect -6696 99074 -6096 99076
rect 114840 99074 115440 99076
rect 0 96396 108831 98756
rect -4816 96076 -4216 96078
rect 112960 96076 113560 96078
rect -4816 95474 -4216 95476
rect 112960 95474 113560 95476
rect 0 92748 108831 95156
rect -2936 92428 -2336 92430
rect 111080 92428 111680 92430
rect -2936 91826 -2336 91828
rect 111080 91826 111680 91828
rect 0 85596 108831 91508
rect -7636 85276 -7036 85278
rect 115780 85276 116380 85278
rect -7636 84674 -7036 84676
rect 115780 84674 116380 84676
rect 0 81996 108831 84356
rect -5756 81676 -5156 81678
rect 113900 81676 114500 81678
rect -5756 81074 -5156 81076
rect 113900 81074 114500 81076
rect 0 78396 108831 80756
rect -3876 78076 -3276 78078
rect 112020 78076 112620 78078
rect -3876 77474 -3276 77476
rect 112020 77474 112620 77476
rect 0 74748 108831 77156
rect -1996 74428 -1396 74430
rect 110140 74428 110740 74430
rect -1996 73826 -1396 73828
rect 110140 73826 110740 73828
rect 0 67596 108831 73508
rect -8576 67276 -7976 67278
rect 116720 67276 117320 67278
rect -8576 66674 -7976 66676
rect 116720 66674 117320 66676
rect 0 63996 108831 66356
rect -6696 63676 -6096 63678
rect 114840 63676 115440 63678
rect -6696 63074 -6096 63076
rect 114840 63074 115440 63076
rect 0 60396 108831 62756
rect -4816 60076 -4216 60078
rect 112960 60076 113560 60078
rect -4816 59474 -4216 59476
rect 112960 59474 113560 59476
rect 0 56748 108831 59156
rect -2936 56428 -2336 56430
rect 111080 56428 111680 56430
rect -2936 55826 -2336 55828
rect 111080 55826 111680 55828
rect 0 49596 108831 55508
rect -7636 49276 -7036 49278
rect 115780 49276 116380 49278
rect -7636 48674 -7036 48676
rect 115780 48674 116380 48676
rect 0 45996 108831 48356
rect -5756 45676 -5156 45678
rect 113900 45676 114500 45678
rect -5756 45074 -5156 45076
rect 113900 45074 114500 45076
rect 0 42396 108831 44756
rect -3876 42076 -3276 42078
rect 112020 42076 112620 42078
rect -3876 41474 -3276 41476
rect 112020 41474 112620 41476
rect 0 38748 108831 41156
rect -1996 38428 -1396 38430
rect 110140 38428 110740 38430
rect -1996 37826 -1396 37828
rect 110140 37826 110740 37828
rect 0 31596 108831 37508
rect -8576 31276 -7976 31278
rect 116720 31276 117320 31278
rect -8576 30674 -7976 30676
rect 116720 30674 117320 30676
rect 0 27996 108831 30356
rect -6696 27676 -6096 27678
rect 114840 27676 115440 27678
rect -6696 27074 -6096 27076
rect 114840 27074 115440 27076
rect 0 24396 108831 26756
rect -4816 24076 -4216 24078
rect 112960 24076 113560 24078
rect -4816 23474 -4216 23476
rect 112960 23474 113560 23476
rect 0 20748 108831 23156
rect -2936 20428 -2336 20430
rect 111080 20428 111680 20430
rect -2936 19826 -2336 19828
rect 111080 19826 111680 19828
rect 0 13596 108831 19508
rect -7636 13276 -7036 13278
rect 115780 13276 116380 13278
rect -7636 12674 -7036 12676
rect 115780 12674 116380 12676
rect 0 9996 108831 12356
rect -5756 9676 -5156 9678
rect 113900 9676 114500 9678
rect -5756 9074 -5156 9076
rect 113900 9074 114500 9076
rect 0 6396 108831 8756
rect -3876 6076 -3276 6078
rect 112020 6076 112620 6078
rect -3876 5474 -3276 5476
rect 112020 5474 112620 5476
rect 0 2748 108831 5156
rect -1996 2428 -1396 2430
rect 110140 2428 110740 2430
rect -1996 1826 -1396 1828
rect 110140 1826 110740 1828
rect 0 0 108831 1508
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 110140 -324 110740 -322
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 110140 -926 110740 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 111080 -1264 111680 -1262
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 111080 -1866 111680 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112020 -2204 112620 -2202
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112020 -2806 112620 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 112960 -3144 113560 -3142
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 112960 -3746 113560 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 113900 -4084 114500 -4082
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 113900 -4686 114500 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 114840 -5024 115440 -5022
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 114840 -5626 115440 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 115780 -5964 116380 -5962
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 115780 -6566 116380 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 116720 -6904 117320 -6902
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 116720 -7506 117320 -7504
<< labels >>
rlabel metal2 s 2778 110175 2834 110975 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 108031 85688 108831 85808 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 84658 0 84714 800 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal3 s 0 105408 800 105528 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal3 s 108031 87048 108831 87168 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 97078 0 97134 800 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal3 s 0 78888 800 79008 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 5538 0 5594 800 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 74078 0 74134 800 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal2 s 58898 0 58954 800 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 65798 110175 65854 110975 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal2 s 102138 0 102194 800 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 0 1368 800 1488 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal2 s 64418 0 64474 800 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 108031 45568 108831 45688 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 71318 110175 71374 110975 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal2 s 66718 0 66774 800 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal2 s 80978 110175 81034 110975 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal2 s 6458 0 6514 800 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 0 36048 800 36168 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 108031 72088 108831 72208 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 0 47608 800 47728 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 108031 102688 108831 102808 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal2 s 69018 0 69074 800 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 0 106088 800 106208 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal2 s 31298 0 31354 800 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal2 s 51998 0 52054 800 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 87878 110175 87934 110975 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal3 s 108031 57808 108831 57928 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal2 s 98458 0 98514 800 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 io_in[10]
port 31 nsew signal input
rlabel metal2 s 101218 110175 101274 110975 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 io_in[12]
port 33 nsew signal input
rlabel metal2 s 37738 110175 37794 110975 6 io_in[13]
port 34 nsew signal input
rlabel metal2 s 19338 110175 19394 110975 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 io_in[15]
port 36 nsew signal input
rlabel metal3 s 0 70048 800 70168 6 io_in[16]
port 37 nsew signal input
rlabel metal3 s 108031 65288 108831 65408 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 97078 110175 97134 110975 6 io_in[18]
port 39 nsew signal input
rlabel metal3 s 108031 2728 108831 2848 6 io_in[19]
port 40 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 63498 110175 63554 110975 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 66718 110175 66774 110975 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40958 110175 41014 110975 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 io_in[24]
port 46 nsew signal input
rlabel metal3 s 108031 52368 108831 52488 6 io_in[25]
port 47 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 io_in[26]
port 48 nsew signal input
rlabel metal2 s 27618 110175 27674 110975 6 io_in[27]
port 49 nsew signal input
rlabel metal2 s 28538 110175 28594 110975 6 io_in[28]
port 50 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 io_in[29]
port 51 nsew signal input
rlabel metal2 s 90178 110175 90234 110975 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s 108031 10208 108831 10328 6 io_in[30]
port 53 nsew signal input
rlabel metal3 s 108031 6808 108831 6928 6 io_in[31]
port 54 nsew signal input
rlabel metal2 s 8298 110175 8354 110975 6 io_in[32]
port 55 nsew signal input
rlabel metal3 s 0 109488 800 109608 6 io_in[33]
port 56 nsew signal input
rlabel metal3 s 108031 82288 108831 82408 6 io_in[34]
port 57 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 io_in[35]
port 58 nsew signal input
rlabel metal2 s 50618 110175 50674 110975 6 io_in[36]
port 59 nsew signal input
rlabel metal2 s 13818 110175 13874 110975 6 io_in[37]
port 60 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 io_in[3]
port 61 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 108031 18368 108831 18488 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 0 91808 800 91928 6 io_in[6]
port 64 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 io_in[7]
port 65 nsew signal input
rlabel metal2 s 101678 110175 101734 110975 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 108031 97928 108831 98048 6 io_in[9]
port 67 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 io_oeb[0]
port 68 nsew signal output
rlabel metal2 s 100758 0 100814 800 6 io_oeb[10]
port 69 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 io_oeb[11]
port 70 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 io_oeb[12]
port 71 nsew signal output
rlabel metal2 s 35898 110175 35954 110975 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 108031 63248 108831 63368 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 94778 110175 94834 110975 6 io_oeb[15]
port 74 nsew signal output
rlabel metal3 s 108031 25168 108831 25288 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 99378 110175 99434 110975 6 io_oeb[18]
port 77 nsew signal output
rlabel metal3 s 108031 41488 108831 41608 6 io_oeb[19]
port 78 nsew signal output
rlabel metal2 s 80058 0 80114 800 6 io_oeb[1]
port 79 nsew signal output
rlabel metal3 s 108031 66648 108831 66768 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 8758 110175 8814 110975 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 94778 0 94834 800 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s 108031 19728 108831 19848 6 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s 0 104048 800 104168 6 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 io_oeb[26]
port 86 nsew signal output
rlabel metal2 s 48778 110175 48834 110975 6 io_oeb[27]
port 87 nsew signal output
rlabel metal2 s 22098 110175 22154 110975 6 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 io_oeb[29]
port 89 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s 0 83648 800 83768 6 io_oeb[30]
port 91 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 io_oeb[31]
port 92 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s 108031 16328 108831 16448 6 io_oeb[33]
port 94 nsew signal output
rlabel metal2 s 31758 110175 31814 110975 6 io_oeb[34]
port 95 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 io_oeb[36]
port 97 nsew signal output
rlabel metal2 s 14738 110175 14794 110975 6 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 108031 688 108831 808 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 io_oeb[4]
port 100 nsew signal output
rlabel metal2 s 93858 0 93914 800 6 io_oeb[5]
port 101 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 io_oeb[6]
port 102 nsew signal output
rlabel metal2 s 23018 110175 23074 110975 6 io_oeb[7]
port 103 nsew signal output
rlabel metal2 s 68558 0 68614 800 6 io_oeb[8]
port 104 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 io_oeb[9]
port 105 nsew signal output
rlabel metal2 s 49698 110175 49754 110975 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 io_out[10]
port 107 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 108031 68008 108831 68128 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 0 65288 800 65408 6 io_out[13]
port 110 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 95238 110175 95294 110975 6 io_out[15]
port 112 nsew signal output
rlabel metal3 s 108031 106088 108831 106208 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 5998 110175 6054 110975 6 io_out[17]
port 114 nsew signal output
rlabel metal3 s 108031 17008 108831 17128 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 0 95208 800 95328 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 73158 110175 73214 110975 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 47858 110175 47914 110975 6 io_out[21]
port 119 nsew signal output
rlabel metal3 s 0 80248 800 80368 6 io_out[22]
port 120 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s 108031 94528 108831 94648 6 io_out[24]
port 122 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 io_out[25]
port 123 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 io_out[26]
port 124 nsew signal output
rlabel metal2 s 98918 110175 98974 110975 6 io_out[27]
port 125 nsew signal output
rlabel metal2 s 92938 0 92994 800 6 io_out[28]
port 126 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 io_out[29]
port 127 nsew signal output
rlabel metal2 s 76378 0 76434 800 6 io_out[2]
port 128 nsew signal output
rlabel metal2 s 38198 110175 38254 110975 6 io_out[30]
port 129 nsew signal output
rlabel metal3 s 108031 65968 108831 66088 6 io_out[31]
port 130 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 io_out[32]
port 131 nsew signal output
rlabel metal2 s 42338 110175 42394 110975 6 io_out[33]
port 132 nsew signal output
rlabel metal2 s 1858 110175 1914 110975 6 io_out[34]
port 133 nsew signal output
rlabel metal3 s 108031 49648 108831 49768 6 io_out[35]
port 134 nsew signal output
rlabel metal2 s 6918 110175 6974 110975 6 io_out[36]
port 135 nsew signal output
rlabel metal3 s 0 61888 800 62008 6 io_out[37]
port 136 nsew signal output
rlabel metal2 s 105358 110175 105414 110975 6 io_out[3]
port 137 nsew signal output
rlabel metal2 s 85118 110175 85174 110975 6 io_out[4]
port 138 nsew signal output
rlabel metal2 s 103058 110175 103114 110975 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 0 63248 800 63368 6 io_out[6]
port 140 nsew signal output
rlabel metal2 s 96158 110175 96214 110975 6 io_out[7]
port 141 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 io_out[9]
port 143 nsew signal output
rlabel metal3 s 0 90448 800 90568 6 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_data_in[100]
port 145 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 la_data_in[101]
port 146 nsew signal input
rlabel metal3 s 108031 28568 108831 28688 6 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 80058 110175 80114 110975 6 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_data_in[104]
port 149 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 la_data_in[105]
port 150 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 la_data_in[106]
port 151 nsew signal input
rlabel metal3 s 108031 84328 108831 84448 6 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 la_data_in[109]
port 154 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 la_data_in[10]
port 155 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 la_data_in[110]
port 156 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 la_data_in[111]
port 157 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 57978 110175 58034 110975 6 la_data_in[114]
port 160 nsew signal input
rlabel metal3 s 108031 25848 108831 25968 6 la_data_in[115]
port 161 nsew signal input
rlabel metal3 s 108031 69368 108831 69488 6 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 938 0 994 800 6 la_data_in[118]
port 164 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 la_data_in[119]
port 165 nsew signal input
rlabel metal3 s 108031 44208 108831 44328 6 la_data_in[11]
port 166 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 86498 110175 86554 110975 6 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 33138 110175 33194 110975 6 la_data_in[124]
port 171 nsew signal input
rlabel metal3 s 108031 12928 108831 13048 6 la_data_in[125]
port 172 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 11518 110175 11574 110975 6 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 47398 110175 47454 110975 6 la_data_in[12]
port 175 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 la_data_in[13]
port 176 nsew signal input
rlabel metal3 s 108031 106768 108831 106888 6 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 la_data_in[15]
port 178 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 478 110175 534 110975 6 la_data_in[17]
port 180 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 7838 110175 7894 110975 6 la_data_in[19]
port 182 nsew signal input
rlabel metal3 s 108031 46248 108831 46368 6 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 78678 110175 78734 110975 6 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 66258 110175 66314 110975 6 la_data_in[21]
port 185 nsew signal input
rlabel metal3 s 108031 48968 108831 49088 6 la_data_in[22]
port 186 nsew signal input
rlabel metal3 s 108031 100648 108831 100768 6 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 72698 110175 72754 110975 6 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_data_in[27]
port 191 nsew signal input
rlabel metal3 s 108031 21088 108831 21208 6 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 57518 110175 57574 110975 6 la_data_in[2]
port 194 nsew signal input
rlabel metal3 s 108031 37408 108831 37528 6 la_data_in[30]
port 195 nsew signal input
rlabel metal3 s 108031 10888 108831 11008 6 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 20718 110175 20774 110975 6 la_data_in[32]
port 197 nsew signal input
rlabel metal3 s 108031 101328 108831 101448 6 la_data_in[33]
port 198 nsew signal input
rlabel metal3 s 108031 40808 108831 40928 6 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 87418 110175 87474 110975 6 la_data_in[35]
port 200 nsew signal input
rlabel metal3 s 108031 22448 108831 22568 6 la_data_in[36]
port 201 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 la_data_in[37]
port 202 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 104438 110175 104494 110975 6 la_data_in[39]
port 204 nsew signal input
rlabel metal3 s 108031 27888 108831 28008 6 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 92018 110175 92074 110975 6 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 la_data_in[41]
port 207 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 34058 110175 34114 110975 6 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 77298 110175 77354 110975 6 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 54298 110175 54354 110975 6 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 25318 110175 25374 110975 6 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 17958 110175 18014 110975 6 la_data_in[47]
port 213 nsew signal input
rlabel metal3 s 108031 93848 108831 93968 6 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 3698 110175 3754 110975 6 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_data_in[4]
port 216 nsew signal input
rlabel metal3 s 108031 68688 108831 68808 6 la_data_in[50]
port 217 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 50158 110175 50214 110975 6 la_data_in[52]
port 219 nsew signal input
rlabel metal3 s 108031 79568 108831 79688 6 la_data_in[53]
port 220 nsew signal input
rlabel metal3 s 108031 95888 108831 96008 6 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 36358 110175 36414 110975 6 la_data_in[55]
port 222 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 38658 110175 38714 110975 6 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 100758 110175 100814 110975 6 la_data_in[59]
port 226 nsew signal input
rlabel metal3 s 108031 39448 108831 39568 6 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 96618 110175 96674 110975 6 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 53378 110175 53434 110975 6 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 94318 110175 94374 110975 6 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 46018 110175 46074 110975 6 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 55218 110175 55274 110975 6 la_data_in[65]
port 233 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 la_data_in[67]
port 235 nsew signal input
rlabel metal3 s 108031 31968 108831 32088 6 la_data_in[68]
port 236 nsew signal input
rlabel metal3 s 108031 108128 108831 108248 6 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 la_data_in[6]
port 238 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 la_data_in[70]
port 239 nsew signal input
rlabel metal3 s 108031 89088 108831 89208 6 la_data_in[71]
port 240 nsew signal input
rlabel metal3 s 108031 97248 108831 97368 6 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 71778 110175 71834 110975 6 la_data_in[73]
port 242 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 la_data_in[74]
port 243 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 23938 110175 23994 110975 6 la_data_in[78]
port 247 nsew signal input
rlabel metal3 s 108031 56448 108831 56568 6 la_data_in[79]
port 248 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 12438 110175 12494 110975 6 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 92938 110175 92994 110975 6 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 107658 110175 107714 110975 6 la_data_in[84]
port 254 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 60278 110175 60334 110975 6 la_data_in[86]
port 256 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 17498 110175 17554 110975 6 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 58898 110175 58954 110975 6 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_data_in[8]
port 260 nsew signal input
rlabel metal3 s 108031 71408 108831 71528 6 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 81898 110175 81954 110975 6 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 39118 110175 39174 110975 6 la_data_in[93]
port 264 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 78218 110175 78274 110975 6 la_data_in[98]
port 269 nsew signal input
rlabel metal3 s 108031 61208 108831 61328 6 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 91558 110175 91614 110975 6 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 la_data_out[100]
port 273 nsew signal output
rlabel metal3 s 0 46928 800 47048 6 la_data_out[101]
port 274 nsew signal output
rlabel metal3 s 108031 75488 108831 75608 6 la_data_out[102]
port 275 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 61658 110175 61714 110975 6 la_data_out[104]
port 277 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 la_data_out[107]
port 280 nsew signal output
rlabel metal3 s 108031 1368 108831 1488 6 la_data_out[108]
port 281 nsew signal output
rlabel metal3 s 0 91128 800 91248 6 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 32218 110175 32274 110975 6 la_data_out[10]
port 283 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 20258 110175 20314 110975 6 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 86958 110175 87014 110975 6 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 68558 110175 68614 110975 6 la_data_out[114]
port 288 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 la_data_out[115]
port 289 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 28998 110175 29054 110975 6 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 26238 110175 26294 110975 6 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 108118 110175 108174 110975 6 la_data_out[119]
port 293 nsew signal output
rlabel metal3 s 108031 82968 108831 83088 6 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 la_data_out[120]
port 295 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 la_data_out[121]
port 296 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 106278 110175 106334 110975 6 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 104438 0 104494 800 6 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 la_data_out[125]
port 300 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 la_data_out[126]
port 301 nsew signal output
rlabel metal3 s 0 101328 800 101448 6 la_data_out[127]
port 302 nsew signal output
rlabel metal3 s 108031 62568 108831 62688 6 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 96618 0 96674 800 6 la_data_out[13]
port 304 nsew signal output
rlabel metal3 s 108031 48288 108831 48408 6 la_data_out[14]
port 305 nsew signal output
rlabel metal3 s 0 76848 800 76968 6 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 105818 0 105874 800 6 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 36818 110175 36874 110975 6 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 80518 110175 80574 110975 6 la_data_out[21]
port 313 nsew signal output
rlabel metal3 s 108031 80248 108831 80368 6 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 43258 110175 43314 110975 6 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 40038 110175 40094 110975 6 la_data_out[24]
port 316 nsew signal output
rlabel metal3 s 108031 99288 108831 99408 6 la_data_out[25]
port 317 nsew signal output
rlabel metal3 s 108031 7488 108831 7608 6 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 78218 0 78274 800 6 la_data_out[27]
port 319 nsew signal output
rlabel metal3 s 108031 30608 108831 30728 6 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 la_data_out[2]
port 322 nsew signal output
rlabel metal3 s 108031 51008 108831 51128 6 la_data_out[30]
port 323 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 la_data_out[31]
port 324 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 21638 110175 21694 110975 6 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 la_data_out[34]
port 327 nsew signal output
rlabel metal3 s 108031 53048 108831 53168 6 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 105358 0 105414 800 6 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 103978 110175 104034 110975 6 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 la_data_out[39]
port 332 nsew signal output
rlabel metal3 s 0 92488 800 92608 6 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 la_data_out[41]
port 335 nsew signal output
rlabel metal3 s 108031 59168 108831 59288 6 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 la_data_out[45]
port 339 nsew signal output
rlabel metal3 s 108031 24488 108831 24608 6 la_data_out[46]
port 340 nsew signal output
rlabel metal3 s 108031 14968 108831 15088 6 la_data_out[47]
port 341 nsew signal output
rlabel metal3 s 108031 6128 108831 6248 6 la_data_out[48]
port 342 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 la_data_out[49]
port 343 nsew signal output
rlabel metal3 s 108031 64608 108831 64728 6 la_data_out[4]
port 344 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 76378 110175 76434 110975 6 la_data_out[51]
port 346 nsew signal output
rlabel metal3 s 108031 55768 108831 55888 6 la_data_out[52]
port 347 nsew signal output
rlabel metal3 s 108031 107448 108831 107568 6 la_data_out[53]
port 348 nsew signal output
rlabel metal3 s 108031 110168 108831 110288 6 la_data_out[54]
port 349 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 92018 0 92074 800 6 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 47858 0 47914 800 6 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 46938 110175 46994 110975 6 la_data_out[58]
port 353 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 93858 110175 93914 110975 6 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 la_data_out[61]
port 357 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 la_data_out[62]
port 358 nsew signal output
rlabel metal3 s 108031 31288 108831 31408 6 la_data_out[63]
port 359 nsew signal output
rlabel metal3 s 108031 38768 108831 38888 6 la_data_out[64]
port 360 nsew signal output
rlabel metal3 s 108031 17688 108831 17808 6 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 59818 110175 59874 110975 6 la_data_out[66]
port 362 nsew signal output
rlabel metal3 s 108031 21768 108831 21888 6 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 59358 110175 59414 110975 6 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 la_data_out[69]
port 365 nsew signal output
rlabel metal3 s 0 93848 800 93968 6 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 31298 110175 31354 110975 6 la_data_out[70]
port 367 nsew signal output
rlabel metal3 s 108031 99968 108831 100088 6 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 103518 110175 103574 110975 6 la_data_out[72]
port 369 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 la_data_out[73]
port 370 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 35898 0 35954 800 6 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 40038 0 40094 800 6 la_data_out[77]
port 374 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 62578 110175 62634 110975 6 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 105818 110175 105874 110975 6 la_data_out[7]
port 377 nsew signal output
rlabel metal3 s 108031 73448 108831 73568 6 la_data_out[80]
port 378 nsew signal output
rlabel metal3 s 108031 20408 108831 20528 6 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 51998 110175 52054 110975 6 la_data_out[82]
port 380 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 56598 0 56654 800 6 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 89718 0 89774 800 6 la_data_out[85]
port 383 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 la_data_out[86]
port 384 nsew signal output
rlabel metal3 s 108031 42848 108831 42968 6 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 98458 110175 98514 110975 6 la_data_out[88]
port 386 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 75458 110175 75514 110975 6 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 17038 110175 17094 110975 6 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 15198 110175 15254 110975 6 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 74998 110175 75054 110975 6 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 84198 110175 84254 110975 6 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 1398 0 1454 800 6 la_data_out[94]
port 393 nsew signal output
rlabel metal3 s 108031 38088 108831 38208 6 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 34518 110175 34574 110975 6 la_data_out[96]
port 395 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 62118 0 62174 800 6 la_data_out[98]
port 397 nsew signal output
rlabel metal3 s 108031 80928 108831 81048 6 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 la_oenb[100]
port 401 nsew signal input
rlabel metal3 s 108031 4768 108831 4888 6 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 26698 110175 26754 110975 6 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 la_oenb[104]
port 405 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 la_oenb[105]
port 406 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 la_oenb[106]
port 407 nsew signal input
rlabel metal3 s 0 56448 800 56568 6 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 63958 110175 64014 110975 6 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 30838 110175 30894 110975 6 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 41418 110175 41474 110975 6 la_oenb[110]
port 412 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 la_oenb[111]
port 413 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_oenb[113]
port 415 nsew signal input
rlabel metal3 s 108031 104048 108831 104168 6 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 la_oenb[115]
port 417 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 33598 110175 33654 110975 6 la_oenb[117]
port 419 nsew signal input
rlabel metal3 s 108031 90448 108831 90568 6 la_oenb[118]
port 420 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 97538 110175 97594 110975 6 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_oenb[120]
port 423 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 la_oenb[121]
port 424 nsew signal input
rlabel metal3 s 108031 76848 108831 76968 6 la_oenb[122]
port 425 nsew signal input
rlabel metal3 s 108031 11568 108831 11688 6 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 4158 110175 4214 110975 6 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 la_oenb[127]
port 430 nsew signal input
rlabel metal3 s 108031 89768 108831 89888 6 la_oenb[12]
port 431 nsew signal input
rlabel metal3 s 108031 74808 108831 74928 6 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 88338 110175 88394 110975 6 la_oenb[14]
port 433 nsew signal input
rlabel metal3 s 108031 76168 108831 76288 6 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 12898 110175 12954 110975 6 la_oenb[17]
port 436 nsew signal input
rlabel metal3 s 108031 70048 108831 70168 6 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_oenb[19]
port 438 nsew signal input
rlabel metal3 s 0 108808 800 108928 6 la_oenb[1]
port 439 nsew signal input
rlabel metal3 s 108031 58488 108831 58608 6 la_oenb[20]
port 440 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 56598 110175 56654 110975 6 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 40498 110175 40554 110975 6 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 84658 110175 84714 110975 6 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 9218 110175 9274 110975 6 la_oenb[27]
port 447 nsew signal input
rlabel metal3 s 108031 9528 108831 9648 6 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_oenb[29]
port 449 nsew signal input
rlabel metal3 s 108031 59848 108831 59968 6 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 la_oenb[31]
port 452 nsew signal input
rlabel metal3 s 108031 44888 108831 45008 6 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 55678 110175 55734 110975 6 la_oenb[33]
port 454 nsew signal input
rlabel metal3 s 108031 35368 108831 35488 6 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_oenb[37]
port 458 nsew signal input
rlabel metal3 s 108031 96568 108831 96688 6 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 la_oenb[39]
port 460 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 la_oenb[3]
port 461 nsew signal input
rlabel metal3 s 0 75488 800 75608 6 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 67178 110175 67234 110975 6 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_oenb[42]
port 464 nsew signal input
rlabel metal3 s 108031 47608 108831 47728 6 la_oenb[43]
port 465 nsew signal input
rlabel metal3 s 0 97928 800 98048 6 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 la_oenb[45]
port 467 nsew signal input
rlabel metal3 s 108031 42168 108831 42288 6 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 102138 110175 102194 110975 6 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 43718 110175 43774 110975 6 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 478 0 534 800 6 la_oenb[4]
port 472 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 938 110175 994 110975 6 la_oenb[51]
port 474 nsew signal input
rlabel metal3 s 108031 23808 108831 23928 6 la_oenb[52]
port 475 nsew signal input
rlabel metal3 s 108031 54408 108831 54528 6 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_oenb[54]
port 477 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 24858 110175 24914 110975 6 la_oenb[56]
port 479 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 57058 110175 57114 110975 6 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 73618 110175 73674 110975 6 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_oenb[60]
port 484 nsew signal input
rlabel metal3 s 108031 34688 108831 34808 6 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 la_oenb[62]
port 486 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 la_oenb[63]
port 487 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 la_oenb[64]
port 488 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 6458 110175 6514 110975 6 la_oenb[66]
port 490 nsew signal input
rlabel metal3 s 108031 14288 108831 14408 6 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 62118 110175 62174 110975 6 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 77758 110175 77814 110975 6 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 29918 110175 29974 110975 6 la_oenb[71]
port 496 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 48318 110175 48374 110975 6 la_oenb[74]
port 499 nsew signal input
rlabel metal3 s 0 102688 800 102808 6 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 11058 110175 11114 110975 6 la_oenb[76]
port 501 nsew signal input
rlabel metal3 s 108031 4088 108831 4208 6 la_oenb[77]
port 502 nsew signal input
rlabel metal3 s 0 108128 800 108248 6 la_oenb[78]
port 503 nsew signal input
rlabel metal3 s 108031 27208 108831 27328 6 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 la_oenb[7]
port 505 nsew signal input
rlabel metal3 s 108031 92488 108831 92608 6 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 82358 110175 82414 110975 6 la_oenb[81]
port 507 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oenb[83]
port 509 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 la_oenb[84]
port 510 nsew signal input
rlabel metal3 s 108031 51688 108831 51808 6 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 92478 110175 92534 110975 6 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 45558 110175 45614 110975 6 la_oenb[87]
port 513 nsew signal input
rlabel metal3 s 108031 104728 108831 104848 6 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 la_oenb[89]
port 515 nsew signal input
rlabel metal3 s 108031 83648 108831 83768 6 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 69478 110175 69534 110975 6 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 106738 110175 106794 110975 6 la_oenb[93]
port 520 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 la_oenb[94]
port 521 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_oenb[96]
port 523 nsew signal input
rlabel metal3 s 108031 91128 108831 91248 6 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 54758 110175 54814 110975 6 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 90638 110175 90694 110975 6 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 user_clock2
port 528 nsew signal input
rlabel metal2 s 15658 110175 15714 110975 6 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 79598 110175 79654 110975 6 user_irq[2]
port 531 nsew signal output
rlabel metal2 s 52458 110175 52514 110975 6 wb_clk_i
port 532 nsew signal input
rlabel metal3 s 108031 3408 108831 3528 6 wb_rst_i
port 533 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 wbs_ack_o
port 534 nsew signal output
rlabel metal2 s 51078 110175 51134 110975 6 wbs_adr_i[0]
port 535 nsew signal input
rlabel metal3 s 108031 32648 108831 32768 6 wbs_adr_i[10]
port 536 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 wbs_adr_i[11]
port 537 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 wbs_adr_i[12]
port 538 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 wbs_adr_i[13]
port 539 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 wbs_adr_i[14]
port 540 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 wbs_adr_i[15]
port 541 nsew signal input
rlabel metal3 s 108031 86368 108831 86488 6 wbs_adr_i[16]
port 542 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 wbs_adr_i[17]
port 543 nsew signal input
rlabel metal3 s 108031 8168 108831 8288 6 wbs_adr_i[18]
port 544 nsew signal input
rlabel metal2 s 64878 110175 64934 110975 6 wbs_adr_i[19]
port 545 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_adr_i[1]
port 546 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 wbs_adr_i[20]
port 547 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_adr_i[21]
port 548 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 wbs_adr_i[22]
port 549 nsew signal input
rlabel metal2 s 44638 110175 44694 110975 6 wbs_adr_i[23]
port 550 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_adr_i[24]
port 551 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 wbs_adr_i[25]
port 552 nsew signal input
rlabel metal3 s 0 85008 800 85128 6 wbs_adr_i[26]
port 553 nsew signal input
rlabel metal2 s 70398 110175 70454 110975 6 wbs_adr_i[27]
port 554 nsew signal input
rlabel metal2 s 5538 110175 5594 110975 6 wbs_adr_i[28]
port 555 nsew signal input
rlabel metal3 s 108031 109488 108831 109608 6 wbs_adr_i[29]
port 556 nsew signal input
rlabel metal2 s 13358 110175 13414 110975 6 wbs_adr_i[2]
port 557 nsew signal input
rlabel metal2 s 42798 110175 42854 110975 6 wbs_adr_i[30]
port 558 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_adr_i[31]
port 559 nsew signal input
rlabel metal3 s 108031 61888 108831 62008 6 wbs_adr_i[3]
port 560 nsew signal input
rlabel metal2 s 22558 110175 22614 110975 6 wbs_adr_i[4]
port 561 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 wbs_adr_i[5]
port 562 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 wbs_adr_i[6]
port 563 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 wbs_adr_i[7]
port 564 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wbs_adr_i[8]
port 565 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 wbs_adr_i[9]
port 566 nsew signal input
rlabel metal2 s 52918 110175 52974 110975 6 wbs_cyc_i
port 567 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 wbs_dat_i[0]
port 568 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 wbs_dat_i[10]
port 569 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 wbs_dat_i[11]
port 570 nsew signal input
rlabel metal2 s 89258 110175 89314 110975 6 wbs_dat_i[12]
port 571 nsew signal input
rlabel metal3 s 108031 93168 108831 93288 6 wbs_dat_i[13]
port 572 nsew signal input
rlabel metal3 s 108031 34008 108831 34128 6 wbs_dat_i[14]
port 573 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_dat_i[15]
port 574 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 wbs_dat_i[16]
port 575 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 wbs_dat_i[17]
port 576 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 wbs_dat_i[18]
port 577 nsew signal input
rlabel metal2 s 74078 110175 74134 110975 6 wbs_dat_i[19]
port 578 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 wbs_dat_i[1]
port 579 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 wbs_dat_i[20]
port 580 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_i[21]
port 581 nsew signal input
rlabel metal2 s 99838 110175 99894 110975 6 wbs_dat_i[22]
port 582 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 wbs_dat_i[23]
port 583 nsew signal input
rlabel metal2 s 10598 110175 10654 110975 6 wbs_dat_i[24]
port 584 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_i[25]
port 585 nsew signal input
rlabel metal3 s 108031 13608 108831 13728 6 wbs_dat_i[26]
port 586 nsew signal input
rlabel metal3 s 108031 36048 108831 36168 6 wbs_dat_i[27]
port 587 nsew signal input
rlabel metal2 s 35438 110175 35494 110975 6 wbs_dat_i[28]
port 588 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 wbs_dat_i[29]
port 589 nsew signal input
rlabel metal3 s 108031 103368 108831 103488 6 wbs_dat_i[2]
port 590 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wbs_dat_i[30]
port 591 nsew signal input
rlabel metal2 s 27158 110175 27214 110975 6 wbs_dat_i[31]
port 592 nsew signal input
rlabel metal2 s 70858 110175 70914 110975 6 wbs_dat_i[3]
port 593 nsew signal input
rlabel metal3 s 0 95888 800 96008 6 wbs_dat_i[4]
port 594 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_i[5]
port 595 nsew signal input
rlabel metal2 s 85578 110175 85634 110975 6 wbs_dat_i[6]
port 596 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_i[7]
port 597 nsew signal input
rlabel metal2 s 68098 110175 68154 110975 6 wbs_dat_i[8]
port 598 nsew signal input
rlabel metal3 s 0 99288 800 99408 6 wbs_dat_i[9]
port 599 nsew signal input
rlabel metal2 s 3238 110175 3294 110975 6 wbs_dat_o[0]
port 600 nsew signal output
rlabel metal3 s 108031 87728 108831 87848 6 wbs_dat_o[10]
port 601 nsew signal output
rlabel metal2 s 70398 0 70454 800 6 wbs_dat_o[11]
port 602 nsew signal output
rlabel metal2 s 101678 0 101734 800 6 wbs_dat_o[12]
port 603 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_o[13]
port 604 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 wbs_dat_o[14]
port 605 nsew signal output
rlabel metal2 s 103518 0 103574 800 6 wbs_dat_o[15]
port 606 nsew signal output
rlabel metal2 s 83278 110175 83334 110975 6 wbs_dat_o[16]
port 607 nsew signal output
rlabel metal2 s 1398 110175 1454 110975 6 wbs_dat_o[17]
port 608 nsew signal output
rlabel metal3 s 108031 55088 108831 55208 6 wbs_dat_o[18]
port 609 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 wbs_dat_o[19]
port 610 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 wbs_dat_o[1]
port 611 nsew signal output
rlabel metal2 s 45098 110175 45154 110975 6 wbs_dat_o[20]
port 612 nsew signal output
rlabel metal2 s 24398 110175 24454 110975 6 wbs_dat_o[21]
port 613 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 wbs_dat_o[22]
port 614 nsew signal output
rlabel metal2 s 5078 110175 5134 110975 6 wbs_dat_o[23]
port 615 nsew signal output
rlabel metal2 s 69018 110175 69074 110975 6 wbs_dat_o[24]
port 616 nsew signal output
rlabel metal3 s 108031 72768 108831 72888 6 wbs_dat_o[25]
port 617 nsew signal output
rlabel metal2 s 75918 110175 75974 110975 6 wbs_dat_o[26]
port 618 nsew signal output
rlabel metal2 s 89718 110175 89774 110975 6 wbs_dat_o[27]
port 619 nsew signal output
rlabel metal3 s 108031 29248 108831 29368 6 wbs_dat_o[28]
port 620 nsew signal output
rlabel metal2 s 16118 110175 16174 110975 6 wbs_dat_o[29]
port 621 nsew signal output
rlabel metal3 s 0 67328 800 67448 6 wbs_dat_o[2]
port 622 nsew signal output
rlabel metal2 s 82818 110175 82874 110975 6 wbs_dat_o[30]
port 623 nsew signal output
rlabel metal2 s 29458 110175 29514 110975 6 wbs_dat_o[31]
port 624 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 wbs_dat_o[3]
port 625 nsew signal output
rlabel metal2 s 18418 110175 18474 110975 6 wbs_dat_o[4]
port 626 nsew signal output
rlabel metal2 s 64418 110175 64474 110975 6 wbs_dat_o[5]
port 627 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 wbs_dat_o[6]
port 628 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_o[7]
port 629 nsew signal output
rlabel metal3 s 108031 78208 108831 78328 6 wbs_dat_o[8]
port 630 nsew signal output
rlabel metal3 s 108031 78888 108831 79008 6 wbs_dat_o[9]
port 631 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 wbs_sel_i[0]
port 632 nsew signal input
rlabel metal2 s 10138 110175 10194 110975 6 wbs_sel_i[1]
port 633 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 wbs_sel_i[2]
port 634 nsew signal input
rlabel metal2 s 19798 110175 19854 110975 6 wbs_sel_i[3]
port 635 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 wbs_stb_i
port 636 nsew signal input
rlabel metal2 s 61198 110175 61254 110975 6 wbs_we_i
port 637 nsew signal input
rlabel metal4 s 72804 -1864 73404 112296 6 vccd1
port 638 nsew power bidirectional
rlabel metal4 s 36804 -1864 37404 112296 6 vccd1
port 639 nsew power bidirectional
rlabel metal4 s 804 -1864 1404 112296 6 vccd1
port 640 nsew power bidirectional
rlabel metal4 s 110140 -924 110740 111356 6 vccd1
port 641 nsew power bidirectional
rlabel metal4 s -1996 -924 -1396 111356 4 vccd1
port 642 nsew power bidirectional
rlabel metal5 s -1996 110756 110740 111356 6 vccd1
port 643 nsew power bidirectional
rlabel metal5 s -2936 73828 111680 74428 6 vccd1
port 644 nsew power bidirectional
rlabel metal5 s -2936 37828 111680 38428 6 vccd1
port 645 nsew power bidirectional
rlabel metal5 s -2936 1828 111680 2428 6 vccd1
port 646 nsew power bidirectional
rlabel metal5 s -1996 -924 110740 -324 8 vccd1
port 647 nsew power bidirectional
rlabel metal4 s 111080 -1864 111680 112296 6 vssd1
port 648 nsew ground bidirectional
rlabel metal4 s 90804 -1864 91404 112296 6 vssd1
port 649 nsew ground bidirectional
rlabel metal4 s 54804 -1864 55404 112296 6 vssd1
port 650 nsew ground bidirectional
rlabel metal4 s 18804 -1864 19404 112296 6 vssd1
port 651 nsew ground bidirectional
rlabel metal4 s -2936 -1864 -2336 112296 4 vssd1
port 652 nsew ground bidirectional
rlabel metal5 s -2936 111696 111680 112296 6 vssd1
port 653 nsew ground bidirectional
rlabel metal5 s -2936 91828 111680 92428 6 vssd1
port 654 nsew ground bidirectional
rlabel metal5 s -2936 55828 111680 56428 6 vssd1
port 655 nsew ground bidirectional
rlabel metal5 s -2936 19828 111680 20428 6 vssd1
port 656 nsew ground bidirectional
rlabel metal5 s -2936 -1864 111680 -1264 8 vssd1
port 657 nsew ground bidirectional
rlabel metal4 s 76404 -3744 77004 114176 6 vccd2
port 658 nsew power bidirectional
rlabel metal4 s 40404 -3744 41004 114176 6 vccd2
port 659 nsew power bidirectional
rlabel metal4 s 4404 -3744 5004 114176 6 vccd2
port 660 nsew power bidirectional
rlabel metal4 s 112020 -2804 112620 113236 6 vccd2
port 661 nsew power bidirectional
rlabel metal4 s -3876 -2804 -3276 113236 4 vccd2
port 662 nsew power bidirectional
rlabel metal5 s -3876 112636 112620 113236 6 vccd2
port 663 nsew power bidirectional
rlabel metal5 s -4816 77476 113560 78076 6 vccd2
port 664 nsew power bidirectional
rlabel metal5 s -4816 41476 113560 42076 6 vccd2
port 665 nsew power bidirectional
rlabel metal5 s -4816 5476 113560 6076 6 vccd2
port 666 nsew power bidirectional
rlabel metal5 s -3876 -2804 112620 -2204 8 vccd2
port 667 nsew power bidirectional
rlabel metal4 s 112960 -3744 113560 114176 6 vssd2
port 668 nsew ground bidirectional
rlabel metal4 s 94404 -3744 95004 114176 6 vssd2
port 669 nsew ground bidirectional
rlabel metal4 s 58404 -3744 59004 114176 6 vssd2
port 670 nsew ground bidirectional
rlabel metal4 s 22404 -3744 23004 114176 6 vssd2
port 671 nsew ground bidirectional
rlabel metal4 s -4816 -3744 -4216 114176 4 vssd2
port 672 nsew ground bidirectional
rlabel metal5 s -4816 113576 113560 114176 6 vssd2
port 673 nsew ground bidirectional
rlabel metal5 s -4816 95476 113560 96076 6 vssd2
port 674 nsew ground bidirectional
rlabel metal5 s -4816 59476 113560 60076 6 vssd2
port 675 nsew ground bidirectional
rlabel metal5 s -4816 23476 113560 24076 6 vssd2
port 676 nsew ground bidirectional
rlabel metal5 s -4816 -3744 113560 -3144 8 vssd2
port 677 nsew ground bidirectional
rlabel metal4 s 80004 -5624 80604 116056 6 vdda1
port 678 nsew power bidirectional
rlabel metal4 s 44004 -5624 44604 116056 6 vdda1
port 679 nsew power bidirectional
rlabel metal4 s 8004 -5624 8604 116056 6 vdda1
port 680 nsew power bidirectional
rlabel metal4 s 113900 -4684 114500 115116 6 vdda1
port 681 nsew power bidirectional
rlabel metal4 s -5756 -4684 -5156 115116 4 vdda1
port 682 nsew power bidirectional
rlabel metal5 s -5756 114516 114500 115116 6 vdda1
port 683 nsew power bidirectional
rlabel metal5 s -6696 81076 115440 81676 6 vdda1
port 684 nsew power bidirectional
rlabel metal5 s -6696 45076 115440 45676 6 vdda1
port 685 nsew power bidirectional
rlabel metal5 s -6696 9076 115440 9676 6 vdda1
port 686 nsew power bidirectional
rlabel metal5 s -5756 -4684 114500 -4084 8 vdda1
port 687 nsew power bidirectional
rlabel metal4 s 114840 -5624 115440 116056 6 vssa1
port 688 nsew ground bidirectional
rlabel metal4 s 98004 -5624 98604 116056 6 vssa1
port 689 nsew ground bidirectional
rlabel metal4 s 62004 -5624 62604 116056 6 vssa1
port 690 nsew ground bidirectional
rlabel metal4 s 26004 -5624 26604 116056 6 vssa1
port 691 nsew ground bidirectional
rlabel metal4 s -6696 -5624 -6096 116056 4 vssa1
port 692 nsew ground bidirectional
rlabel metal5 s -6696 115456 115440 116056 6 vssa1
port 693 nsew ground bidirectional
rlabel metal5 s -6696 99076 115440 99676 6 vssa1
port 694 nsew ground bidirectional
rlabel metal5 s -6696 63076 115440 63676 6 vssa1
port 695 nsew ground bidirectional
rlabel metal5 s -6696 27076 115440 27676 6 vssa1
port 696 nsew ground bidirectional
rlabel metal5 s -6696 -5624 115440 -5024 8 vssa1
port 697 nsew ground bidirectional
rlabel metal4 s 83604 -7504 84204 117936 6 vdda2
port 698 nsew power bidirectional
rlabel metal4 s 47604 -7504 48204 117936 6 vdda2
port 699 nsew power bidirectional
rlabel metal4 s 11604 -7504 12204 117936 6 vdda2
port 700 nsew power bidirectional
rlabel metal4 s 115780 -6564 116380 116996 6 vdda2
port 701 nsew power bidirectional
rlabel metal4 s -7636 -6564 -7036 116996 4 vdda2
port 702 nsew power bidirectional
rlabel metal5 s -7636 116396 116380 116996 6 vdda2
port 703 nsew power bidirectional
rlabel metal5 s -8576 84676 117320 85276 6 vdda2
port 704 nsew power bidirectional
rlabel metal5 s -8576 48676 117320 49276 6 vdda2
port 705 nsew power bidirectional
rlabel metal5 s -8576 12676 117320 13276 6 vdda2
port 706 nsew power bidirectional
rlabel metal5 s -7636 -6564 116380 -5964 8 vdda2
port 707 nsew power bidirectional
rlabel metal4 s 116720 -7504 117320 117936 6 vssa2
port 708 nsew ground bidirectional
rlabel metal4 s 101604 -7504 102204 117936 6 vssa2
port 709 nsew ground bidirectional
rlabel metal4 s 65604 -7504 66204 117936 6 vssa2
port 710 nsew ground bidirectional
rlabel metal4 s 29604 -7504 30204 117936 6 vssa2
port 711 nsew ground bidirectional
rlabel metal4 s -8576 -7504 -7976 117936 4 vssa2
port 712 nsew ground bidirectional
rlabel metal5 s -8576 117336 117320 117936 6 vssa2
port 713 nsew ground bidirectional
rlabel metal5 s -8576 102676 117320 103276 6 vssa2
port 714 nsew ground bidirectional
rlabel metal5 s -8576 66676 117320 67276 6 vssa2
port 715 nsew ground bidirectional
rlabel metal5 s -8576 30676 117320 31276 6 vssa2
port 716 nsew ground bidirectional
rlabel metal5 s -8576 -7504 117320 -6904 8 vssa2
port 717 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 108831 110975
string LEFview TRUE
string GDS_FILE /project/openlane/user_project_wrapper/runs/user_project_wrapper/results/magic/user_project_wrapper.gds
string GDS_END 25610182
string GDS_START 130
<< end >>

