VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 898.465 BY 909.185 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 905.185 23.370 909.185 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 700.440 898.465 701.040 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.990 0.000 697.270 4.000 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 714.040 898.465 714.640 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 0.000 800.770 4.000 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 905.185 543.170 909.185 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.190 0.000 844.470 4.000 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 370.640 898.465 371.240 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 905.185 591.470 909.185 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 0.000 550.070 4.000 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 905.185 671.970 909.185 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 588.240 898.465 588.840 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 839.840 898.465 840.440 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.190 0.000 568.470 4.000 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.240 4.000 877.840 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 0.000 428.170 4.000 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.890 905.185 727.170 909.185 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 469.240 898.465 469.840 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 0.000 809.970 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 905.185 837.570 909.185 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 905.185 313.170 909.185 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 905.185 161.370 909.185 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 0.000 715.670 4.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 530.440 898.465 531.040 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.790 905.185 803.070 909.185 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 13.640 898.465 14.240 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 0.000 508.670 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 905.185 524.770 909.185 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 905.185 552.370 909.185 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 905.185 340.770 909.185 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 428.440 898.465 429.040 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 905.185 232.670 909.185 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 905.185 237.270 909.185 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.590 905.185 747.870 909.185 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 78.240 898.465 78.840 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 51.040 898.465 51.640 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 905.185 71.670 909.185 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 904.440 4.000 905.040 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 673.240 898.465 673.840 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.390 0.000 876.670 4.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 905.185 421.270 909.185 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 905.185 117.670 909.185 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 146.240 898.465 146.840 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 0.000 487.970 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.890 905.185 842.170 909.185 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 805.840 898.465 806.440 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.990 0.000 536.270 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 0.000 828.370 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.990 0.000 743.270 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 905.185 297.070 909.185 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 516.840 898.465 517.440 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 905.185 784.670 909.185 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 204.040 898.465 204.640 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.490 905.185 823.770 909.185 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 336.640 898.465 337.240 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 0.000 658.170 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 547.440 898.465 548.040 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 905.185 76.270 909.185 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 0.000 782.370 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 153.040 898.465 153.640 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.440 4.000 854.040 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 905.185 407.470 909.185 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 905.185 184.370 909.185 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 125.840 898.465 126.440 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 905.185 264.870 909.185 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 0.000 366.070 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 905.185 122.270 909.185 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.790 0.000 895.070 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 0.000 773.170 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 905.185 193.570 909.185 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 905.185 412.070 909.185 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 554.240 898.465 554.840 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.790 0.000 527.070 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 905.185 789.270 909.185 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 867.040 898.465 867.640 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 905.185 50.970 909.185 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 132.640 898.465 133.240 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 0.000 437.370 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 905.185 605.270 909.185 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 905.185 398.270 909.185 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 775.240 898.465 775.840 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 0.000 389.070 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 0.000 384.470 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.890 905.185 819.170 909.185 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.290 0.000 768.570 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 0.000 540.870 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 0.000 630.570 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 905.185 317.770 909.185 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 540.640 898.465 541.240 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 905.185 349.970 909.185 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 905.185 18.770 909.185 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 404.640 898.465 405.240 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 905.185 62.470 909.185 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 905.185 869.770 909.185 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 905.185 704.170 909.185 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.090 905.185 851.370 909.185 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 905.185 793.870 909.185 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 0.000 814.570 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 0.000 805.370 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 231.240 898.465 231.840 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 905.185 662.770 909.185 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 0.000 545.470 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 693.640 898.465 694.240 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 0.000 706.470 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.890 0.000 819.170 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 905.185 483.370 909.185 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 210.840 898.465 211.440 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 567.840 898.465 568.440 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 357.040 898.465 357.640 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 0.000 205.070 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 905.185 713.370 909.185 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 905.185 274.070 909.185 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 98.640 898.465 99.240 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 905.185 99.270 909.185 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 905.185 391.370 909.185 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 873.840 898.465 874.440 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 905.185 4.970 909.185 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 905.185 67.070 909.185 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 377.440 898.465 378.040 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 905.185 653.570 909.185 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 905.185 547.770 909.185 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 397.840 898.465 398.440 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 826.240 898.465 826.840 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.390 905.185 600.670 909.185 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.790 0.000 711.070 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 0.000 343.070 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 170.040 898.465 170.640 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 905.185 476.470 909.185 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 302.640 898.465 303.240 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 85.040 898.465 85.640 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 905.185 175.170 909.185 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 833.040 898.465 833.640 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 329.840 898.465 330.440 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.290 905.185 722.570 909.185 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 183.640 898.465 184.240 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.890 905.185 865.170 909.185 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 224.440 898.465 225.040 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.390 905.185 761.670 909.185 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 905.185 283.270 909.185 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 905.185 637.470 909.185 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 905.185 448.870 909.185 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 905.185 211.970 909.185 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 905.185 152.170 909.185 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 768.440 898.465 769.040 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 905.185 32.570 909.185 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 561.040 898.465 561.640 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 905.185 416.670 909.185 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 649.440 898.465 650.040 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 785.440 898.465 786.040 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 905.185 301.670 909.185 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 905.185 322.370 909.185 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 0.000 849.070 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.690 905.185 832.970 909.185 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 323.040 898.465 323.640 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 905.185 798.470 909.185 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 905.185 444.270 909.185 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.790 905.185 780.070 909.185 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.490 0.000 501.770 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 905.185 382.170 909.185 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 905.185 458.070 909.185 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.990 0.000 559.270 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 258.440 898.465 259.040 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 887.440 898.465 888.040 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 727.640 898.465 728.240 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 799.040 898.465 799.640 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 905.185 596.070 909.185 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 0.000 582.270 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 905.185 198.170 909.185 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 462.440 898.465 463.040 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 905.185 103.870 909.185 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.590 905.185 770.870 909.185 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.890 905.185 888.170 909.185 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.490 905.185 501.770 909.185 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 905.185 147.570 909.185 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 905.185 487.970 909.185 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 0.000 692.670 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 581.440 898.465 582.040 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 905.185 676.570 909.185 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 905.185 326.970 909.185 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.790 0.000 734.070 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 0.000 885.870 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 905.185 648.970 909.185 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 496.440 898.465 497.040 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 905.185 757.070 909.185 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.790 0.000 688.070 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 0.000 441.970 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 615.440 898.465 616.040 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 905.185 510.970 909.185 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.240 4.000 826.840 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 0.000 625.970 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 0.000 361.470 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 6.840 898.465 7.440 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 751.440 4.000 752.040 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 905.185 269.470 909.185 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 905.185 170.570 909.185 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 0.000 517.870 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 905.185 717.970 909.185 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.190 905.185 568.470 909.185 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.840 4.000 500.440 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 905.185 241.870 909.185 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 905.185 216.570 909.185 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.490 905.185 892.770 909.185 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 680.040 898.465 680.640 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.240 4.000 860.840 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.690 905.185 878.970 909.185 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.590 0.000 862.870 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 0.000 299.370 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.040 4.000 833.640 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 510.040 898.465 510.640 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 0.000 796.170 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 391.040 898.465 391.640 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.790 0.000 872.070 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 905.185 306.270 909.185 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 0.000 621.370 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 905.185 667.370 909.185 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 656.240 898.465 656.840 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 905.185 359.170 909.185 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 905.185 331.570 909.185 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 812.640 898.465 813.240 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 57.840 898.465 58.440 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 244.840 898.465 245.440 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 414.840 898.465 415.440 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 905.185 179.770 909.185 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 435.240 898.465 435.840 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.190 0.000 867.470 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.190 0.000 752.470 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.290 905.185 860.570 909.185 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 0.000 593.770 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 482.840 898.465 483.440 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.490 0.000 823.770 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 197.240 898.465 197.840 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 119.040 898.465 119.640 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 44.240 898.465 44.840 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 523.640 898.465 524.240 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.590 905.185 632.870 909.185 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 455.640 898.465 456.240 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 880.640 898.465 881.240 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 901.040 898.465 901.640 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 0.000 759.370 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 905.185 386.770 909.185 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.190 905.185 775.470 909.185 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.490 0.000 777.770 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 251.640 898.465 252.240 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 316.240 898.465 316.840 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 139.440 898.465 140.040 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 905.185 497.170 909.185 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 176.840 898.465 177.440 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 905.185 492.570 909.185 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 905.185 260.270 909.185 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 819.440 898.465 820.040 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 905.185 855.970 909.185 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 608.640 4.000 609.240 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 905.185 520.170 909.185 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.090 905.185 874.370 909.185 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 601.840 898.465 602.440 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 159.840 898.465 160.440 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 905.185 430.470 909.185 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 0.000 464.970 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.390 0.000 738.670 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 350.240 898.465 350.840 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 905.185 814.570 909.185 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 615.440 4.000 616.040 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.390 905.185 623.670 909.185 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 905.185 140.670 909.185 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 905.185 126.870 909.185 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 905.185 619.070 909.185 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.690 905.185 694.970 909.185 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 309.440 898.465 310.040 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 905.185 287.870 909.185 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 0.000 513.270 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 666.440 898.465 667.040 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 0.000 478.770 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 34.040 898.465 34.640 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 905.185 221.170 909.185 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 905.185 529.370 909.185 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.490 0.000 639.770 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 905.185 255.670 909.185 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 905.185 345.370 909.185 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.990 0.000 720.270 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 853.440 898.465 854.040 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 905.185 278.670 909.185 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 741.240 898.465 741.840 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.390 905.185 807.670 909.185 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.590 0.000 747.870 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 629.040 898.465 629.640 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 91.840 898.465 92.440 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.990 0.000 858.270 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 905.185 37.170 909.185 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 734.440 898.465 735.040 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 608.640 898.465 609.240 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.790 905.185 734.070 909.185 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 622.240 898.465 622.840 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 0.000 356.870 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 905.185 108.470 909.185 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 574.640 898.465 575.240 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 0.000 786.970 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 476.040 898.465 476.640 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 778.640 4.000 779.240 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 905.185 467.270 909.185 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 905.185 336.170 909.185 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 905.185 699.570 909.185 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 0.000 554.670 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 905.185 80.870 909.185 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 71.440 898.465 72.040 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 0.000 667.370 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 489.640 898.465 490.240 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 363.840 898.465 364.440 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 905.185 462.670 909.185 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 285.640 898.465 286.240 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.190 0.000 890.470 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 792.240 898.465 792.840 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 905.185 556.970 909.185 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 384.240 898.465 384.840 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.840 4.000 806.440 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.190 0.000 729.470 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 343.440 898.465 344.040 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.490 905.185 846.770 909.185 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 905.185 363.770 909.185 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 905.185 9.570 909.185 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 190.440 898.465 191.040 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 442.040 898.465 442.640 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 0.000 474.170 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 905.185 207.370 909.185 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 0.000 763.970 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 905.185 471.870 909.185 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 905.185 609.870 909.185 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 0.000 616.770 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 278.840 898.465 279.440 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 905.185 55.570 909.185 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 112.240 898.465 112.840 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 0.000 460.370 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 905.185 515.570 909.185 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.590 0.000 701.870 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 905.185 642.070 909.185 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 905.185 251.070 909.185 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 0.000 674.270 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 905.185 402.870 909.185 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 4.000 847.240 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 905.185 94.670 909.185 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 27.240 898.465 27.840 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.840 4.000 891.440 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 217.640 898.465 218.240 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 0.000 416.670 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 754.840 898.465 755.440 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.890 905.185 681.170 909.185 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.590 0.000 678.870 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 421.640 898.465 422.240 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 905.185 766.270 909.185 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 905.185 377.570 909.185 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 860.240 898.465 860.840 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 686.840 898.465 687.440 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 0.000 412.070 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 905.185 577.670 909.185 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 905.185 883.570 909.185 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 0.000 573.070 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 748.040 898.465 748.640 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 905.185 453.470 909.185 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.190 905.185 752.470 909.185 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 905.185 131.470 909.185 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 905.185 658.170 909.185 ;
    END
  END user_irq[2]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 905.185 435.070 909.185 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 20.440 898.465 21.040 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 0.000 589.170 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 905.185 425.870 909.185 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 265.240 898.465 265.840 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.990 0.000 881.270 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 0.000 492.570 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 707.240 898.465 707.840 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 64.640 898.465 65.240 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 905.185 538.570 909.185 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 0.000 648.970 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 905.185 368.370 909.185 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.690 0.000 832.970 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 905.185 582.270 909.185 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 905.185 46.370 909.185 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 894.240 898.465 894.840 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 905.185 113.070 909.185 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 905.185 354.570 909.185 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 503.240 898.465 503.840 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 905.185 188.970 909.185 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 0.000 683.470 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.290 0.000 791.570 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 905.185 439.670 909.185 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.390 905.185 738.670 909.185 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 761.640 898.465 762.240 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 272.040 898.465 272.640 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.290 0.000 607.570 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 905.185 614.470 909.185 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 905.185 828.370 909.185 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 0.000 635.170 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 905.185 90.070 909.185 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 105.440 898.465 106.040 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 295.840 898.465 296.440 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 905.185 292.470 909.185 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 846.640 898.465 847.240 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 905.185 228.070 909.185 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 905.185 586.870 909.185 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 905.185 708.770 909.185 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 905.185 563.870 909.185 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 819.440 4.000 820.040 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 905.185 27.970 909.185 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 720.840 898.465 721.440 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 0.000 577.670 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.590 0.000 839.870 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 0.000 853.670 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 905.185 690.370 909.185 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 905.185 14.170 909.185 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 448.840 898.465 449.440 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 0.000 469.570 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 905.185 372.970 909.185 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 905.185 202.770 909.185 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 0.000 662.770 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 905.185 41.770 909.185 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 905.185 573.070 909.185 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 595.040 898.465 595.640 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 905.185 628.270 909.185 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.990 905.185 743.270 909.185 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 238.040 898.465 238.640 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 905.185 136.070 909.185 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 905.185 685.770 909.185 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 905.185 246.470 909.185 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 905.185 156.770 909.185 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 905.185 533.970 909.185 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 0.000 398.270 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 635.840 898.465 636.440 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 894.465 642.640 898.465 643.240 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 905.185 85.470 909.185 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 905.185 165.970 909.185 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 0.000 602.970 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 905.185 506.370 909.185 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 724.020 -9.320 727.020 917.800 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 544.020 -9.320 547.020 917.800 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 364.020 -9.320 367.020 917.800 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.020 -9.320 187.020 917.800 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 4.020 -9.320 7.020 917.800 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 905.360 -4.620 908.360 913.100 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 913.100 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -9.980 910.100 908.360 913.100 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 729.140 913.060 732.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 549.140 913.060 552.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 369.140 913.060 372.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 189.140 913.060 192.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 9.140 913.060 12.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -9.980 -4.620 908.360 -1.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 910.060 -9.320 913.060 917.800 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 814.020 -9.320 817.020 917.800 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 634.020 -9.320 637.020 917.800 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 454.020 -9.320 457.020 917.800 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 274.020 -9.320 277.020 917.800 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 94.020 -9.320 97.020 917.800 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 917.800 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 914.800 913.060 917.800 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 819.140 913.060 822.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 639.140 913.060 642.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 459.140 913.060 462.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 279.140 913.060 282.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 99.140 913.060 102.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 -9.320 913.060 -6.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 742.020 -18.720 745.020 927.200 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 562.020 -18.720 565.020 927.200 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 382.020 -18.720 385.020 927.200 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 202.020 -18.720 205.020 927.200 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.020 -18.720 25.020 927.200 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 914.760 -14.020 917.760 922.500 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 922.500 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -19.380 919.500 917.760 922.500 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 747.380 922.460 750.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 567.380 922.460 570.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 387.380 922.460 390.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 207.380 922.460 210.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 27.380 922.460 30.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -19.380 -14.020 917.760 -11.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 919.460 -18.720 922.460 927.200 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 832.020 -18.720 835.020 927.200 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 652.020 -18.720 655.020 927.200 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 472.020 -18.720 475.020 927.200 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 292.020 -18.720 295.020 927.200 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 112.020 -18.720 115.020 927.200 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 927.200 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 924.200 922.460 927.200 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 837.380 922.460 840.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 657.380 922.460 660.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 477.380 922.460 480.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 297.380 922.460 300.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 117.380 922.460 120.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 -18.720 922.460 -15.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 760.020 -28.120 763.020 936.600 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 580.020 -28.120 583.020 936.600 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 400.020 -28.120 403.020 936.600 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 220.020 -28.120 223.020 936.600 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 40.020 -28.120 43.020 936.600 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 924.160 -23.420 927.160 931.900 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 931.900 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -28.780 928.900 927.160 931.900 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 765.380 931.860 768.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 585.380 931.860 588.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 405.380 931.860 408.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 225.380 931.860 228.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 45.380 931.860 48.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -28.780 -23.420 927.160 -20.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 928.860 -28.120 931.860 936.600 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 850.020 -28.120 853.020 936.600 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 670.020 -28.120 673.020 936.600 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 490.020 -28.120 493.020 936.600 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 310.020 -28.120 313.020 936.600 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 130.020 -28.120 133.020 936.600 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 936.600 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 933.600 931.860 936.600 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 855.380 931.860 858.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 675.380 931.860 678.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 495.380 931.860 498.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 315.380 931.860 318.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 135.380 931.860 138.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 -28.120 931.860 -25.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 778.020 -37.520 781.020 946.000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 598.020 -37.520 601.020 946.000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 418.020 -37.520 421.020 946.000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 238.020 -37.520 241.020 946.000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 58.020 -37.520 61.020 946.000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 933.560 -32.820 936.560 941.300 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 941.300 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -38.180 938.300 936.560 941.300 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 783.380 941.260 786.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 603.380 941.260 606.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 423.380 941.260 426.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 243.380 941.260 246.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 63.380 941.260 66.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -38.180 -32.820 936.560 -29.820 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 938.260 -37.520 941.260 946.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 868.020 -37.520 871.020 946.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 688.020 -37.520 691.020 946.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 508.020 -37.520 511.020 946.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 328.020 -37.520 331.020 946.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 148.020 -37.520 151.020 946.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 946.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 943.000 941.260 946.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 873.380 941.260 876.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 693.380 941.260 696.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 513.380 941.260 516.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 333.380 941.260 336.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 153.380 941.260 156.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 -37.520 941.260 -34.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 4.745 8.585 892.255 896.835 ;
      LAYER met1 ;
        RECT 4.685 8.540 895.090 897.840 ;
      LAYER met2 ;
        RECT 5.610 904.905 9.010 905.185 ;
        RECT 9.850 904.905 13.610 905.185 ;
        RECT 14.450 904.905 18.210 905.185 ;
        RECT 19.050 904.905 22.810 905.185 ;
        RECT 23.650 904.905 27.410 905.185 ;
        RECT 28.250 904.905 32.010 905.185 ;
        RECT 32.850 904.905 36.610 905.185 ;
        RECT 37.450 904.905 41.210 905.185 ;
        RECT 42.050 904.905 45.810 905.185 ;
        RECT 46.650 904.905 50.410 905.185 ;
        RECT 51.250 904.905 55.010 905.185 ;
        RECT 55.850 904.905 61.910 905.185 ;
        RECT 62.750 904.905 66.510 905.185 ;
        RECT 67.350 904.905 71.110 905.185 ;
        RECT 71.950 904.905 75.710 905.185 ;
        RECT 76.550 904.905 80.310 905.185 ;
        RECT 81.150 904.905 84.910 905.185 ;
        RECT 85.750 904.905 89.510 905.185 ;
        RECT 90.350 904.905 94.110 905.185 ;
        RECT 94.950 904.905 98.710 905.185 ;
        RECT 99.550 904.905 103.310 905.185 ;
        RECT 104.150 904.905 107.910 905.185 ;
        RECT 108.750 904.905 112.510 905.185 ;
        RECT 113.350 904.905 117.110 905.185 ;
        RECT 117.950 904.905 121.710 905.185 ;
        RECT 122.550 904.905 126.310 905.185 ;
        RECT 127.150 904.905 130.910 905.185 ;
        RECT 131.750 904.905 135.510 905.185 ;
        RECT 136.350 904.905 140.110 905.185 ;
        RECT 140.950 904.905 147.010 905.185 ;
        RECT 147.850 904.905 151.610 905.185 ;
        RECT 152.450 904.905 156.210 905.185 ;
        RECT 157.050 904.905 160.810 905.185 ;
        RECT 161.650 904.905 165.410 905.185 ;
        RECT 166.250 904.905 170.010 905.185 ;
        RECT 170.850 904.905 174.610 905.185 ;
        RECT 175.450 904.905 179.210 905.185 ;
        RECT 180.050 904.905 183.810 905.185 ;
        RECT 184.650 904.905 188.410 905.185 ;
        RECT 189.250 904.905 193.010 905.185 ;
        RECT 193.850 904.905 197.610 905.185 ;
        RECT 198.450 904.905 202.210 905.185 ;
        RECT 203.050 904.905 206.810 905.185 ;
        RECT 207.650 904.905 211.410 905.185 ;
        RECT 212.250 904.905 216.010 905.185 ;
        RECT 216.850 904.905 220.610 905.185 ;
        RECT 221.450 904.905 227.510 905.185 ;
        RECT 228.350 904.905 232.110 905.185 ;
        RECT 232.950 904.905 236.710 905.185 ;
        RECT 237.550 904.905 241.310 905.185 ;
        RECT 242.150 904.905 245.910 905.185 ;
        RECT 246.750 904.905 250.510 905.185 ;
        RECT 251.350 904.905 255.110 905.185 ;
        RECT 255.950 904.905 259.710 905.185 ;
        RECT 260.550 904.905 264.310 905.185 ;
        RECT 265.150 904.905 268.910 905.185 ;
        RECT 269.750 904.905 273.510 905.185 ;
        RECT 274.350 904.905 278.110 905.185 ;
        RECT 278.950 904.905 282.710 905.185 ;
        RECT 283.550 904.905 287.310 905.185 ;
        RECT 288.150 904.905 291.910 905.185 ;
        RECT 292.750 904.905 296.510 905.185 ;
        RECT 297.350 904.905 301.110 905.185 ;
        RECT 301.950 904.905 305.710 905.185 ;
        RECT 306.550 904.905 312.610 905.185 ;
        RECT 313.450 904.905 317.210 905.185 ;
        RECT 318.050 904.905 321.810 905.185 ;
        RECT 322.650 904.905 326.410 905.185 ;
        RECT 327.250 904.905 331.010 905.185 ;
        RECT 331.850 904.905 335.610 905.185 ;
        RECT 336.450 904.905 340.210 905.185 ;
        RECT 341.050 904.905 344.810 905.185 ;
        RECT 345.650 904.905 349.410 905.185 ;
        RECT 350.250 904.905 354.010 905.185 ;
        RECT 354.850 904.905 358.610 905.185 ;
        RECT 359.450 904.905 363.210 905.185 ;
        RECT 364.050 904.905 367.810 905.185 ;
        RECT 368.650 904.905 372.410 905.185 ;
        RECT 373.250 904.905 377.010 905.185 ;
        RECT 377.850 904.905 381.610 905.185 ;
        RECT 382.450 904.905 386.210 905.185 ;
        RECT 387.050 904.905 390.810 905.185 ;
        RECT 391.650 904.905 397.710 905.185 ;
        RECT 398.550 904.905 402.310 905.185 ;
        RECT 403.150 904.905 406.910 905.185 ;
        RECT 407.750 904.905 411.510 905.185 ;
        RECT 412.350 904.905 416.110 905.185 ;
        RECT 416.950 904.905 420.710 905.185 ;
        RECT 421.550 904.905 425.310 905.185 ;
        RECT 426.150 904.905 429.910 905.185 ;
        RECT 430.750 904.905 434.510 905.185 ;
        RECT 435.350 904.905 439.110 905.185 ;
        RECT 439.950 904.905 443.710 905.185 ;
        RECT 444.550 904.905 448.310 905.185 ;
        RECT 449.150 904.905 452.910 905.185 ;
        RECT 453.750 904.905 457.510 905.185 ;
        RECT 458.350 904.905 462.110 905.185 ;
        RECT 462.950 904.905 466.710 905.185 ;
        RECT 467.550 904.905 471.310 905.185 ;
        RECT 472.150 904.905 475.910 905.185 ;
        RECT 476.750 904.905 482.810 905.185 ;
        RECT 483.650 904.905 487.410 905.185 ;
        RECT 488.250 904.905 492.010 905.185 ;
        RECT 492.850 904.905 496.610 905.185 ;
        RECT 497.450 904.905 501.210 905.185 ;
        RECT 502.050 904.905 505.810 905.185 ;
        RECT 506.650 904.905 510.410 905.185 ;
        RECT 511.250 904.905 515.010 905.185 ;
        RECT 515.850 904.905 519.610 905.185 ;
        RECT 520.450 904.905 524.210 905.185 ;
        RECT 525.050 904.905 528.810 905.185 ;
        RECT 529.650 904.905 533.410 905.185 ;
        RECT 534.250 904.905 538.010 905.185 ;
        RECT 538.850 904.905 542.610 905.185 ;
        RECT 543.450 904.905 547.210 905.185 ;
        RECT 548.050 904.905 551.810 905.185 ;
        RECT 552.650 904.905 556.410 905.185 ;
        RECT 557.250 904.905 563.310 905.185 ;
        RECT 564.150 904.905 567.910 905.185 ;
        RECT 568.750 904.905 572.510 905.185 ;
        RECT 573.350 904.905 577.110 905.185 ;
        RECT 577.950 904.905 581.710 905.185 ;
        RECT 582.550 904.905 586.310 905.185 ;
        RECT 587.150 904.905 590.910 905.185 ;
        RECT 591.750 904.905 595.510 905.185 ;
        RECT 596.350 904.905 600.110 905.185 ;
        RECT 600.950 904.905 604.710 905.185 ;
        RECT 605.550 904.905 609.310 905.185 ;
        RECT 610.150 904.905 613.910 905.185 ;
        RECT 614.750 904.905 618.510 905.185 ;
        RECT 619.350 904.905 623.110 905.185 ;
        RECT 623.950 904.905 627.710 905.185 ;
        RECT 628.550 904.905 632.310 905.185 ;
        RECT 633.150 904.905 636.910 905.185 ;
        RECT 637.750 904.905 641.510 905.185 ;
        RECT 642.350 904.905 648.410 905.185 ;
        RECT 649.250 904.905 653.010 905.185 ;
        RECT 653.850 904.905 657.610 905.185 ;
        RECT 658.450 904.905 662.210 905.185 ;
        RECT 663.050 904.905 666.810 905.185 ;
        RECT 667.650 904.905 671.410 905.185 ;
        RECT 672.250 904.905 676.010 905.185 ;
        RECT 676.850 904.905 680.610 905.185 ;
        RECT 681.450 904.905 685.210 905.185 ;
        RECT 686.050 904.905 689.810 905.185 ;
        RECT 690.650 904.905 694.410 905.185 ;
        RECT 695.250 904.905 699.010 905.185 ;
        RECT 699.850 904.905 703.610 905.185 ;
        RECT 704.450 904.905 708.210 905.185 ;
        RECT 709.050 904.905 712.810 905.185 ;
        RECT 713.650 904.905 717.410 905.185 ;
        RECT 718.250 904.905 722.010 905.185 ;
        RECT 722.850 904.905 726.610 905.185 ;
        RECT 727.450 904.905 733.510 905.185 ;
        RECT 734.350 904.905 738.110 905.185 ;
        RECT 738.950 904.905 742.710 905.185 ;
        RECT 743.550 904.905 747.310 905.185 ;
        RECT 748.150 904.905 751.910 905.185 ;
        RECT 752.750 904.905 756.510 905.185 ;
        RECT 757.350 904.905 761.110 905.185 ;
        RECT 761.950 904.905 765.710 905.185 ;
        RECT 766.550 904.905 770.310 905.185 ;
        RECT 771.150 904.905 774.910 905.185 ;
        RECT 775.750 904.905 779.510 905.185 ;
        RECT 780.350 904.905 784.110 905.185 ;
        RECT 784.950 904.905 788.710 905.185 ;
        RECT 789.550 904.905 793.310 905.185 ;
        RECT 794.150 904.905 797.910 905.185 ;
        RECT 798.750 904.905 802.510 905.185 ;
        RECT 803.350 904.905 807.110 905.185 ;
        RECT 807.950 904.905 814.010 905.185 ;
        RECT 814.850 904.905 818.610 905.185 ;
        RECT 819.450 904.905 823.210 905.185 ;
        RECT 824.050 904.905 827.810 905.185 ;
        RECT 828.650 904.905 832.410 905.185 ;
        RECT 833.250 904.905 837.010 905.185 ;
        RECT 837.850 904.905 841.610 905.185 ;
        RECT 842.450 904.905 846.210 905.185 ;
        RECT 847.050 904.905 850.810 905.185 ;
        RECT 851.650 904.905 855.410 905.185 ;
        RECT 856.250 904.905 860.010 905.185 ;
        RECT 860.850 904.905 864.610 905.185 ;
        RECT 865.450 904.905 869.210 905.185 ;
        RECT 870.050 904.905 873.810 905.185 ;
        RECT 874.650 904.905 878.410 905.185 ;
        RECT 879.250 904.905 883.010 905.185 ;
        RECT 883.850 904.905 887.610 905.185 ;
        RECT 888.450 904.905 892.210 905.185 ;
        RECT 893.050 904.905 895.060 905.185 ;
        RECT 5.610 4.280 895.060 904.905 ;
        RECT 5.610 4.000 6.710 4.280 ;
        RECT 7.550 4.000 11.310 4.280 ;
        RECT 12.150 4.000 15.910 4.280 ;
        RECT 16.750 4.000 20.510 4.280 ;
        RECT 21.350 4.000 25.110 4.280 ;
        RECT 25.950 4.000 29.710 4.280 ;
        RECT 30.550 4.000 34.310 4.280 ;
        RECT 35.150 4.000 38.910 4.280 ;
        RECT 39.750 4.000 43.510 4.280 ;
        RECT 44.350 4.000 48.110 4.280 ;
        RECT 48.950 4.000 52.710 4.280 ;
        RECT 53.550 4.000 57.310 4.280 ;
        RECT 58.150 4.000 61.910 4.280 ;
        RECT 62.750 4.000 66.510 4.280 ;
        RECT 67.350 4.000 71.110 4.280 ;
        RECT 71.950 4.000 75.710 4.280 ;
        RECT 76.550 4.000 80.310 4.280 ;
        RECT 81.150 4.000 87.210 4.280 ;
        RECT 88.050 4.000 91.810 4.280 ;
        RECT 92.650 4.000 96.410 4.280 ;
        RECT 97.250 4.000 101.010 4.280 ;
        RECT 101.850 4.000 105.610 4.280 ;
        RECT 106.450 4.000 110.210 4.280 ;
        RECT 111.050 4.000 114.810 4.280 ;
        RECT 115.650 4.000 119.410 4.280 ;
        RECT 120.250 4.000 124.010 4.280 ;
        RECT 124.850 4.000 128.610 4.280 ;
        RECT 129.450 4.000 133.210 4.280 ;
        RECT 134.050 4.000 137.810 4.280 ;
        RECT 138.650 4.000 142.410 4.280 ;
        RECT 143.250 4.000 147.010 4.280 ;
        RECT 147.850 4.000 151.610 4.280 ;
        RECT 152.450 4.000 156.210 4.280 ;
        RECT 157.050 4.000 160.810 4.280 ;
        RECT 161.650 4.000 165.410 4.280 ;
        RECT 166.250 4.000 172.310 4.280 ;
        RECT 173.150 4.000 176.910 4.280 ;
        RECT 177.750 4.000 181.510 4.280 ;
        RECT 182.350 4.000 186.110 4.280 ;
        RECT 186.950 4.000 190.710 4.280 ;
        RECT 191.550 4.000 195.310 4.280 ;
        RECT 196.150 4.000 199.910 4.280 ;
        RECT 200.750 4.000 204.510 4.280 ;
        RECT 205.350 4.000 209.110 4.280 ;
        RECT 209.950 4.000 213.710 4.280 ;
        RECT 214.550 4.000 218.310 4.280 ;
        RECT 219.150 4.000 222.910 4.280 ;
        RECT 223.750 4.000 227.510 4.280 ;
        RECT 228.350 4.000 232.110 4.280 ;
        RECT 232.950 4.000 236.710 4.280 ;
        RECT 237.550 4.000 241.310 4.280 ;
        RECT 242.150 4.000 245.910 4.280 ;
        RECT 246.750 4.000 250.510 4.280 ;
        RECT 251.350 4.000 257.410 4.280 ;
        RECT 258.250 4.000 262.010 4.280 ;
        RECT 262.850 4.000 266.610 4.280 ;
        RECT 267.450 4.000 271.210 4.280 ;
        RECT 272.050 4.000 275.810 4.280 ;
        RECT 276.650 4.000 280.410 4.280 ;
        RECT 281.250 4.000 285.010 4.280 ;
        RECT 285.850 4.000 289.610 4.280 ;
        RECT 290.450 4.000 294.210 4.280 ;
        RECT 295.050 4.000 298.810 4.280 ;
        RECT 299.650 4.000 303.410 4.280 ;
        RECT 304.250 4.000 308.010 4.280 ;
        RECT 308.850 4.000 312.610 4.280 ;
        RECT 313.450 4.000 317.210 4.280 ;
        RECT 318.050 4.000 321.810 4.280 ;
        RECT 322.650 4.000 326.410 4.280 ;
        RECT 327.250 4.000 331.010 4.280 ;
        RECT 331.850 4.000 337.910 4.280 ;
        RECT 338.750 4.000 342.510 4.280 ;
        RECT 343.350 4.000 347.110 4.280 ;
        RECT 347.950 4.000 351.710 4.280 ;
        RECT 352.550 4.000 356.310 4.280 ;
        RECT 357.150 4.000 360.910 4.280 ;
        RECT 361.750 4.000 365.510 4.280 ;
        RECT 366.350 4.000 370.110 4.280 ;
        RECT 370.950 4.000 374.710 4.280 ;
        RECT 375.550 4.000 379.310 4.280 ;
        RECT 380.150 4.000 383.910 4.280 ;
        RECT 384.750 4.000 388.510 4.280 ;
        RECT 389.350 4.000 393.110 4.280 ;
        RECT 393.950 4.000 397.710 4.280 ;
        RECT 398.550 4.000 402.310 4.280 ;
        RECT 403.150 4.000 406.910 4.280 ;
        RECT 407.750 4.000 411.510 4.280 ;
        RECT 412.350 4.000 416.110 4.280 ;
        RECT 416.950 4.000 423.010 4.280 ;
        RECT 423.850 4.000 427.610 4.280 ;
        RECT 428.450 4.000 432.210 4.280 ;
        RECT 433.050 4.000 436.810 4.280 ;
        RECT 437.650 4.000 441.410 4.280 ;
        RECT 442.250 4.000 446.010 4.280 ;
        RECT 446.850 4.000 450.610 4.280 ;
        RECT 451.450 4.000 455.210 4.280 ;
        RECT 456.050 4.000 459.810 4.280 ;
        RECT 460.650 4.000 464.410 4.280 ;
        RECT 465.250 4.000 469.010 4.280 ;
        RECT 469.850 4.000 473.610 4.280 ;
        RECT 474.450 4.000 478.210 4.280 ;
        RECT 479.050 4.000 482.810 4.280 ;
        RECT 483.650 4.000 487.410 4.280 ;
        RECT 488.250 4.000 492.010 4.280 ;
        RECT 492.850 4.000 496.610 4.280 ;
        RECT 497.450 4.000 501.210 4.280 ;
        RECT 502.050 4.000 508.110 4.280 ;
        RECT 508.950 4.000 512.710 4.280 ;
        RECT 513.550 4.000 517.310 4.280 ;
        RECT 518.150 4.000 521.910 4.280 ;
        RECT 522.750 4.000 526.510 4.280 ;
        RECT 527.350 4.000 531.110 4.280 ;
        RECT 531.950 4.000 535.710 4.280 ;
        RECT 536.550 4.000 540.310 4.280 ;
        RECT 541.150 4.000 544.910 4.280 ;
        RECT 545.750 4.000 549.510 4.280 ;
        RECT 550.350 4.000 554.110 4.280 ;
        RECT 554.950 4.000 558.710 4.280 ;
        RECT 559.550 4.000 563.310 4.280 ;
        RECT 564.150 4.000 567.910 4.280 ;
        RECT 568.750 4.000 572.510 4.280 ;
        RECT 573.350 4.000 577.110 4.280 ;
        RECT 577.950 4.000 581.710 4.280 ;
        RECT 582.550 4.000 588.610 4.280 ;
        RECT 589.450 4.000 593.210 4.280 ;
        RECT 594.050 4.000 597.810 4.280 ;
        RECT 598.650 4.000 602.410 4.280 ;
        RECT 603.250 4.000 607.010 4.280 ;
        RECT 607.850 4.000 611.610 4.280 ;
        RECT 612.450 4.000 616.210 4.280 ;
        RECT 617.050 4.000 620.810 4.280 ;
        RECT 621.650 4.000 625.410 4.280 ;
        RECT 626.250 4.000 630.010 4.280 ;
        RECT 630.850 4.000 634.610 4.280 ;
        RECT 635.450 4.000 639.210 4.280 ;
        RECT 640.050 4.000 643.810 4.280 ;
        RECT 644.650 4.000 648.410 4.280 ;
        RECT 649.250 4.000 653.010 4.280 ;
        RECT 653.850 4.000 657.610 4.280 ;
        RECT 658.450 4.000 662.210 4.280 ;
        RECT 663.050 4.000 666.810 4.280 ;
        RECT 667.650 4.000 673.710 4.280 ;
        RECT 674.550 4.000 678.310 4.280 ;
        RECT 679.150 4.000 682.910 4.280 ;
        RECT 683.750 4.000 687.510 4.280 ;
        RECT 688.350 4.000 692.110 4.280 ;
        RECT 692.950 4.000 696.710 4.280 ;
        RECT 697.550 4.000 701.310 4.280 ;
        RECT 702.150 4.000 705.910 4.280 ;
        RECT 706.750 4.000 710.510 4.280 ;
        RECT 711.350 4.000 715.110 4.280 ;
        RECT 715.950 4.000 719.710 4.280 ;
        RECT 720.550 4.000 724.310 4.280 ;
        RECT 725.150 4.000 728.910 4.280 ;
        RECT 729.750 4.000 733.510 4.280 ;
        RECT 734.350 4.000 738.110 4.280 ;
        RECT 738.950 4.000 742.710 4.280 ;
        RECT 743.550 4.000 747.310 4.280 ;
        RECT 748.150 4.000 751.910 4.280 ;
        RECT 752.750 4.000 758.810 4.280 ;
        RECT 759.650 4.000 763.410 4.280 ;
        RECT 764.250 4.000 768.010 4.280 ;
        RECT 768.850 4.000 772.610 4.280 ;
        RECT 773.450 4.000 777.210 4.280 ;
        RECT 778.050 4.000 781.810 4.280 ;
        RECT 782.650 4.000 786.410 4.280 ;
        RECT 787.250 4.000 791.010 4.280 ;
        RECT 791.850 4.000 795.610 4.280 ;
        RECT 796.450 4.000 800.210 4.280 ;
        RECT 801.050 4.000 804.810 4.280 ;
        RECT 805.650 4.000 809.410 4.280 ;
        RECT 810.250 4.000 814.010 4.280 ;
        RECT 814.850 4.000 818.610 4.280 ;
        RECT 819.450 4.000 823.210 4.280 ;
        RECT 824.050 4.000 827.810 4.280 ;
        RECT 828.650 4.000 832.410 4.280 ;
        RECT 833.250 4.000 839.310 4.280 ;
        RECT 840.150 4.000 843.910 4.280 ;
        RECT 844.750 4.000 848.510 4.280 ;
        RECT 849.350 4.000 853.110 4.280 ;
        RECT 853.950 4.000 857.710 4.280 ;
        RECT 858.550 4.000 862.310 4.280 ;
        RECT 863.150 4.000 866.910 4.280 ;
        RECT 867.750 4.000 871.510 4.280 ;
        RECT 872.350 4.000 876.110 4.280 ;
        RECT 876.950 4.000 880.710 4.280 ;
        RECT 881.550 4.000 885.310 4.280 ;
        RECT 886.150 4.000 889.910 4.280 ;
        RECT 890.750 4.000 894.510 4.280 ;
      LAYER met3 ;
        RECT 4.000 900.640 894.065 901.505 ;
        RECT 4.000 898.640 894.465 900.640 ;
        RECT 4.400 897.240 894.465 898.640 ;
        RECT 4.000 895.240 894.465 897.240 ;
        RECT 4.000 893.840 894.065 895.240 ;
        RECT 4.000 891.840 894.465 893.840 ;
        RECT 4.400 890.440 894.465 891.840 ;
        RECT 4.000 888.440 894.465 890.440 ;
        RECT 4.000 887.040 894.065 888.440 ;
        RECT 4.000 885.040 894.465 887.040 ;
        RECT 4.400 883.640 894.465 885.040 ;
        RECT 4.000 881.640 894.465 883.640 ;
        RECT 4.000 880.240 894.065 881.640 ;
        RECT 4.000 878.240 894.465 880.240 ;
        RECT 4.400 876.840 894.465 878.240 ;
        RECT 4.000 874.840 894.465 876.840 ;
        RECT 4.000 873.440 894.065 874.840 ;
        RECT 4.000 871.440 894.465 873.440 ;
        RECT 4.400 870.040 894.465 871.440 ;
        RECT 4.000 868.040 894.465 870.040 ;
        RECT 4.000 866.640 894.065 868.040 ;
        RECT 4.000 861.240 894.465 866.640 ;
        RECT 4.400 859.840 894.065 861.240 ;
        RECT 4.000 854.440 894.465 859.840 ;
        RECT 4.400 853.040 894.065 854.440 ;
        RECT 4.000 847.640 894.465 853.040 ;
        RECT 4.400 846.240 894.065 847.640 ;
        RECT 4.000 840.840 894.465 846.240 ;
        RECT 4.400 839.440 894.065 840.840 ;
        RECT 4.000 834.040 894.465 839.440 ;
        RECT 4.400 832.640 894.065 834.040 ;
        RECT 4.000 827.240 894.465 832.640 ;
        RECT 4.400 825.840 894.065 827.240 ;
        RECT 4.000 820.440 894.465 825.840 ;
        RECT 4.400 819.040 894.065 820.440 ;
        RECT 4.000 813.640 894.465 819.040 ;
        RECT 4.400 812.240 894.065 813.640 ;
        RECT 4.000 806.840 894.465 812.240 ;
        RECT 4.400 805.440 894.065 806.840 ;
        RECT 4.000 800.040 894.465 805.440 ;
        RECT 4.400 798.640 894.065 800.040 ;
        RECT 4.000 793.240 894.465 798.640 ;
        RECT 4.400 791.840 894.065 793.240 ;
        RECT 4.000 786.440 894.465 791.840 ;
        RECT 4.400 785.040 894.065 786.440 ;
        RECT 4.000 779.640 894.465 785.040 ;
        RECT 4.400 778.240 894.465 779.640 ;
        RECT 4.000 776.240 894.465 778.240 ;
        RECT 4.000 774.840 894.065 776.240 ;
        RECT 4.000 772.840 894.465 774.840 ;
        RECT 4.400 771.440 894.465 772.840 ;
        RECT 4.000 769.440 894.465 771.440 ;
        RECT 4.000 768.040 894.065 769.440 ;
        RECT 4.000 766.040 894.465 768.040 ;
        RECT 4.400 764.640 894.465 766.040 ;
        RECT 4.000 762.640 894.465 764.640 ;
        RECT 4.000 761.240 894.065 762.640 ;
        RECT 4.000 759.240 894.465 761.240 ;
        RECT 4.400 757.840 894.465 759.240 ;
        RECT 4.000 755.840 894.465 757.840 ;
        RECT 4.000 754.440 894.065 755.840 ;
        RECT 4.000 752.440 894.465 754.440 ;
        RECT 4.400 751.040 894.465 752.440 ;
        RECT 4.000 749.040 894.465 751.040 ;
        RECT 4.000 747.640 894.065 749.040 ;
        RECT 4.000 742.240 894.465 747.640 ;
        RECT 4.400 740.840 894.065 742.240 ;
        RECT 4.000 735.440 894.465 740.840 ;
        RECT 4.400 734.040 894.065 735.440 ;
        RECT 4.000 728.640 894.465 734.040 ;
        RECT 4.400 727.240 894.065 728.640 ;
        RECT 4.000 721.840 894.465 727.240 ;
        RECT 4.400 720.440 894.065 721.840 ;
        RECT 4.000 715.040 894.465 720.440 ;
        RECT 4.400 713.640 894.065 715.040 ;
        RECT 4.000 708.240 894.465 713.640 ;
        RECT 4.400 706.840 894.065 708.240 ;
        RECT 4.000 701.440 894.465 706.840 ;
        RECT 4.400 700.040 894.065 701.440 ;
        RECT 4.000 694.640 894.465 700.040 ;
        RECT 4.400 693.240 894.065 694.640 ;
        RECT 4.000 687.840 894.465 693.240 ;
        RECT 4.400 686.440 894.065 687.840 ;
        RECT 4.000 681.040 894.465 686.440 ;
        RECT 4.400 679.640 894.065 681.040 ;
        RECT 4.000 674.240 894.465 679.640 ;
        RECT 4.400 672.840 894.065 674.240 ;
        RECT 4.000 667.440 894.465 672.840 ;
        RECT 4.400 666.040 894.065 667.440 ;
        RECT 4.000 660.640 894.465 666.040 ;
        RECT 4.400 659.240 894.465 660.640 ;
        RECT 4.000 657.240 894.465 659.240 ;
        RECT 4.000 655.840 894.065 657.240 ;
        RECT 4.000 653.840 894.465 655.840 ;
        RECT 4.400 652.440 894.465 653.840 ;
        RECT 4.000 650.440 894.465 652.440 ;
        RECT 4.000 649.040 894.065 650.440 ;
        RECT 4.000 647.040 894.465 649.040 ;
        RECT 4.400 645.640 894.465 647.040 ;
        RECT 4.000 643.640 894.465 645.640 ;
        RECT 4.000 642.240 894.065 643.640 ;
        RECT 4.000 640.240 894.465 642.240 ;
        RECT 4.400 638.840 894.465 640.240 ;
        RECT 4.000 636.840 894.465 638.840 ;
        RECT 4.000 635.440 894.065 636.840 ;
        RECT 4.000 633.440 894.465 635.440 ;
        RECT 4.400 632.040 894.465 633.440 ;
        RECT 4.000 630.040 894.465 632.040 ;
        RECT 4.000 628.640 894.065 630.040 ;
        RECT 4.000 626.640 894.465 628.640 ;
        RECT 4.400 625.240 894.465 626.640 ;
        RECT 4.000 623.240 894.465 625.240 ;
        RECT 4.000 621.840 894.065 623.240 ;
        RECT 4.000 616.440 894.465 621.840 ;
        RECT 4.400 615.040 894.065 616.440 ;
        RECT 4.000 609.640 894.465 615.040 ;
        RECT 4.400 608.240 894.065 609.640 ;
        RECT 4.000 602.840 894.465 608.240 ;
        RECT 4.400 601.440 894.065 602.840 ;
        RECT 4.000 596.040 894.465 601.440 ;
        RECT 4.400 594.640 894.065 596.040 ;
        RECT 4.000 589.240 894.465 594.640 ;
        RECT 4.400 587.840 894.065 589.240 ;
        RECT 4.000 582.440 894.465 587.840 ;
        RECT 4.400 581.040 894.065 582.440 ;
        RECT 4.000 575.640 894.465 581.040 ;
        RECT 4.400 574.240 894.065 575.640 ;
        RECT 4.000 568.840 894.465 574.240 ;
        RECT 4.400 567.440 894.065 568.840 ;
        RECT 4.000 562.040 894.465 567.440 ;
        RECT 4.400 560.640 894.065 562.040 ;
        RECT 4.000 555.240 894.465 560.640 ;
        RECT 4.400 553.840 894.065 555.240 ;
        RECT 4.000 548.440 894.465 553.840 ;
        RECT 4.400 547.040 894.065 548.440 ;
        RECT 4.000 541.640 894.465 547.040 ;
        RECT 4.400 540.240 894.065 541.640 ;
        RECT 4.000 534.840 894.465 540.240 ;
        RECT 4.400 533.440 894.465 534.840 ;
        RECT 4.000 531.440 894.465 533.440 ;
        RECT 4.000 530.040 894.065 531.440 ;
        RECT 4.000 528.040 894.465 530.040 ;
        RECT 4.400 526.640 894.465 528.040 ;
        RECT 4.000 524.640 894.465 526.640 ;
        RECT 4.000 523.240 894.065 524.640 ;
        RECT 4.000 521.240 894.465 523.240 ;
        RECT 4.400 519.840 894.465 521.240 ;
        RECT 4.000 517.840 894.465 519.840 ;
        RECT 4.000 516.440 894.065 517.840 ;
        RECT 4.000 514.440 894.465 516.440 ;
        RECT 4.400 513.040 894.465 514.440 ;
        RECT 4.000 511.040 894.465 513.040 ;
        RECT 4.000 509.640 894.065 511.040 ;
        RECT 4.000 507.640 894.465 509.640 ;
        RECT 4.400 506.240 894.465 507.640 ;
        RECT 4.000 504.240 894.465 506.240 ;
        RECT 4.000 502.840 894.065 504.240 ;
        RECT 4.000 500.840 894.465 502.840 ;
        RECT 4.400 499.440 894.465 500.840 ;
        RECT 4.000 497.440 894.465 499.440 ;
        RECT 4.000 496.040 894.065 497.440 ;
        RECT 4.000 490.640 894.465 496.040 ;
        RECT 4.400 489.240 894.065 490.640 ;
        RECT 4.000 483.840 894.465 489.240 ;
        RECT 4.400 482.440 894.065 483.840 ;
        RECT 4.000 477.040 894.465 482.440 ;
        RECT 4.400 475.640 894.065 477.040 ;
        RECT 4.000 470.240 894.465 475.640 ;
        RECT 4.400 468.840 894.065 470.240 ;
        RECT 4.000 463.440 894.465 468.840 ;
        RECT 4.400 462.040 894.065 463.440 ;
        RECT 4.000 456.640 894.465 462.040 ;
        RECT 4.400 455.240 894.065 456.640 ;
        RECT 4.000 449.840 894.465 455.240 ;
        RECT 4.400 448.440 894.065 449.840 ;
        RECT 4.000 443.040 894.465 448.440 ;
        RECT 4.400 441.640 894.065 443.040 ;
        RECT 4.000 436.240 894.465 441.640 ;
        RECT 4.400 434.840 894.065 436.240 ;
        RECT 4.000 429.440 894.465 434.840 ;
        RECT 4.400 428.040 894.065 429.440 ;
        RECT 4.000 422.640 894.465 428.040 ;
        RECT 4.400 421.240 894.065 422.640 ;
        RECT 4.000 415.840 894.465 421.240 ;
        RECT 4.400 414.440 894.065 415.840 ;
        RECT 4.000 409.040 894.465 414.440 ;
        RECT 4.400 407.640 894.465 409.040 ;
        RECT 4.000 405.640 894.465 407.640 ;
        RECT 4.000 404.240 894.065 405.640 ;
        RECT 4.000 402.240 894.465 404.240 ;
        RECT 4.400 400.840 894.465 402.240 ;
        RECT 4.000 398.840 894.465 400.840 ;
        RECT 4.000 397.440 894.065 398.840 ;
        RECT 4.000 395.440 894.465 397.440 ;
        RECT 4.400 394.040 894.465 395.440 ;
        RECT 4.000 392.040 894.465 394.040 ;
        RECT 4.000 390.640 894.065 392.040 ;
        RECT 4.000 388.640 894.465 390.640 ;
        RECT 4.400 387.240 894.465 388.640 ;
        RECT 4.000 385.240 894.465 387.240 ;
        RECT 4.000 383.840 894.065 385.240 ;
        RECT 4.000 381.840 894.465 383.840 ;
        RECT 4.400 380.440 894.465 381.840 ;
        RECT 4.000 378.440 894.465 380.440 ;
        RECT 4.000 377.040 894.065 378.440 ;
        RECT 4.000 371.640 894.465 377.040 ;
        RECT 4.400 370.240 894.065 371.640 ;
        RECT 4.000 364.840 894.465 370.240 ;
        RECT 4.400 363.440 894.065 364.840 ;
        RECT 4.000 358.040 894.465 363.440 ;
        RECT 4.400 356.640 894.065 358.040 ;
        RECT 4.000 351.240 894.465 356.640 ;
        RECT 4.400 349.840 894.065 351.240 ;
        RECT 4.000 344.440 894.465 349.840 ;
        RECT 4.400 343.040 894.065 344.440 ;
        RECT 4.000 337.640 894.465 343.040 ;
        RECT 4.400 336.240 894.065 337.640 ;
        RECT 4.000 330.840 894.465 336.240 ;
        RECT 4.400 329.440 894.065 330.840 ;
        RECT 4.000 324.040 894.465 329.440 ;
        RECT 4.400 322.640 894.065 324.040 ;
        RECT 4.000 317.240 894.465 322.640 ;
        RECT 4.400 315.840 894.065 317.240 ;
        RECT 4.000 310.440 894.465 315.840 ;
        RECT 4.400 309.040 894.065 310.440 ;
        RECT 4.000 303.640 894.465 309.040 ;
        RECT 4.400 302.240 894.065 303.640 ;
        RECT 4.000 296.840 894.465 302.240 ;
        RECT 4.400 295.440 894.065 296.840 ;
        RECT 4.000 290.040 894.465 295.440 ;
        RECT 4.400 288.640 894.465 290.040 ;
        RECT 4.000 286.640 894.465 288.640 ;
        RECT 4.000 285.240 894.065 286.640 ;
        RECT 4.000 283.240 894.465 285.240 ;
        RECT 4.400 281.840 894.465 283.240 ;
        RECT 4.000 279.840 894.465 281.840 ;
        RECT 4.000 278.440 894.065 279.840 ;
        RECT 4.000 276.440 894.465 278.440 ;
        RECT 4.400 275.040 894.465 276.440 ;
        RECT 4.000 273.040 894.465 275.040 ;
        RECT 4.000 271.640 894.065 273.040 ;
        RECT 4.000 269.640 894.465 271.640 ;
        RECT 4.400 268.240 894.465 269.640 ;
        RECT 4.000 266.240 894.465 268.240 ;
        RECT 4.000 264.840 894.065 266.240 ;
        RECT 4.000 262.840 894.465 264.840 ;
        RECT 4.400 261.440 894.465 262.840 ;
        RECT 4.000 259.440 894.465 261.440 ;
        RECT 4.000 258.040 894.065 259.440 ;
        RECT 4.000 256.040 894.465 258.040 ;
        RECT 4.400 254.640 894.465 256.040 ;
        RECT 4.000 252.640 894.465 254.640 ;
        RECT 4.000 251.240 894.065 252.640 ;
        RECT 4.000 245.840 894.465 251.240 ;
        RECT 4.400 244.440 894.065 245.840 ;
        RECT 4.000 239.040 894.465 244.440 ;
        RECT 4.400 237.640 894.065 239.040 ;
        RECT 4.000 232.240 894.465 237.640 ;
        RECT 4.400 230.840 894.065 232.240 ;
        RECT 4.000 225.440 894.465 230.840 ;
        RECT 4.400 224.040 894.065 225.440 ;
        RECT 4.000 218.640 894.465 224.040 ;
        RECT 4.400 217.240 894.065 218.640 ;
        RECT 4.000 211.840 894.465 217.240 ;
        RECT 4.400 210.440 894.065 211.840 ;
        RECT 4.000 205.040 894.465 210.440 ;
        RECT 4.400 203.640 894.065 205.040 ;
        RECT 4.000 198.240 894.465 203.640 ;
        RECT 4.400 196.840 894.065 198.240 ;
        RECT 4.000 191.440 894.465 196.840 ;
        RECT 4.400 190.040 894.065 191.440 ;
        RECT 4.000 184.640 894.465 190.040 ;
        RECT 4.400 183.240 894.065 184.640 ;
        RECT 4.000 177.840 894.465 183.240 ;
        RECT 4.400 176.440 894.065 177.840 ;
        RECT 4.000 171.040 894.465 176.440 ;
        RECT 4.400 169.640 894.065 171.040 ;
        RECT 4.000 164.240 894.465 169.640 ;
        RECT 4.400 162.840 894.465 164.240 ;
        RECT 4.000 160.840 894.465 162.840 ;
        RECT 4.000 159.440 894.065 160.840 ;
        RECT 4.000 157.440 894.465 159.440 ;
        RECT 4.400 156.040 894.465 157.440 ;
        RECT 4.000 154.040 894.465 156.040 ;
        RECT 4.000 152.640 894.065 154.040 ;
        RECT 4.000 150.640 894.465 152.640 ;
        RECT 4.400 149.240 894.465 150.640 ;
        RECT 4.000 147.240 894.465 149.240 ;
        RECT 4.000 145.840 894.065 147.240 ;
        RECT 4.000 143.840 894.465 145.840 ;
        RECT 4.400 142.440 894.465 143.840 ;
        RECT 4.000 140.440 894.465 142.440 ;
        RECT 4.000 139.040 894.065 140.440 ;
        RECT 4.000 137.040 894.465 139.040 ;
        RECT 4.400 135.640 894.465 137.040 ;
        RECT 4.000 133.640 894.465 135.640 ;
        RECT 4.000 132.240 894.065 133.640 ;
        RECT 4.000 130.240 894.465 132.240 ;
        RECT 4.400 128.840 894.465 130.240 ;
        RECT 4.000 126.840 894.465 128.840 ;
        RECT 4.000 125.440 894.065 126.840 ;
        RECT 4.000 120.040 894.465 125.440 ;
        RECT 4.400 118.640 894.065 120.040 ;
        RECT 4.000 113.240 894.465 118.640 ;
        RECT 4.400 111.840 894.065 113.240 ;
        RECT 4.000 106.440 894.465 111.840 ;
        RECT 4.400 105.040 894.065 106.440 ;
        RECT 4.000 99.640 894.465 105.040 ;
        RECT 4.400 98.240 894.065 99.640 ;
        RECT 4.000 92.840 894.465 98.240 ;
        RECT 4.400 91.440 894.065 92.840 ;
        RECT 4.000 86.040 894.465 91.440 ;
        RECT 4.400 84.640 894.065 86.040 ;
        RECT 4.000 79.240 894.465 84.640 ;
        RECT 4.400 77.840 894.065 79.240 ;
        RECT 4.000 72.440 894.465 77.840 ;
        RECT 4.400 71.040 894.065 72.440 ;
        RECT 4.000 65.640 894.465 71.040 ;
        RECT 4.400 64.240 894.065 65.640 ;
        RECT 4.000 58.840 894.465 64.240 ;
        RECT 4.400 57.440 894.065 58.840 ;
        RECT 4.000 52.040 894.465 57.440 ;
        RECT 4.400 50.640 894.065 52.040 ;
        RECT 4.000 45.240 894.465 50.640 ;
        RECT 4.400 43.840 894.065 45.240 ;
        RECT 4.000 38.440 894.465 43.840 ;
        RECT 4.400 37.040 894.465 38.440 ;
        RECT 4.000 35.040 894.465 37.040 ;
        RECT 4.000 33.640 894.065 35.040 ;
        RECT 4.000 31.640 894.465 33.640 ;
        RECT 4.400 30.240 894.465 31.640 ;
        RECT 4.000 28.240 894.465 30.240 ;
        RECT 4.000 26.840 894.065 28.240 ;
        RECT 4.000 24.840 894.465 26.840 ;
        RECT 4.400 23.440 894.465 24.840 ;
        RECT 4.000 21.440 894.465 23.440 ;
        RECT 4.000 20.040 894.065 21.440 ;
        RECT 4.000 18.040 894.465 20.040 ;
        RECT 4.400 16.640 894.465 18.040 ;
        RECT 4.000 14.640 894.465 16.640 ;
        RECT 4.000 13.240 894.065 14.640 ;
        RECT 4.000 11.240 894.465 13.240 ;
        RECT 4.400 9.840 894.465 11.240 ;
        RECT 4.000 7.840 894.465 9.840 ;
        RECT 4.000 6.975 894.065 7.840 ;
      LAYER met4 ;
        RECT 16.855 15.135 21.620 889.945 ;
        RECT 25.420 15.135 39.620 889.945 ;
        RECT 43.420 15.135 57.620 889.945 ;
        RECT 61.420 15.135 93.620 889.945 ;
        RECT 97.420 15.135 111.620 889.945 ;
        RECT 115.420 15.135 129.620 889.945 ;
        RECT 133.420 15.135 147.620 889.945 ;
        RECT 151.420 15.135 183.620 889.945 ;
        RECT 187.420 15.135 201.620 889.945 ;
        RECT 205.420 15.135 219.620 889.945 ;
        RECT 223.420 15.135 237.620 889.945 ;
        RECT 241.420 15.135 273.620 889.945 ;
        RECT 277.420 15.135 291.620 889.945 ;
        RECT 295.420 15.135 309.620 889.945 ;
        RECT 313.420 15.135 327.620 889.945 ;
        RECT 331.420 15.135 363.620 889.945 ;
        RECT 367.420 15.135 381.620 889.945 ;
        RECT 385.420 15.135 399.620 889.945 ;
        RECT 403.420 15.135 417.620 889.945 ;
        RECT 421.420 15.135 453.620 889.945 ;
        RECT 457.420 15.135 471.620 889.945 ;
        RECT 475.420 15.135 489.620 889.945 ;
        RECT 493.420 15.135 507.620 889.945 ;
        RECT 511.420 15.135 543.620 889.945 ;
        RECT 547.420 15.135 561.620 889.945 ;
        RECT 565.420 15.135 579.620 889.945 ;
        RECT 583.420 15.135 597.620 889.945 ;
        RECT 601.420 15.135 633.620 889.945 ;
        RECT 637.420 15.135 651.620 889.945 ;
        RECT 655.420 15.135 669.620 889.945 ;
        RECT 673.420 15.135 687.620 889.945 ;
        RECT 691.420 15.135 723.620 889.945 ;
        RECT 727.420 15.135 741.620 889.945 ;
        RECT 745.420 15.135 759.620 889.945 ;
        RECT 763.420 15.135 777.620 889.945 ;
        RECT 781.420 15.135 813.620 889.945 ;
        RECT 817.420 15.135 826.785 889.945 ;
      LAYER met5 ;
        RECT -42.880 946.000 -39.880 946.010 ;
        RECT 148.020 946.000 151.020 946.010 ;
        RECT 328.020 946.000 331.020 946.010 ;
        RECT 508.020 946.000 511.020 946.010 ;
        RECT 688.020 946.000 691.020 946.010 ;
        RECT 868.020 946.000 871.020 946.010 ;
        RECT 938.260 946.000 941.260 946.010 ;
        RECT -42.880 942.990 -39.880 943.000 ;
        RECT 148.020 942.990 151.020 943.000 ;
        RECT 328.020 942.990 331.020 943.000 ;
        RECT 508.020 942.990 511.020 943.000 ;
        RECT 688.020 942.990 691.020 943.000 ;
        RECT 868.020 942.990 871.020 943.000 ;
        RECT 938.260 942.990 941.260 943.000 ;
        RECT -38.180 941.300 -35.180 941.310 ;
        RECT 58.020 941.300 61.020 941.310 ;
        RECT 238.020 941.300 241.020 941.310 ;
        RECT 418.020 941.300 421.020 941.310 ;
        RECT 598.020 941.300 601.020 941.310 ;
        RECT 778.020 941.300 781.020 941.310 ;
        RECT 933.560 941.300 936.560 941.310 ;
        RECT -38.180 938.290 -35.180 938.300 ;
        RECT 58.020 938.290 61.020 938.300 ;
        RECT 238.020 938.290 241.020 938.300 ;
        RECT 418.020 938.290 421.020 938.300 ;
        RECT 598.020 938.290 601.020 938.300 ;
        RECT 778.020 938.290 781.020 938.300 ;
        RECT 933.560 938.290 936.560 938.300 ;
        RECT -33.480 936.600 -30.480 936.610 ;
        RECT 130.020 936.600 133.020 936.610 ;
        RECT 310.020 936.600 313.020 936.610 ;
        RECT 490.020 936.600 493.020 936.610 ;
        RECT 670.020 936.600 673.020 936.610 ;
        RECT 850.020 936.600 853.020 936.610 ;
        RECT 928.860 936.600 931.860 936.610 ;
        RECT -33.480 933.590 -30.480 933.600 ;
        RECT 130.020 933.590 133.020 933.600 ;
        RECT 310.020 933.590 313.020 933.600 ;
        RECT 490.020 933.590 493.020 933.600 ;
        RECT 670.020 933.590 673.020 933.600 ;
        RECT 850.020 933.590 853.020 933.600 ;
        RECT 928.860 933.590 931.860 933.600 ;
        RECT -28.780 931.900 -25.780 931.910 ;
        RECT 40.020 931.900 43.020 931.910 ;
        RECT 220.020 931.900 223.020 931.910 ;
        RECT 400.020 931.900 403.020 931.910 ;
        RECT 580.020 931.900 583.020 931.910 ;
        RECT 760.020 931.900 763.020 931.910 ;
        RECT 924.160 931.900 927.160 931.910 ;
        RECT -28.780 928.890 -25.780 928.900 ;
        RECT 40.020 928.890 43.020 928.900 ;
        RECT 220.020 928.890 223.020 928.900 ;
        RECT 400.020 928.890 403.020 928.900 ;
        RECT 580.020 928.890 583.020 928.900 ;
        RECT 760.020 928.890 763.020 928.900 ;
        RECT 924.160 928.890 927.160 928.900 ;
        RECT -24.080 927.200 -21.080 927.210 ;
        RECT 112.020 927.200 115.020 927.210 ;
        RECT 292.020 927.200 295.020 927.210 ;
        RECT 472.020 927.200 475.020 927.210 ;
        RECT 652.020 927.200 655.020 927.210 ;
        RECT 832.020 927.200 835.020 927.210 ;
        RECT 919.460 927.200 922.460 927.210 ;
        RECT -24.080 924.190 -21.080 924.200 ;
        RECT 112.020 924.190 115.020 924.200 ;
        RECT 292.020 924.190 295.020 924.200 ;
        RECT 472.020 924.190 475.020 924.200 ;
        RECT 652.020 924.190 655.020 924.200 ;
        RECT 832.020 924.190 835.020 924.200 ;
        RECT 919.460 924.190 922.460 924.200 ;
        RECT -19.380 922.500 -16.380 922.510 ;
        RECT 22.020 922.500 25.020 922.510 ;
        RECT 202.020 922.500 205.020 922.510 ;
        RECT 382.020 922.500 385.020 922.510 ;
        RECT 562.020 922.500 565.020 922.510 ;
        RECT 742.020 922.500 745.020 922.510 ;
        RECT 914.760 922.500 917.760 922.510 ;
        RECT -19.380 919.490 -16.380 919.500 ;
        RECT 22.020 919.490 25.020 919.500 ;
        RECT 202.020 919.490 205.020 919.500 ;
        RECT 382.020 919.490 385.020 919.500 ;
        RECT 562.020 919.490 565.020 919.500 ;
        RECT 742.020 919.490 745.020 919.500 ;
        RECT 914.760 919.490 917.760 919.500 ;
        RECT -14.680 917.800 -11.680 917.810 ;
        RECT 94.020 917.800 97.020 917.810 ;
        RECT 274.020 917.800 277.020 917.810 ;
        RECT 454.020 917.800 457.020 917.810 ;
        RECT 634.020 917.800 637.020 917.810 ;
        RECT 814.020 917.800 817.020 917.810 ;
        RECT 910.060 917.800 913.060 917.810 ;
        RECT -14.680 914.790 -11.680 914.800 ;
        RECT 94.020 914.790 97.020 914.800 ;
        RECT 274.020 914.790 277.020 914.800 ;
        RECT 454.020 914.790 457.020 914.800 ;
        RECT 634.020 914.790 637.020 914.800 ;
        RECT 814.020 914.790 817.020 914.800 ;
        RECT 910.060 914.790 913.060 914.800 ;
        RECT -9.980 913.100 -6.980 913.110 ;
        RECT 4.020 913.100 7.020 913.110 ;
        RECT 184.020 913.100 187.020 913.110 ;
        RECT 364.020 913.100 367.020 913.110 ;
        RECT 544.020 913.100 547.020 913.110 ;
        RECT 724.020 913.100 727.020 913.110 ;
        RECT 905.360 913.100 908.360 913.110 ;
        RECT -9.980 910.090 -6.980 910.100 ;
        RECT 4.020 910.090 7.020 910.100 ;
        RECT 184.020 910.090 187.020 910.100 ;
        RECT 364.020 910.090 367.020 910.100 ;
        RECT 544.020 910.090 547.020 910.100 ;
        RECT 724.020 910.090 727.020 910.100 ;
        RECT 905.360 910.090 908.360 910.100 ;
        RECT 0.000 877.980 898.465 908.500 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 938.260 876.380 941.260 876.390 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 938.260 873.370 941.260 873.380 ;
        RECT 0.000 859.980 898.465 871.780 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 928.860 858.380 931.860 858.390 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 928.860 855.370 931.860 855.380 ;
        RECT 0.000 841.980 898.465 853.780 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 919.460 840.380 922.460 840.390 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 919.460 837.370 922.460 837.380 ;
        RECT 0.000 823.740 898.465 835.780 ;
        RECT -14.680 822.140 -11.680 822.150 ;
        RECT 910.060 822.140 913.060 822.150 ;
        RECT -14.680 819.130 -11.680 819.140 ;
        RECT 910.060 819.130 913.060 819.140 ;
        RECT 0.000 787.980 898.465 817.540 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 933.560 786.380 936.560 786.390 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 933.560 783.370 936.560 783.380 ;
        RECT 0.000 769.980 898.465 781.780 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 924.160 768.380 927.160 768.390 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 924.160 765.370 927.160 765.380 ;
        RECT 0.000 751.980 898.465 763.780 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 914.760 750.380 917.760 750.390 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 914.760 747.370 917.760 747.380 ;
        RECT 0.000 733.740 898.465 745.780 ;
        RECT -9.980 732.140 -6.980 732.150 ;
        RECT 905.360 732.140 908.360 732.150 ;
        RECT -9.980 729.130 -6.980 729.140 ;
        RECT 905.360 729.130 908.360 729.140 ;
        RECT 0.000 697.980 898.465 727.540 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 938.260 696.380 941.260 696.390 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 938.260 693.370 941.260 693.380 ;
        RECT 0.000 679.980 898.465 691.780 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 928.860 678.380 931.860 678.390 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 928.860 675.370 931.860 675.380 ;
        RECT 0.000 661.980 898.465 673.780 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 919.460 660.380 922.460 660.390 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 919.460 657.370 922.460 657.380 ;
        RECT 0.000 643.740 898.465 655.780 ;
        RECT -14.680 642.140 -11.680 642.150 ;
        RECT 910.060 642.140 913.060 642.150 ;
        RECT -14.680 639.130 -11.680 639.140 ;
        RECT 910.060 639.130 913.060 639.140 ;
        RECT 0.000 607.980 898.465 637.540 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 933.560 606.380 936.560 606.390 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 933.560 603.370 936.560 603.380 ;
        RECT 0.000 589.980 898.465 601.780 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 924.160 588.380 927.160 588.390 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 924.160 585.370 927.160 585.380 ;
        RECT 0.000 571.980 898.465 583.780 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 914.760 570.380 917.760 570.390 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 914.760 567.370 917.760 567.380 ;
        RECT 0.000 553.740 898.465 565.780 ;
        RECT -9.980 552.140 -6.980 552.150 ;
        RECT 905.360 552.140 908.360 552.150 ;
        RECT -9.980 549.130 -6.980 549.140 ;
        RECT 905.360 549.130 908.360 549.140 ;
        RECT 0.000 517.980 898.465 547.540 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 938.260 516.380 941.260 516.390 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 938.260 513.370 941.260 513.380 ;
        RECT 0.000 499.980 898.465 511.780 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 928.860 498.380 931.860 498.390 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 928.860 495.370 931.860 495.380 ;
        RECT 0.000 481.980 898.465 493.780 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 919.460 480.380 922.460 480.390 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 919.460 477.370 922.460 477.380 ;
        RECT 0.000 463.740 898.465 475.780 ;
        RECT -14.680 462.140 -11.680 462.150 ;
        RECT 910.060 462.140 913.060 462.150 ;
        RECT -14.680 459.130 -11.680 459.140 ;
        RECT 910.060 459.130 913.060 459.140 ;
        RECT 0.000 427.980 898.465 457.540 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 933.560 426.380 936.560 426.390 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 933.560 423.370 936.560 423.380 ;
        RECT 0.000 409.980 898.465 421.780 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 924.160 408.380 927.160 408.390 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 924.160 405.370 927.160 405.380 ;
        RECT 0.000 391.980 898.465 403.780 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 914.760 390.380 917.760 390.390 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 914.760 387.370 917.760 387.380 ;
        RECT 0.000 373.740 898.465 385.780 ;
        RECT -9.980 372.140 -6.980 372.150 ;
        RECT 905.360 372.140 908.360 372.150 ;
        RECT -9.980 369.130 -6.980 369.140 ;
        RECT 905.360 369.130 908.360 369.140 ;
        RECT 0.000 337.980 898.465 367.540 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 938.260 336.380 941.260 336.390 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 938.260 333.370 941.260 333.380 ;
        RECT 0.000 319.980 898.465 331.780 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 928.860 318.380 931.860 318.390 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 928.860 315.370 931.860 315.380 ;
        RECT 0.000 301.980 898.465 313.780 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 919.460 300.380 922.460 300.390 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 919.460 297.370 922.460 297.380 ;
        RECT 0.000 283.740 898.465 295.780 ;
        RECT -14.680 282.140 -11.680 282.150 ;
        RECT 910.060 282.140 913.060 282.150 ;
        RECT -14.680 279.130 -11.680 279.140 ;
        RECT 910.060 279.130 913.060 279.140 ;
        RECT 0.000 247.980 898.465 277.540 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 933.560 246.380 936.560 246.390 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 933.560 243.370 936.560 243.380 ;
        RECT 0.000 229.980 898.465 241.780 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 924.160 228.380 927.160 228.390 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 924.160 225.370 927.160 225.380 ;
        RECT 0.000 211.980 898.465 223.780 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 914.760 210.380 917.760 210.390 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 914.760 207.370 917.760 207.380 ;
        RECT 0.000 193.740 898.465 205.780 ;
        RECT -9.980 192.140 -6.980 192.150 ;
        RECT 905.360 192.140 908.360 192.150 ;
        RECT -9.980 189.130 -6.980 189.140 ;
        RECT 905.360 189.130 908.360 189.140 ;
        RECT 0.000 157.980 898.465 187.540 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 938.260 156.380 941.260 156.390 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 938.260 153.370 941.260 153.380 ;
        RECT 0.000 139.980 898.465 151.780 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 928.860 138.380 931.860 138.390 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 928.860 135.370 931.860 135.380 ;
        RECT 0.000 121.980 898.465 133.780 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 919.460 120.380 922.460 120.390 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 919.460 117.370 922.460 117.380 ;
        RECT 0.000 103.740 898.465 115.780 ;
        RECT -14.680 102.140 -11.680 102.150 ;
        RECT 910.060 102.140 913.060 102.150 ;
        RECT -14.680 99.130 -11.680 99.140 ;
        RECT 910.060 99.130 913.060 99.140 ;
        RECT 0.000 67.980 898.465 97.540 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 933.560 66.380 936.560 66.390 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 933.560 63.370 936.560 63.380 ;
        RECT 0.000 49.980 898.465 61.780 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 924.160 48.380 927.160 48.390 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 924.160 45.370 927.160 45.380 ;
        RECT 0.000 31.980 898.465 43.780 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 914.760 30.380 917.760 30.390 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 914.760 27.370 917.760 27.380 ;
        RECT 0.000 13.740 898.465 25.780 ;
        RECT -9.980 12.140 -6.980 12.150 ;
        RECT 905.360 12.140 908.360 12.150 ;
        RECT -9.980 9.130 -6.980 9.140 ;
        RECT 905.360 9.130 908.360 9.140 ;
        RECT 0.000 0.000 898.465 7.540 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 905.360 -1.620 908.360 -1.610 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 905.360 -4.630 908.360 -4.620 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 910.060 -6.320 913.060 -6.310 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 910.060 -9.330 913.060 -9.320 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 914.760 -11.020 917.760 -11.010 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 914.760 -14.030 917.760 -14.020 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 919.460 -15.720 922.460 -15.710 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 919.460 -18.730 922.460 -18.720 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 924.160 -20.420 927.160 -20.410 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 924.160 -23.430 927.160 -23.420 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 928.860 -25.120 931.860 -25.110 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 928.860 -28.130 931.860 -28.120 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 933.560 -29.820 936.560 -29.810 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 933.560 -32.830 936.560 -32.820 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 938.260 -34.520 941.260 -34.510 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 938.260 -37.530 941.260 -37.520 ;
  END
END user_project_wrapper
END LIBRARY

